��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8����"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v�Ӛ�U
�"���3�v������/$��C~a�TS��=��W��z�yW�9M��4R؞+�HR�|OZ�=���.OL11b���䍟5o�HF�pw��%�U	��+.�jw���٬�������O�X�Z�����]g*��s>�ql���U!����[�D����r?�M �®�m�;Y�+��م�HK8D;���p�E����yʵT��7ӹC��fD����NwR�S(l���ے��J�R���d�������?�.2�P�)O����գ����)�uVS���Ԁj#L֏3�����l+�o(��3�!ٿ>N�^Y(K�j�r�(�I+(��k�o��X��4A>h�]�k�e��A����,�'�F_H[q)|{���7hE_&��+Մ����i��`�0��_��]��(���h#`��h��2sK�Nl��b�v��/}i��2�T.��i[e�-<����f.J����� ��ě�:/��$�2[��.��F4��v?]0A��`�ђ�W7"�
���G��0�H��k�e�'51ȝF�����+l��ұSA��	�uҟc��AK20�&B{��G�}K���U֩ҋi�;2� e.�.��q[��D@H��~{L=��GOtM���g���ۣ�kj�c92�>���煒����<����I~Q˲�F��$`��7r�2�<���#١��0�Co�T��u�2)���>S[UD;���P��Юf�7Vd���m޶���VB�����sx/�1�oU����<�9�#@P��j����o���Lҽ���J�ɪexˁ|�2���@/զ�ļ����!
�OFvV�k�3�Ξ��=���,a�h]�R�����*U��W���a���Cb�I�0��N��zM�h��fJ�9���t��:(=��N��ז�U��c�Y8��ej앋z:)�-��ic�� �|�>4(��=^��]����6.����)��_~��&+��:�B�H���+u)\<�E�v�28���
��\Ï���n���08�>�w������|��K�{Y/B�o�o�J�������k^�V� �R�.ߒT޺I�ekÒ��@�m����*�k���DD�F��>3BC]�hY�;�z�����`@��Xd�.gop@�n�-<�W��z��Op˗,��0G����@����n�����>�i�.pu��6	�d��ԴS1����'��Ou^Fs���aYP���5�}N6�\f�$�/:���͖��r���QmA#:���я��z�,z�uHJ\��FNg(�����{��\�g5�Fo?(^�����!y�F9-%�ś.C|����b�f��!�p5�+�A�,�JO��[+��M�'ޕ7�mz�k�Н��?�Z=�qV�!�2�$�\�1�n���]`A-��D�'G�:*��#���ϨL�l�w(u����}�P�b��rp�°�yj��5* �Jg>1��~���WOQ�D�a�
��i�1;�@���!?�`Y�W��:V8�c�&Ĝ>�y!m!�M�)�*b+�*^��;X�g[���B���<^2g����$�S-	iI�]���=h}*�U�}���@㶊~��+5��Z�8]�:���`�����(�=���w]Tq���͎b[�r0�ۧ1(�c&�6ʈ.��>*�"p)N0ܶ���N,~=o}Ӎ��Sd�+��24ʓ.(tz�O|�����3�<S�D�Q]�䬩����~���N�K���пƙ-Z,x�8J�|��ŝBgNC�^M�Pt�η3��[p��<����.l�X���i+��7˰�����:�pDn����e<+=51B���)�ߙ����g�[���)b��Ǡ�Z�i~ƀ��E�T��!�7����b���r����}v�s���˨P޿�m��]wȁ�R��@b����P�2��<4$w���͕�p�:N&�L�I���_���pn��UK�k���j��!�Вjգ�����pp�6Pi�R�>�����6�gD��OXk+=�M�<��^��׬Q y�9�m!�yQ3
��� u�)�:�l�*���'+O�_���|'7y��3[L��T<�Ù��N�o��e�����K�V�o��e�g��]T������S�>3>N������`�ԓɿ(�z�-l�q츏3��G]�d�,u��?MS�Z�L�Pg���ﰊ�T�}�-.>��#��ذ�x�~�[�{�N��,���"�k��UE�;�(�_u�ʈ)�B:#�%a�ДbYZCg�ppm�V�Q�ܺ����A{�>�P�d�i᝾$u��nQ.�u�[�g�E)��#3�Ns��F@eO�j�G/�0��p͌��3�>��=p/��D!�&�S+��3�w>�cڼy_um�B69g(�����ls�"j~,��}��7H�L�:��!��(�g����e H�U[˻�]_F�D6��*&�׬���c�i�g��`T4p�i�,��SЁ�Y���0h�1%^)k>�TN���%_^ۋ���\�bTu�'����[� �'�H1�ό��r��NRA�g���5C�������[-���*Yd�N�w������T�Q*[��M��� �Z������N�l�kd�n�c_�d� �����	(��g�����m�rO0l
k�)8�Pf��U�V�׽2r(��xp�J/+N!����Ԏ1��瘲�4��BM�x˹<?}�,�ـv���#�Y�N�'�jl*�;;��⫾8>�@d]�rW��}B"ݤ�ѧ<���ox���d��t��o�dc:@��R
e�:V�����)�iX�Y!�T��`
0�N��r�{�7Dr���W����E�]��jn�O8�--B��D�T-iBs��DDj�����̧���YS��^�ͺޒ�
�#K���)�����Ĉ 4\X��E�aY����G�q��D��e�)M�s�`��f;� �������2�;������w��%J�J\3.����Iz�)iC�r���1��h�"9��oE����c���G~�;a�LE�yB)�������+�1���L݃�v����U.�t�mX�'�r0G���ˣ콐�\ݘ�H����,�(���ZG�*},M��I����Ddl��)H�!ő4:���4�w���_�Fs_������y�a��/%ѱ�gG��^���=tUx~&E�\]|��x��h��/����Wt�g�V��@�G�WV���օw�Tk�$0���S���$�X�֏��6㌞�����e߇>�:��-e{֑�ѵ������AN�/�c�{�W>�r�(�5�T�j[�%�_Ѳ��ؽG������Q]>nH�͡����>H9�q>�_�- �$��ީ^�S�&�g�I�:b�n������E:��
�>��ߛ�����]��p:�à�&���`������p��_=��=�f�]"t҃����30<1�%}H0�X*��=��1�\B�;:���&`D���J��Lsh"�sv��t�g	��	�XS��R0�1��i~����͜I�P��+�w,�)OjR����-�����~���
����#��<���R�[��zZ�J��hʽ�*¡��}HE;3��:��g��f1툤�]�_����`&�\�:�>7r��I�i������+b���f)�!YB[4Ba�W���g1E��+-��Uy��f=�z�; ���;�~�	!��ki�lɝ��6�'BB�$.I���ՠ?���ZP4\-1��Z����L��Q�"�j�`evd�#!��q+[�~^4'��~Tg��ho�6rwѿ�����b<�g�!՚��a�+�\��c��RoJ�X}�H�o�����XX&!�������G+Hl$A9��bl5|�'v�z6��">���_�uj����y�3,�U8���95a��=�G���k�.l\���p�э�Ly?�Z�c�����-K�I0�v '���ynZV7��6%��7���g�����̹ݿ�������i��.�$z)�h~�l���
��g�ۏ�=��B=S@6���)�$�8��S�C�+�7pu����=�_,�VʰU(k�Ccz[,�y�-�e	g���\^T�P���s�=P����N��q�Ň�0�sR_��V�u"^�c!�l
@�s1(�,vuV��־":He������	R���S����,��eWَ,֩��ov�F�R���<�%��-����In�,9������F7��R��^&�*�4����_��Kc�Lּ���*q\:r ��(I�{d!fǰ���E=LK:�_/X�O���up+W��d�Ͷ%6nԷ\O��e�0Cr3f'pH/�72�A��I+0o�Qŭn	��v�'�`c��p�T��,Ԛ��R�������=�`�ˑ�,jR�ߚ�6�)
�ϱhi�(q}<�ec�gMx�t�MM֕�Ƞ
��D��'�lͅ��`Dz���6{>�,"X"L�;`�M��S�3��i��^e�	w���|�E���K1b�ڈ�n�GX=�� ��g11�F���geA
�H��O��&����pa/Y�%��H�{r�ZS���dV���T	��~��t˵w#����[n ��q�]1�T#�<"k_��z�u
Ҕ� ,�u����G���nb��=�YMM��q͜�$�U�Quhv-Ի�u���AD�5�P�L��`�V۩�!t�+���)�Vg�y�W�y���u��ŵ�� ��ރs�X��aN8�^�z��$�ߕ?�yP����1*Þ,?�L��~��XJ���*��p�5z�kl� ���n���N]�ײL
T���C�1��9�� 	���땫��ڼ		ܙ��Uj��{X�r$9=>=$n ���~�D3��cd��ݕ��z<v?�ԻI9����@�$�g�Uz�g������ЇhHod7��B_�R�c�%|4K�}i�]{j�l�/'_c{�{�%���D���_nQh��s��+{*��)�Ey,���5�����)�1K����ë����=��y�IWr�R|G:F�|0��zOaN�x&Du��NAȜ/�NY��9���'���z��g:/h���4�hgH�
}�}�EK��)�����t���\���Ć���8�WѼs$B&�����h�	��9��6��g骦_�b�"Y0���Ro�]��]�u�)a7m͑��P�AoeHUZ*a�1��I{S���]Ć��9W�[�'b�uF��F�|�,\CH��7Q��+�����U�)l��l���sQ��@�|��b���u�
:��c�Bl=r+x@�*7�[�;���ě�z���8~���&n(En� ^�0�<�y�#�����v�ux0=��\R���Tl��Q��rR2�T��>E|�h}.����[�xt�D�\��zXL�wRc�6FJq5qw>�)VLR�b1Q^�qX�̥�>5]׸!�V�j��QIp���)i�És�����ubY�B�����K��r�Z��r>��P�m�A4�ʎ�{�t��XoJ(9,������8��*����\������d�e��_b���7AM=�5ٻ�h;;F�,T�XI�������4�!��MN6���?��hp�O��@�ƞ��D�+��M�;:�O%���@s6��vq�y��M=R}�գ�i�n䍖��\R�u��|3����E�|�Wt��	�2+���Γ��Pv�uh�T���jܔ�a��� ����-��6ȕ\�|�S1Mz���'r%��|�MN9��Z�rI���<��Q�M� ��)��L�c�c��J��.��8]H����y��z�W,������bC����3Pz�(��k���'EG(�z�*Y_�%��BTmy�!�ę����*|
X�K�V��q����o��<�{��0��)L��~rd_�q������{�%�ReI�k�F��/B�i8Z�$ ͈���n��5
��tэM��f��+��^����*��(�-�\��:�!��>GT)���˕eY������2�%>�4�>S�g���9�>"@=�� �Utܞ����@�訋tU�(	k�V����H�Ȅҏ�vPJ��<�v�&.�ekC�<��/�>\�%�ϥ�������}S�X�;�o\���,�� �x����|�k[�.�d���GrI|�\�@dh��m���/F��`�U��M��7�`�.�
�!5���!�-��߭�������2mz9�h�5��;�I�p�-�*��B��]ֻB9��o
�� X�t0}̗��>.k�,'4/=��Pv�G%�yd�!S�oE|�Hv�H�l��/Av>"�YCo��h8Y����N��.����S�x�)!ݑ�tl�׏O�.��p1��4*P�����0k����p���eՎ���G-���T%��-I�0���1�{3q�;N��c��u�s�n�l������d��2i��ӿ��� ��=4v�	����K��:]y�$2�F4�� ;΃Ëqa�1Ĵ��Ѫ[�����xEhh�?ѡ�$q�f'���3��}V����������U�	�+L{�n��3��i��J�O~
n��7!���'ex�%5t�٦��.t���z�E;��VZ���0�_Iƶ�=m>��������(�Op>�py򇡛�K��Sv̢�����=Q�TҎu�8�ܜ5DĶ�u@� ���1Cz�!�>�� ���g#��&;���h <c+dv��3T��O �9�ꇓ�f]�
�� ot.Cs&i�W:�j�r��eD5�0�͚�uN8�|��I���$�׳1�����r�u�R�0`\��Nq���/�0[�������{Y�I~�V��p9e��豆=�S�+z
��-�]�#@�c���IM��p&Y����+�i��P�(��=�qO�f[O���?�O_^������F�>���̮aK*�kR�/��H�u��#��L1��Z�i�����Ab�?{���X�N|������ϵG�nTď5��&�@E.Uy�8
���dm�4\�����訐T[��Ԭ=��z���5��?]k��Y�0�����F�{'��/!!*n�+~j��ϭ�ȳ��%ݠ%���nH�i��*2�f�Ϲ �COB�������P/���'�p���x=�ׇc�'�q���}x}���H��wE ?6J��IjV��C���#�˺B>��V䗯�(W�`�n��A���r$�{�� J.�*A�/$^e�C5;cլJ�0 w�'�GpbZ�y�Am�.�� ���3���7���e��9���T��da<5{�X�J�S8 ҥke�"fP��.s����ԡ;P,S�h2yF,��s�W�5bP��x�SN"Ð�QH#�:a�D���j�D=zn�$v AoE�$w��T��M��U֊Y1{EJN�Fo�#����G`Lc�tV�k=������j�/Dl,"�3��xsR�!�G&?��=����W�o/�;���R��1��m���~ݪ)���s\���v�z��o�p�CU����H #��e���b��`}rX�g�ٸ�J$[7��D�Zp.��;#�Ø�T���>r��d2���(F���>t��eW���x��~e�z
�y����#���Q1���.8���+�D_�5�����R6˪����Ja�+22Xڦ�P�ܭk���pdnwC ���5����1�ӧ~�%/�91�������A��+4<]�9�_�����u�Oyi���h�|�f��� #M�����g5����e�mf���� �n�D���L�/���D9ea�Ofȿ
��ɚ.L�L诗�)�z(E�-j�j|�����:�<����-�v�k[����u�elc�Q��5���tI��M �I�t4�� ��1b}�X 7n�Ck V�T	�]+�W�*+L9G�P�
O�)A�:0SQ���PK���c���q��!l]���h?�^�O�j�h4��������3GН:̘�VH��b,ރ�KvZ�X�
��d�#�ľ)����A���	�w�~��	>�����'����~���'��ˑo4T�X\�q��s��I�R��@�Bbw.t�3e�P'��Q�݊�-����
�+E�+�\�#���By|Тv�ȝX
��To�[��'�����ߨh��HO�Nt�C���`Q�)2d�<5�=ط2��ϐc�Q��@����n�Y;Gׇ+m^L��L�?������˯�J���j�5�-}���^��$�~���U5a����\�I&����^r�j��ӏ ��
������{u�W�Ю7�a)Or�!�;�cm�A7f3�.(�
�5k��C�b}6�8���Ls@ O�=;�#�<EX/et��[�� �}���d��sU��
.y�uh;.� ���{�ۀ�*/���Y�l#[v�lտ�~=�a�l�v	Y�\�S�	�6&h�;+�xnG&|G�F���L�#rȒ2�����������n�-i��#�o}�z�p6���Q{uX�������l�laT�F]��߿�����ܜ����i��Hti׏7G�6N!_?y��o5˳�殱�X���1�J ��i���=P>�����`dB�۹���`���R�i��g.`0����W-��S|>ػK�Wu�B�4\��Z�ۯ���<��}D���I+oe[m|���B���:K�$h��2<�T�	|��oay�+��[i��=+��ù��p��_e;�Y��9��z�.�뎟la��P���=�;.&J$ƺ.S�`u�I�����_Kȱ.ju���w��X��Y�Sgx�G0ϼɓe�4`�l�j���8�AM����_���J3�Q'���E��q�bKt��PƅD�u�'q�tPv?�D��G_~oQJ5�V��9Z�l�E�I��[�r�_9�!��l�:@��"�*R����uu��&�4�kc��iY^<L`�A�d�z�Q����a6}?�A��nEe�$����0N�8Y����b� �#	���h,ȣ��g�vC�̚�= r9H5�Vf� -aj�� U���K����SI-�Ԇo`21�?��"Q9cx��_���/��`/̿�������}�����.��S��ـX?��RA�2&�|���J>��z�j��-���B٦6���_�ő�����fqȦ��1l7�Z�ZDQ�tPP�Q���-B����ᠠ�0��g��tzlN-_ς�5�;+q-�����nPؤ�Ѯ?]q��]D��˾�E�N��]�K ��<�/�@{�!�4�����]�R��r����n�\ _��@B|5X���a#���@ ��wrO�9X�r�sM'_�VC��e̕a!D:�i�am-�7�L��7ھ�� \5F>�k��VHଆ��?���_c���}���J6��~(|�ex٨���8�̻�<|b��K��� �;Rˮ�l���7���eᑙQ�>�H'�,V���U:�2^� ?��l�oc�H7M;I�`nT̳Ww���U5~�CO�ԍ�^x��jC֎���-�p�lt��瀒�e蜽Q�~��`_�"d���k��,1-L:��ς�Ȁ���Le|����r`D�TY�_!���K�r��Ķ`�1i�y&���k��L[G�U��TcO]X�k�ad3:���=b�>P~x�ӳ0�J��gc�V�}g� w$���%�2�t�5l����V�.���˸���ty�^�`y����<V�>ⷝ&�[�i�?C1�F�*]m� xKUT�7#�o�����0��/D2�9��԰�5 mRgH��^�"9i@>��@��Q���-�w��eZbR$��1�T SޗYHΕE\�rNYp���ڶ ~��cƒ�'H�hn�}
�C���{kZ< ����vK�[���4|�9�ev�Ȋ�M\g�}R���F\��ќ��r���#Ħ��):ɠ�b��Oc(�^N�	�L��+��wf$S�&�����d�r��
Li���x3h��.b��4�~F)��CpJ�͡iP��_���y�q�	���	��:4f�3s���P��(���PX$�E�wy�Y�2�=%~}�'L�Z�(BT�)#
�� ؗ���b�㒤n9��9;�S�N�FJA��[�řN���N�\�����'<���CO/+&�}]@v�߮�N���#�n�,��/�M!٧R���a8�*�ы.�e�>��T���� B_[ЬVC�6~Cl���8�	Q	B\��BHc���-��Tb��ۧ�xT�h�"v�1��2�,3�j�W��J���Q����0>j��'|TX�4Y�<�7#�-�S~���%�1�ƌ��a#��w|���^�F�J�'�U�؍�d:��3�m����#l�9�bۓ/S����.S�P׃_��X�c��!L�u/!��ay��$��R���h� �L�@��+QN�ҶʿBͫ޲�8��s���O�a���w��eƛ�mF���v �ӧ&/3'f�؁Dq2Ϋ�%��ٰWv��JA�b΀��o�h�]r7Ͷ�C|�s5�a��lɃ��5�ـ��7�w��V�b6�c�%�+�8=,Fb��vr�	`˲������6Z�ы�a���4��3��C����h5.�0����Զɖ�X�'f� �c���3G��v)��,+�I!��8�)����QW�%Y�F?3w�*�ٗW2��Fh�o�2�I(�p��;�X������ �`(��4*�SI5Í�����zPĉn�)�ŧGt0t�H1�o�,��g�̬��L�у��Z!��e�����gM�����]w6�h@0P[H���G{����=0m3�⧦&RD�"7 ��"js��kvC�o�m?�]	���І��<�e�zd���z>l�� �S�(� ���_E���OK�v��1�{0T�����������(��ø��HϛkW>��Y$�~�����#nW;��sm�9N�(8��{�P���GФ�ĄC*�C�J�W㈋����v�b%2i�".�[���:P��1���ם����˅;��,�����θ�� K�d
� ��#U�h��D��(V[Ҫ���@�7�=`�~���T���y��"F�ҼS.L���c����1 �Rq��8�G_s'N��q�!�tyT���v����+7�B�ޮ�l+�Po��h�[G�YX���əl�|��t>��G��U�Ӕ�I�&����"��kY;��k��C�&��cј�}��A�#K�j�L������ձ�o\�7� Ł< �>'�ϳ�����PaA,�҃:�]%���3��ӎ٤� �S
�?����	c���m&�WY=lU����Zu�kѪ���:�����f)��sL����R%⊮�B�In�\
�3k3z�=�Aؓv�F\hz�����B8��p#����pr/�Z9�o7mб�TTc�go�g:�8ɏ9�od^�C(��i+p�û7��|�;[SؗK�#i�Yn�scY�dcM�s���3!�bD��ZՊ%OQw�gP�ڶsq TL
�����F�^��캐��a���O������9��Y4�"��;l�G�jԶ���}��-�t� ��ݲitM�T6��o��b����+9g0�`o�r�_]m ٵ2�Oo(���.�{�
i���m�	�c '��Ӂ�\&<J�O7�}CK/���+�i�tQ����z0�����,���]��5��� I&�&�o�����@����{b�R�9CƎx��j69���C)��tɀ� f��l0�(���D/�&��2�1.,��tn����a�>/�G`�}$ܠ� ���\���d�ʐ{����J2b\�t �~����
2Td�g5<�[��פQHT�FH8>��(/��/�p�2�� 9n�^�B���d��V� �\:��G�x2����k�k���xɼ9����H�ƣ��:3t���<L�w�����2,,o,�4˹��-��x�9�O/������Sl��k����I|JM$�}x|�|�K��{ȃ�PX�Bۥ���p��ˏ!i��z_��]T�n.w���0u���O��;v%<���jm�@|���n����1����l��Y��WQ۴܏���&Ϊ݅}��6���������;3a5��F�yN|*~���:��j��^
p�;��
R"X[q���Jd��ErR�V�ͪfzv�X�����)��(fd���,�aR�"��Q����*SH
(�?�C]���Q�3�`�p��:��x�+C<j,C�
��d����W� ���u�C�kk�߼7��e,�Yp)�H��Mo��
�a�%�A����6�o��k5^�]�w���O�Q'��A(,��Sq����=8�^�T�nb���zw�� =u[�6��c�B���c�I~��}�o�i�)N$������"�!��oΒ_�����B(��e���{�[���4��gEA��5�k�m�eF�� H^��� ���v-�q~y�=;�R3�� wfnh�U�7'uk:&6�C�%�=�0���71�������(smI�1�j�jSO�s�T�BdP�����.&�֜d;�Ua�ZB4l���d3��f��ӹ22��@�[l*�����O�3��7��ŦNY:J@���zi�ӷd����������W1p��A�&ʷ�h��?Ep����,AWx��A�P�/�|�!Q�Y6q.@;t+�:;�A��@�s#`sW$�y�s������TV��F�ֱq������	���r:U{����E����N����]����1�=0�r��������;��sk?+ϋ����d�IN[��c��� ���r7%�������b�,������D	{�,��/�D��sLU�;D��F�s�������U
�{'�U�E�&�\Z�>�¤c��<��8���oH���B�2t�7	#Prm�]�\��-���&��oL����-�"�ե��GF��e�ddOb�j��v��Z�����r��bJ����S��Y��c���^�W'8hZ���]���n&�Ȉ��O&���c�x��̢xy��3�q���4�7�9}(�z��h�����S�ߠ��O=pQQE���ycLB�r��FB&ʗ�cs.�h������<)yq��1I�'ȆT8��l�W>'=�}}��JK&H��a�S����s����e�(;/%���eZCǋ��^��H}ssU����<H��B�g�Z�Ne�T��oPզد�����|�Ͳ,k��1��(~M��eRI������C?�7/�[��ŏ:��O�J�8�jn���>]��XV�Ɔ-��u	@<"�4R�v����ʽ�l�{�u������+u9-��ڱI����؏��[p�'M@���������^�<�^1.��;�u��@^���Q /T�F:��2ov��l�|���v�	���i�,IP7���+c�l�+��(Ys(���e��-�`�R�i@fe��O�w�q󰱸h.q��vBl��:QYW=}#�M�Q�|5�uđ�H�B�6�N�c��H�
W����~JŴ�ĺL�8!-@�\��R�B[��'���_�X���.eG��.N�N����fU�Q��a��W�_�g���q�����2��HP��A���p���r���� �r�}%�Ͽ���_H�o%V1��W��È&O�^�!�:DZ�{iCz����I�gN<�D+�Q�C���Ĉ��Nổ�Z/�= �;���ٲ<����w_ߗ��co2v�O}!)o�����>^��`p���?���9F����l0��V-g�>�}�H/���b U/��!�CvM�3�ռ���l�IKg;\p�N	�Nt���4d_O��zKl^������/��C���Dz�<�o��^s�M�
���h���,fy���F�'.����.��E��E��}�%���\:�^Xw6]ؘ�{,��<��Q-@)P
$�y�.(ك\ˣ�r��~ݩ���	��� d� �5q�a�B��e���̧��"$ M�tmqu+S���Z1����^n�(�S���)x:{W�z ��a7n�k�{"��ׁ�������?���T�u/��G�GS�/��\����9V�*>u�
t�UA°�iV��b�>)mZ+9� ��u5�h3�3V����|�6���k�s�|�����i����̨)�_����P�XPUs�j���I����|W��Z��ˊ��aX�����+�;�R����.�5M��봪�<uy�	K��(��L���L�]�F�.��Ƹ�;t�M�����	�B5�O�x������`�,;����h�M8�%���%bP����u��f���ݼI�����Ã�
���ѧ��#�'���G������]�(�*iU?�@�N�t�oڈ�]��ʉ��5�Oo�q�ꡏ�O�������͢Gw���iEV�u��`-���N��p'zO��#���n@ʭ��B���}�q,M	���S��甮=�b(~^1Q%�xO�W%�3o4l�B9����׳�(t��f�Z�-['y@�@� �F���@i��?�"O�1	+�q�H�Ӏ����I���-j�d��N7�D���:�ǣ]��hC���w,VeM�d��(�a
��K$l������
��E���b�E����+f&l�;��yem�+mD���!-e>��tk��lO?�3g\b�wC6��ZUi�Stf �o��=j`F��U�O�(6���LD�fn�� �s�1c�a��1DAu�F�Qe�i>nTwɝ<�)��&/[A�m�;���E
��T���$㪏��|P����%K�?�@�6�'կX�x���y��$|ʿ6�S�3���^d��D����I:?�Tۛ���"䛦&�p��8����@���jA�#�r~���Uxr8�4��.���7w	��& ��� ^S�WBf�3�)�V�&���� �x�[g�!l��p�I�Bm�g�N%�ۖ����0�c�A$!E/�m$-�J�\3����yt�c'08R<�M�E� '��u;9~�ԝYh�ש��C_Ĩhj��K��$���sgQq?΋�	Pn�����*~��T
端6p�m*�f-�Ҟ�}�I=h�)�W��`��Gگ��6.}6�_����� �CM��fpa�*�С��*��-��~+�b(�����̍)Unج�隈v�F�S�>�Kj��`��;KnO�[Q��/~��]�C��n�w��1�B�j�n����B��,���W9�%�8�L��ye)ā��:`�l����:��}�K��$g���� CKj�:�d� ��+	a�[U�TUOsΩ"��(��ۃ��i��9qM#ӤRj�PúǸ�B+饄,���}��yn?p���>�*��yhB���m�h���//̡�64Ƭ��xY/��y����kЇ\v����pH���p<�+�Ҹ�$a�w:�K�=�Pbpc�0��[ЁKr��#�{�i*�eB,&P�Fy�IĲܞ+K�;W�������wlqk��Z)����M��X��B����*�dɏ2x#����g=rP��[n�쑑�H!��o�[jc��,�A�/a�Q���I�K�P���D5Xѱs�A�o�R�qU�!�C�s�l\�5R7'�&���%H�Bl�����귷+�jT��ն��>ũj#2�#��ٯ�Q�����ń�����7��$��ހ��69����\�X�'θ�5���d�۱�l�*&�1�ve>QO�l�yΞ�[CVU�㿳�1E ��?i�]�b���_Y����d+)vU�n3.�W��:�71 &[���~�@+�v���� �@,�t���s����G[��q^��)6c2._7y�j傚��;�^��������� 縉b�#��2�=�}�9�������%2N��i��'��r��1��F/�wx��ZG28��Y�
�����38+
]��~��1ki�/Qt�r��WHx�
�R��*���;>�t�ĥ*�#�}�[�8�[�}��\,e���P�o1|lrK>��[��t�ʑO�k�ք�?;�}���w��h����n6��.��hh34a���Ѱ8�.����b����m��y��^�|$%qL�X���)߳�ۯ��&E����Z7DkL�1�zԯ"�ُ����).��r�tP�2�� #Bכ�ҫ��s�v"e�E�1���L��DLWT��xJzn�m��Dϋ�n��H"��<ר��-C�á��Ƴ�/�w�H�
h�y:/��	������������ nK�*�b�;�^�	���9��J��0f�]�L'A��[�_�,���iR)�#��	)T~^�/��3�-`����`����h�~Cr�<0�����Ӳ����ʀ���?`��(.
�3h7�l�Z�q�W�вrU-{�`��B�#��� x���ʉ�'�Hs#�^A�\�7HO / L�'(�nh�,m��^����i�%o��Ұ��8�W}��P�+��-������F��j��*YQw�_�H��^�t��S��6�,��A2L�-�@|4�/�3T�FW�p,40j������O���i>Qՙ���$��g�C�����0_8�����Zp��d!/����*?U.Z3�mAF�n<���+I�yv{q��Y��î�$�o�c� 8n�VE�����TD����l�T��D�6%TbW�k�ϼ#��{��q��ѰY  ���zn�饅�jO)��W��I!����d{��W���L��H��	��'�T~���p@��b=��w"��z���9�뷞�VBY�ǘ?�E9v�_�@:s�Gܽ���{�������zu!qIwb�n�������÷(�XX�^Z��!��>���[&EFK���ڪa��@M���"����� �|�n�0D������+��ZPM2�|���*Ĥ���L��u1�n�y(��4M�I\�c����!�E����֞���%�N���p=2����h��j�K�ч���_ϒ[���,.z�r��K%+���m�f�El)�+eU�o�|�F�����\��_�儇�������O:�i;���f�a����Wiʂ@��mpy�� 	���CS�4������n����JU��2��o��ن�1����`}:�j@�O+-��ұ>�(���2n=8=`d "�9W��D,a[�@�ʹ7���%�R��';w�7c�AHz����=������hU&�kR7f�ZuU��*R��`x�}΁�Fn������孷�\2�(nv���d�$��W��<��l��ig�4��j��t8lyx�n��a��1�pbK(�N�2I!���ӦHM9r��!���u\gEJ�1��ʍH�0�X	V6/Ŝ�gB�]O��C����?��D�MF��S:#��ݧ<���:BG���AjH���&��CM���r���Ly�:�Ğ�Ki�0'ҳ�!��Y�pk�O@�����@Հİ�� }2�<D��'����\������/���J����vo�-�">���?.�V,9S��'v�vS �i�tNxYp�:�a&w�Ɂ�O�ڍ�I��{��ݭ�-A��wW����f[�YܤtN��P�nI�8���IQ�˵���IUs`2�J�������o�O�f��u����82`.qW����O���L��Ў�n�C�w�>0�!:����D�(�pA� c��G�\R�(�u<��7�[޲Vu=O.+œ7Q�_GQ�䲞=�~�C�����.vE�N�x[���S1��2��l�� l�:�/�.?;5%y�=�
�Д��fC�����r�9��ܤpADF����=�I��N��!	9��ܩm�6��!�=Z��1����OC��X�޿Z�Gt�63���]�Ys��^�Z,�]8W젂������OA����IO�v;7+�mg��{�l�%{o�\��D�3 3����:u�*�=�L���\��d���8�k�<�ܓ�	YxZ?���w4�)T��X��P_�B���W�x^�Cץ���M�?����Bڄ�.~f�|]<�e"������&pl(���G��{���Y�k���4��0������]�fU�{gǑ�r-,2ەrk�o-ަ���}�k����T6�>m�*D�V���@��Y��Ŵ��t�c�_d"�E*�ˮzA+����N2��Nt�1���L~<SWV{�����,�܎������_uUd?��б�c�X��^�\��D���`���­�T��@��N7�
���\� ��Ï�ᤓ���k\e{m��m�߷�9Ӥs��q�^΁�Hwfk�U�`�c���UO=cd3�}sW���[��v���
���)z;�Z���3�
�TH����R(��
`n`�7�3��fR��i�׻i.ݍST���9'�#e�hf�6^�N���!�)j�;0l��u�0Q��}5��W�d^2�9 	���g�ϡ���޺�jU���qil���r�W=i���E]�l�$��Q��Fh!��/R�<ZgS�������.dEn����EFϘm�Ĳ�SL#?L��%��V|�SN��ҽ�d�+�L�rIչ�ƹ �]���s�}�K׵���0����ry$E�Q�m��x�'�Un"��s,N����I�$p00W�0U���#�����"�<���'�T�� 
l/�Q��3]"!o\�xt^3cϑ$%�	ֈ��^4�L�zo��G34Ҳ�O���R�T�e��~HB���҉�A�rYE.��_����R>+���S`��)Z����k����P�7��ö�93�+]�W�y�{i�/�qL�a���QU#	�e1�����)�� 2�F���GQW�B�'c� 
ER@��,dE*�`
��P3����B�*X3$�o��32��/�y#��H��
�%���
�����z�H�1�1&�/ڀ�� ��y9 �:l�H�:�X�Ȉ��U�P��U+z��bO�ܕ%��
q�Ї���5�"�3��ݏ=�O���\V�ˡ���A��������;�g�❊�;-�����	��i>�;r�� ��cHk`	C_ Sl��J��$����h��-�͛>9�`מ�����r�oU+�|q*�>-���Q�kOĄ�p�b���mw�;�rB0�F~�|�d��@��W�;P�$��+}�ddXw�>�V�����3�9E��~;�����c�*s��EO΁�//0] ����ґ=��7p�� z\�]��C�¶�^����Y��R�y�4+�V$�%��_�4}LD����1�i>��e��ܭp�C6s}��R����r���+j��e��myI]��]������s�p��!b ��a��z�qz�k�۔�����Z0��(@a7:E��:()��0~t�l�d�S"V��X2�p��[�KNڇ8r�
}|?ak�˲0ZJ�M9\�ͫTWyPt���㷗B��(���<�B��cD�?̟źCl�����򆐲���K84�m�I��h2�miP���q������j?�x�b9�S���r�Y1�S�P�2f<iȡ��]�7c�8��+n5�$��nBr졓;��8��9�y���]
���0� (��L��c�Q��s�2hA��=N� ��g��(q�o�%���������C��'P�g��� #�5n�����'>�O����_�ٚL.���Y#u�����4���>��;Mj?7n�i!���C�-���b�2�'�N�qZ̪-��p8�/_�d�����E<;X��6sFL��Y6_k�K��r>�������k��9*�]��,`
r|�]�u0�G3��k�F`��(-{g'��|�Vh,���_��Y�W��6�[�U�5Bf�K�=�z�4�iť�8j%��!Ί�~�K^�.����sy. ��qg/�P�8���6�ju���X��¦�0�bZ�MK_����Ԃz�Y%`��e�xI��,)]քLEm�m�C���~�b�ٷN
c���M��6�jHφqj�[*~�Ά�3c���U�ѐ�7SNV�!g�������D��k$��+�ɗE2���C녮�i�L�%>�bp-�ɞ�Ҕ.;] `!��:_�vn�ڦ�I ���\�s�} ��Q�A0Gl�<Z�@��M53��iC���}&xӢ�wWiKJ&y���s[�z7T&k��&�=�����Fcdw���XE/%�t!��c�Z�f�a��(a�Xy�w�N�U�o�#k�Kf+��\x�����3{��0�f,w\�F?Y<uҲE$-0N�5�2�J�?�ME�;�wO]�CD� wZ�m�A|."����zA���@p��76A�(d}:WH���P�^0����X�I~�4Q��w���n�Dh��ḣ.���`7��f�p��X���wh?ͥzTq�sefr��NY#*�Z#�r=߁���nՉ�ݤ�lS�AQ�"\栗�l#�۟�C��t�/J���2t y��L 5A�A�U��L(!B�|r�t�����8������~�7O�$j�X�R�1��P7
c�!lyq�]ª����3������"�E���D�%�l�<#Gxh[�4g�;�1IX�}B�ؐ������[2�a�#�/�N�\Fb��ą/�����y�̘i2fF�AP�ܱ����X��S��������У�<iz��?�0�%�W�5�aM����KzK���'����)D���\�c��8Z���WQ�0{���N�-v2����e��@���s�.�r
Ք6C���|��ac�,�vA>fpc�w��w��lT$M�$2�Z���2��e������U���C�u/�#���D1"�mbf�������6�7X�|pA4���ܑ����׵a�k��>Pwq���*����v<��I_B�!X������c�>��>����N�1��ݔ�U.�����"���@���D��Q��Q%"�ǝ��f{����-[�w}��еiR�a+#�Ի�z�2@��N�uZqI�3f�>.����I�; �!�Ҡ�L�!눆E�ΣD��N!?� dJ����EucPh(�]�����#Ά�q�)��D骗-U"�)����E���֕�K��@�������0y2H����͒�>��Hr6��h���n�6El9m���a�_y1�O: �/e:�*�6��i���%�J�Ĥ1���w`Tȧ	�]UC�S���N���]����%�B��MM�5"���S8�F���5���A �~L������[��ht϶�*p�6E
ď�m��� 5ūUE�44��JL����V�g\k�i� L1G���,�W';�
�)�I]g�b�$��*�M*s {��yS +�~�+���;n��^�j��.�����1D��;wW
m��&N	1�O⃬����'�"���m��pKK��ԙ�JS�b��A�*)���N9���3R���F��H��;3*=�ӕ/�C����B|�ʻB���"}׭�1�B?�l9r�8���J4y/�	�7�~��q�(<��2������o�t��w�)O��(��<L�c�u5!�.�{��ǒ�&;	�.I]��4��a�:�@ˍJ ��^��#�E2�P
%"Z���rh��R(�>�)&b�2�ܲ��`G)�U	�q�$K,l�#�O���.�+���3_Vq���
�]ca��y��hl�:�����<�\�'�:Ը��Q7��rV������6�C���E.�C��Q띧*�`i�u��/ 擩ST�w�ɊH�뗖Fsf�]��U_�g�(��|	5�d��苎I�}�&�s,BY�(�洛���]��L=��я��U����Ȯ:�v�w�z}3���h�P�;C��\>��xzB�\�<��������7���`���Ң�WaXQ ���tQs�'Mwq�P�Q�Ki큈��7 �<�={�C�pk[&�qY<=��� ���H"ḳpAT�����f�O����
����;Tc����s_�F�˟K�n�J7��:s�|;��7)�����>����	ᔁ����X�O�e0m��S�~�F�]҇�c�j�ny��YT)u7�:�T�`0r6=��Q�r;ݮ�o�l#Ӕ&s�x@�u��n)�`�}�̼Б��;6ש��9"	%�?.)�\��o��<�r":���P�no-��0L٭���U��Ŭ�7V8�?�xT�d7���h��pݓ�c̔<7�x�g�ޥ�TA��c��p�,1nZ�s��<��'����7oG�OU{���P�O�k$�m����G�%�>���>Ǵ���TX���ז��w��u�c�F�s,$�:�lX����}UKNl�DϹAj��2$�@�_`��՟�g���5߶Ԑ N�g3�J4 㺩�x%���(Z�ĝ+]Ԯ]jX�q<����"W�b�;N���(J���-eR�܁/���l����9��֛h���nB�AP�j���Eh-[x�[�6�����,���zQ~�o;�rK"�@ZD_v,=���į9{�t�jl�p% �"ԃ�fj_���t�����t�ӻ�~w�&EK�����4K�f�������-b|&$2b��&4�\�����5f��K)�,9��\�o.J"��U��0#7���x��L�|Ͳ8Z@v��rk�~V�?w+4ᇷZh�J��K���! �Qe���-Q�gc�T��<-����o��ꃕ��A��t�>C{z,�hj�	d�tHId����7��%g1�[� �ㄣ�ܺTD��
p	��p�2�5���9Dͦz/b��8��E�f-�����lrr����: yu����[�$L�fFUl�ff���<5R�ד���	��.Nċ:Z����s@���W�N���ک]9�;��.8���XN_&�Fdy���{̊��z�rž��UPz���xL3�_e�d�Ʃ	GEo;�0�5��Z�|E�f�N��J�B6��>�|_3��p�g�Z�c�=�x�����J�q�`�[�����B;��+�L��eX�'�#:���
ͯ�i�;����<�5����U��j+�����cSy�-�Bt�h/�*ӲQ�BJH�V�#�W���<RRS9�:P�����?��E$?��Y�͑�ۉ�cY�F��,i:�9�̅-�8���W�9l$np��� Vt~X��bN����z�O� į_�-l��Q
��i��L�?�W�U]{�Ϧ<��J����Be$aE��j�ӛu�J��bh���$3�By��oQb���Cn��R~�. ��BCtZ��2��0��?G�Tk��|:I��M����K&��B�؄�ʹ��`X���׺�������21�Xb,�׾I\��r��4L�t�0'w�*��~��ш��]�a���ӝV�#P ���MT���ST���[R���'��.8�"�7�8�B}Q����I�N�7ȱ̒��.�n�]��1��P$�Ka��B�k��{&���e����p�sf򸡜�i�(֔����(�emI�'���F����n��A�pk�v]�D������tq��A��͟�:�Z�}<6�̦Ҿ�%�F����k�
l�b��Єoq=��g,�[z��۵�w�C���m�8G�/�-�[�˖��\�-���H��|}r����&�L*�������<w����ʀ@��P5�����êy�m�DBE���ښ9�j�	E
O:
~H$��ΠBP�o�E���Ì�Yo8��`__�����]O`���%ʇ�������g"59�wb���{�GH'��)�.��*M�|�k��7�o��'�y2 �W� ,���;z�����0}���O��e��;vFH2��c��S�%�xYd�g�� �+��t�M��n��V6G�+�<�U�P����薿;���u&B�Q�Ϩ��̩�[�!%gk"��	I/�W�.]�4��H�)5�'ֶ�
T�ʱN�z�*�I�s&k�Ư�l@������f��������؝}
VRB!X(mW$61�ϝ��5hY8�X�:����:�T�d�Jv��y�YtF^c�(q���+���ξ��y��/`M�����Z���󘭵�_�8�w�ؖO��<����Ѐ����O�#��^s�W-�Ϙ�8ޟk����'��=�����k��4���a�W��&xW�{=yG��2G�ֱ!�f�����r�=x�,�ƽ48Bg��t���9���թ�9jC�~�ʟ#�<�85��qZ�2���׀�Kk�O2t��m�N�:�o��.|���D;��~*�`]/��V�C����X��_�JԿ[�t.4ZR��`{:���I����ܸl=r�Ӟ4�MO�\�8�u�q��r 2�"6`3X�7(����7N��iS	rv�n�
�S���.�A��/���z�(�E��"��*��=6LUz�Q����nr�C����֯��xp�Oe2�������m(�7{���CULe.�v덷�]0�|%9�4,��U���|�����7��[n�|zf@�/I��)��K����MT@V#��S�aK}&�� ��v��\,T��7nM��,���mF�?NC;U�����S\������)�m�Њ^�O�-T��վ6֣ǋ��Q
)��H�����H]�Qm`,>\Z+&�AH!��ާ,|�`���rc-+�/T�%#���V��8����r��u��e��?n��G�Z�k&M���Hւ��4�$JR���/��|�И�o��aĴ�}�;��Y�M�E������9*��m;��^�QC�8��)|���1�a������C�	�7J� ���!Ę����WY[��y`~���/�z	�:���5.ԇ�`�=]n"�>��ѳ���� ���9�'��sIF�&��*�n�l�}�"л�)��φD�=S>��7S�A��Z�!�����z�d��7�s�R+ԡ�����cF��F㹋S��q�2�In�BDTC�L
Nt����wYO�	)D����"�9oȽEs�!K�	���c�����Q_�8�-���X?��D-.j'ēa��45�odYKe"<�;�`���$QA��]�)]D1Y�?�y��KzQf �}��+[�INߨ`��zX���+3��n �k���5~<�B���f7��W�Jl� �?�;U��1Z�{\S��p(j�-���*�ޝ=�+�g)�dz��«���*J�@�bQ4;X��8Ѥ�&�V㥼c���vl���^�*�(���1 {[���Ѩ��K^de|j�h����ti�j���s�I�>]�pw���Ӟ~`��:��~:���l4��D���0�%��9e�$�gtBW�N)��w��;�7A�u�����pS8{�lI�τ�Tn�|`*��Z�w+�̤�Լ&�FحrP~K�����W���}TW�*ʸԖd�<%�Y��V9�x��"k˒(E�V�=�z�݆�A$ӵW.~(x���,%�8_T��<:/$��*¹i���u|��i�@�N��Kb���K���)N�i ��?�g�7��sIS9{luRh�:kte����*E�q�k��nl�y�P�S�Ii� - ���yZ��H�N�ħ�ۀ1�j�[s���S���� ��Q��2߸��WC3O�D2����<�8+���c����޺ �S�����ٜ�cE�o�5��S)������oʁ��#�;���W�*٪@�E�e�85w���-��j���ҫ�H�L�v�u������X<D�L+����}jf��:�,�d@V4x� �?n.N	Ga*�.-�&1t�ȨȈd��rm��lOBqW�!�&����B�^z?��}�`8����#Х�@��Fjs&���mtn[W�9�hB���C$ݙ�X���-S���{�6+����Y�AS��E6���i�`g���Cswoa�ࠢY�'�
���^l�ٱ���B,,E�G��$D~�6v��Ox?+�";4h�o�t��� l�}�k�!�m	Ĩ䒩�M��d,�
{r�ٰnGc��o��o�X�����Ay�����tV�d���Kv/��z���7G���f���98m��Z�k�|�a_!b6�0��ُxu��ɻ#XV�z�䶈�R���]dwo/�k3��������O��犨Sv��7uBvV-6Hl�w��(}2��IO��)�+\y(_P�f , ���Ay�CIK"���H���b���r�+�*@7ȩ�^�"C�
T��ED�Y�e� RD�s"��>�Յ�ޞ����W#m/�(��'B�d�YM~Bb��>hm��i����#G��B�y��I�!�]�yCl��N[��v�r���*s�4 �9��s��u��Rx5О�;o��ԥw3\�h��r����ԍP��h*dG���.p��G����j���m%I��J�ѷ��_�YM�4�Y���Y\i�uմ���q����𚡠������w)���s�EcVu����%Д�4����{?���3G�4�GV�3�wC�¥��듬�x��3ȬJ���k!��p��8K�h�B��GT��n�hEg��DO:�T���	�<�Ś����l�9�rj�1��W5����g��16Q��趈j�</U%<����6��rW:f�u+O�|81�K��04W�;c�n��/���tb�
Rߡ��nl�t�%�[��x����[��4
��$ �����$�eFδ4�"	�SN�*�ԣ��00�g�D���)1Y�Mw���j���b]�E?�h�d>���;�/b��z��L�|̘Bo(��h� �pmn%$���o�N2[bsDr�Ԑ���p�}=xY�02����˾�ZϾ�S�ߕ�e(C]|/� �q������� '�w��ꮈb��������)p�0�6lدf�0���J�T�do����&>�_��J�8<.=jc}�����*e�W�֢�>a�m��JͰ���,@-o3��<S�Xo���oZ��ِ���g�sL=�G-J71�E�����=���?��'F�>�;��ު+��G�����wt6����[p�n\�5nUk4��n��r�cE���i(�c��Pwq����C�-օ ܓՐ��^Bk��a_�ˇر$V? Ҕ�dY5Π}�]'���h]w?(�e�#$�8`�5��p���uF��uv��
{M�r��!@RCi��.���ͬ(���Ѡ��ӌ�@X��9%�)�"�Dj�;9���<� ��r�^.��{,�U�QFz�?�F)�(���R$����GH=�
nP�Oɟo=�zcCJ��r�J0Q��Lb}GTިXTN�"�C6�f�}��K���;�r�#99m��5��3a~��E�^K�>� D�k�������	��pU!��<�VE��9�(W��4������@q���(�Jy6ǰ���d��
B��-E��ߜ�51		�����{r�3[y��t�rG�bwԉ#mgj[B�������mC�B��{�iᔤR�1!�1���BHNw�H�;�����B��,	͹h�C��
�<r9C��o���i�P-?+a;?�a�(K)���l�/�<��r>��$~d9bSu��ʗ�/��zP�>?~B��	\
�L�($��-��R�	*'��'��Pp�</�Ҥbǟ鱈��!"P���Ezh�L�?�q�yR�-6"|F	Gep Zt�'aV�����P�I �e���-�u��V�]!L cc�����-gЙ�hN>,NSo�(�4��`�aZL�RsF��
����w#<�\-�Ru�IĄ	.�
�A�����H�Q���i��7�܏����|g��q���e��?0�[�=KWT�!����x\j�QƘ�hxsQT���;�`~ʗz�f�$,�y�u*�����{hQe�&L'�uBז�״�����=+�kE?��Ԛ��d�������O�F��3�^�l[[��l�,���sX*�.�(�=y�7-�37��J'�w��/���[rh�.oŪDv gk(�`���!&
=��}E� 6w�tMؙ�����2ܦU�洰�I��%�>m�Dx��-��QCr��6JZ�_��>od'ՌNCO�"�N��.;S�H��cf�fk���P�XBy~\�9����4�YroZu������U��1�>�Swj�fa�y���������Z|�f!�]ݷK�7T��d�4%R��5)40F'�cq�a�R!U�)Ŀi�.� W�O�ɼ}�n�(Y�W�XR���iZy��H�����6:�"��qy�La�x�"2�����h:��a�h��<,k�P�����}\����ě�����\z�����</�T���Ҏ$L��"������r���2��+Am�1E���P�d�W�{�k9����"t��G58W�SX�%�S�,q>���yA���>Og�O�c8�~,&�&���� k���>�/�}��|c,�)9PP�B���]�秃����9��L��m� �K�r�)FD����E���<@�+1�r��{m��H���Z�o�k�ͬ���N�\�鬹&P�@��&ӷ�g �/��]�]�>d�t�D��@5���|tӘ(�i]G�L1TQ�C%-e?�9E�fW�� ��Ns*�����4?ۂ���@�U��v�4o�KunZ�w�)F���l��_�I�~3˃�s�I��,s��0���O9F�[�	~��mƅ
��q�Sw�䥊�iR*b՗Ϗ�S�${rgͳMy^x�!9���9ˇ^��S�� ,�?��.զ��.���q[������jF>lZ\8�
���:�c��JV��W�Zov~SXޡ�g�C���M�,�9h0gw�:E��e瘉�.�s�����@����A�7�T��׆����S�«�ٶ��(����n�}	xH�A0���?]R/�#�T��u�A�|�h���I���VX1�����ܐ��6���ю((�4k��]j�QQƟFQ:Ј7�ˣ���֣���гҒ�,`�*�k#�p{<
�i������aw��uݸG���6��	�ڇh9ة�l�yjM~{�����A+N7Y�V���6{�J�h.N�0�6ō@�x@CQ�x\i^-���iX�m�'�uy��3)�!���g>yv���X��A��j3���t V�δ�Äe:����EL� bpy���U}R-s����h^:ʥ�9���M�|ƃ��H�5y�=�J�����R8>x�Y�E�"��D(��)0{�N����H<�)K��h��ZT{�j��u�0�٤����59p��`�˶�w�5A��[���D���\��1��9Qb�̈&+��x
��z��hE�g>?�=/M��J5y�Ӹ���v�q�h��\bG�v���ҁ$�� �L4G�dS��&3�A���%QI�ch��#.w73�%ĕ��A�_���Q}��� ���Qz Pm�#y3�����v�v4�� \��&#�O{D#�γ�L���1���4�E�U��*\��Hߢ��K�Ym?�J������$
�&L��=W*}�>1��wV�]�*��"uI��T��:e�6%� ��P�"N�L�k6Ik�!%�DE �����U��Ꮐ����AH�L�t}��)��w��ppYʐZu�!�+Hs|�2�V��J����Wb�Ru�G1j��%� ��J�sj�o���^�w���&�i���! X��Q�qW��@򔭪���~=��� P���M-���n���WH�e���-��:�����y�5��9I�V���i��>F`��F���9��ヹ #����

�0J�f�� ,���t�М����"og�U����,t+��:/ѥ��IOV�V�j�����w��yO����eB6�Z��mq!|���WBMz?7���f, ��'��n�}����`���O���l׮����U�K��リ�X�ê�}Z����9g�4x��Q~�U�%��k�I�������#��>�����@��=lH���+��=���i��E ���n�縙�l�i�4��%e�&�[}��o�0V��ޜӖ��p6$}�����#�U6���won"���T�,���r�<J7��7e$��su�μ�7|>�@�]Y�K�6�x^a�Y�#(�-;���O�`���q��XXD�>�us�mwy<��j��~������t���튈�4WhD��b"���;"����T'p�{s���I��^*�P��iTf�*2 ��$@$"�)=�5R.ʖj͝����1���y����� "�A0u��GO�'Y���E��+�e#��o��5�� BXC�V5��K���[,��G�9�4"�Ɲ�
���
�YD�������8��^�#�LAľ������@H֋��� �&��wQ�c� nN]�U�XZz��S�tfx�$*��$}�Jz��_����W@��1��UU �}��D������b�ՆK�*�d��}9��ە9Y��^GHzs�s�r�0��I�.�@�S��e�����?w9�^ ǩoU�`��s���ڏk���=o*%W�է˦��E��mE�I
�� �d[٣�fs"��J����XW��*j]R��N��<��JFf�ַY�r�;X�w�s	0n�y���!�gVM�k�V27@��cWk�ԈBZ��Y�