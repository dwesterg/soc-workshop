��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bdj#E�]�����Ʒb,v�/��L��AQDG�u̝�Jձ��>!;Xמ�?��A��hOM� E݌꜁�4@�7�	dw������-�<�P0���(���\W�^�{u���Zm���Z��a�Do�2&�D{_��lt�-��zV�Bf��74��uy!��m��9/����}!e��etj�l[Xn�Y�����g,L��R�w;�/�Z{\�*�X)mļ�~�r�T�ä�ޘE��"��[�U���Z~
*6����))���A�M
¡ԏ\#ZfQ���;5r�cM^&��C(�^�w�"�=9���JP�����ڿ~Q��g�{h�6��H~*7��T�*�	����}����[?H�fa��s+҈�t4��K�|żD�����ڋ7ە��:�TZ��=='����S9�7��=ᐥ��J�H��@�!
���I¿�";��^Pȋ<�+nZ�O�*�Hi����Nȓ­a�wY��೨��&��+��I�Ⰺl�� f.Ow8L�5x|����NX{���"�|r�<�d�,ps�/�y�`׊MF�Mp�� �nq���,��/��֨^1p��*rHL�DtT{��Y�'1�j���J�(��zpxL���o�,ė(�W]��..Ea��	��V:Ӊg-Ń��V~�,Z�>��OM�-*"���b�w��1~���@6n��;GaF<R���+��@�}G��Rb�+��g��i�m9���=;Э-7aӹ�98' �ϰ7�A�P�`�e/a�8�_^����'��*�mpF��U�������d�GojQm���曗iP��+�C吏o�E�S�b���/�`���D�y�Lz�o;�٣����H �b�n����=h�����
�A�Y����ykGMV�b��f��6gwuqL��p������F����������+��t�]a:��H��~�B] �5ұq��� e��O���ol�� ����-K��.���WX��=I>�]C�
�7��~7�6@M�:lc�j������?��BcY�E�W�I�q��p����(��.L|�$��ᐕFj!�8��k����b0���y�����'�r��нc��8��DY�.Sz/��P^'emV|i���K��xv� ݠ��H���aJk0$�7`*IqH�[��Tu(@`·˱Jk�ۦ��'U�2�:��F���ʆv򺦂��O��LK��]n?��҈n1�^�ڌ�DPkH�%ƀto�d��B6����E��a ��e�����!V�G�"?��R)@�]�xPU_���[��w�����s�_<�c��/������@X�׃iY,�GI�n%�� �W���#s��%Ά¸בa��w�?y����}�!�cg+%&�P6���mR�"OF���vIoIi7R$� Xˏas�T7������tb@^�d���b����(݁����0���Ɍ���|�@�f6��)�V�����.V��I�,~� ���l`�?��Xg��|�-l�s�r����%q����7��T�k4�1l�46-��;;���#��wBoȽ�{'_�e�����J�Y��қ�H��E���.� �F�i�ó㰢!�����޴�3�Φ���-b� �)�Hsa�!�t=�FH7��)PS��⎚�)E1t{8�:`dԹ���U��'�s�^ʋn9�"y�;��n���Z�?#�t�.8\�N����CaĉZ��
�v�[���pY�� <��5���8�#V�T�Y�.�����@o<��s�� !�u��hN��E$�b;܃���1�m|N~�̏S��P��w�^��Ia�Yy�-/�/����!U�����,��6�7Ξ@Q���P�/B�.��;�M�-}�2ف�0�
�h�ňK���C���F��1$�4�4\9�@�`Ub`�ɴ� ���#�]VTXu�m�a�������D��Q���o]'ѕߐ\�G�,��q8���1E���hzN��7��q�/��U�����+�O%j�3��LW7CxT��
�s�L8Q�;�p>�6%	�	f{�
�od3�����F�Cw,�i���D�T�n��~P����@�bR^�|��T�1�Nw=��@��1�f�C�G$i�|��-b&aeK�����m\gTTHs���Z�B�+��G��Q�̑)�
����-��J9�ݙ�[=�u~d�����hːC��n�q���T߆�Sv3K���x"$89��[t���ˇ��OՑ�xp�OT��y4�Yw�)�Y�a̭�?٥�(�:W��<�_�PzMɪDS�E|��b�j�8g�?��t�	f�)Rߝ�����1,��7A�$�~���m����/�A��'�_�Zp���N6��2�[��G��<�y����w���ʡf���K�Y���E0T����i缣jYnj6����rQ������3��$������������?��|Ѻz�~�+B�:�`�z_k��0Nz��:#`j_�'ʄ����@�mY��q$�I���F�S���X,h��e�ߺ��ϝ��w����@|��}h�S�UvW�Pd���^��3c�9��tl�,B���Ԝy�zYZ����BY��e�H1a5�F�z�����3�ǉ�_�apȿ-W0�xHY�4u3��ȱA�|���.���Io(��'�J��6�K��1����3��@q�Ž�K���?�LU���^ݒo���[���K�1�������L�]r$�H�B��E8J�|�-	�������c�W���̤ݸ{lk���ѻ'A����D�~T�21���?�����[����%�n�7����4gAΝ~�U4j�d`X�������):�׹�)ai'7�@ݶ�-O0,�j�#�L���/k<yG<���S��ޭȳ���{��#��?�/Bڱu@;����oLO#�h�C��T�� Rj�I�*{��r�Z�F��T��h�-�l�#�<��{L�Y�v&��A�e'S>5�'�25��V�`̠CQ�`��h~���צRa����E�P����{���G�Q+K��:=Jn$ɾ�y�K�+�`�3��G#\-O��,�6���O�~���9~)�r�MK-�u���^k�ol���I��O����~8�C�ݡ�Xx\� �"���sBKh��p��uTw�To�ә[�@ȼ�����	�g5l�K�6��y*�|��M�l�~�нz��w�o��y'hwJ�}�%�ؼ�-؊Y?2
P���b;������c�H�:b$�f ��mybG�����%q������������H}78�i���l�d���dD��˫��u_�hg�%E h��4�f���k-��5�����k��T���IȺ=�{
���ӧ�a~1�,>vg�"f5��ME�3�U��K�R�ʒfx��y���1R���.�1�qU���׶f�&#��A�8�3�R��-�}HyRZ�m���y��c̰����d���L���UC��2]�2�<�1��زJ����8T8K#�)I�!��&��8*�����!2�}B��|O-QU#~��4����ٮ�U����!��'�f1�����c|દ��j(p���)�>Ae�.�Y_Z�4�8����sD3��Ǳ���s�gT ����$P0}޲�1��A�6�˗xab�Npa�@N�
Ū���Z�h-���?r���v?�e�ؗ�R�*%E}�y���mNu m�IQu@�������{�q\�mf��Aݴ ���U �k�� ?{7B�e��I�x%�Юs-�G*�l��/���h�yA��j�-K��C.��3\��xWw��+0�;FQ; � �0�0��y�#΅�Is)��V}Z����8��⩎7Vjx��\�M�xT��:����MٳMq��L��Xl&_k�0�P��=%�Һp}���ۛC}��W��o��e�awN塬}�Ab Gm�Cy���~l}�ZG�߽��ZRlR��lO�#(+6�MLI�!��r9d�H��Yeq��(��VReUWK�f �ǣ0*�{�pO	" �P8x�CN�-�L-�	@��\u�5� n�?:�AJ�N^M��E���>9�㳢�K�w�Av҆�f ��%d��n@�6�T$�������1��'��*�'�����c�NY=LJ ^�YY`=29���KY(DR�d�(��T�2O��Ux�b��No�y��/���e먜=z�<@d�E�+�W����B�
����-9$(U����KV��d4Xf��PŬ��j��w:*��$�[���ǘ6�.=�w�G��� �Q��u,�~�⥂�_�RM���-Mی��&�+&�Z[k��Wg?7(���?]o>Ǭr�B��s3�hN���(���D��>W�2��#��� �j
ʠv)!���	Nv y)����ͱ]	���F�俤ϸ���<�F�>���LA�M�ĉ:z�W���!(3�ma�~��L��;<z�hO;�0IgΎ	uz4R�ڍS����x����)°
��X,�&�z�ϼ;�6 �^[q@�pL`-���N�n����_����ܰ��H-�e�7��{�͘!�����q���캳�ծ���.L+�Fsb�n�!]\J�V��(�H�$l�n�)�VX?8t�o�Zf@�x䢬���� ��x���)�7򦆾#V>��O�5��~���N���Y�MI:��[����L�Z�`�����T��Q�A���R�JI����q��$����~8g[��V���-Y�»���O���C7�pJ�浃�t@x\����x�����~!�v|�B`��+���Pєד"3��^��UN� {�߅�(�����˰���ࣆ��F�dNpa]�)���k]����}�L$��<�wA�ͽ�#T���l.R �b�Qo��yWo�W 
�J���$%�b"
!ω��JV�n$��wv#g��#�% ?��bD�
�q�d?��: ~_��ĮmX^�y^���i����<��@�i��q��<�EQ��_귐e|��[�GK�MN+��0x�2���s���4�C�$2�"s���e���^i,�Fv��w@)Ɲ��y&
U�UP�]P�&�9���9i�6�＞	�J�&��5Ż�����-C��C��d��+�� ˒b�K�p�������Y��)]�,�֘eX���,D�gk��K�}{�h�F�|{�gDJ��߉qJ��b �3�s0�p9�)�nCW&��G�vP͒�}S���XtsF�����N�ݫ�K����*�,��G�R+L�M
��]��K@΁�!ݡ�t��F��,�a��-����2ǌ05l�>��v��PϐaNXv��G�eY$cDy��$G$��POB���� �.��xՒ��mg�י^6����F���9[u�a8��"Ϫܩ!��Q=l&�q��3t���`5'�5Ѿ�.5�?�#2���Kh�ezFV����װ)��XQ3<J�ACJ@�E�/�ש[�~�K����kʕo�������E���ε>Ƌ�un��|����t�,�����F��o��|��}!�����K�x���^��{}�p���p&M�G�����{�!yQ,j��%Q�6�W�-Wg-�MJX�Ǩs������~t�ʹN�*(-�[#Ï�*P�����μ^zCH�n��_Oza�Ug�S���k����Fi��l*]0p��T�=e"4�e�*I���ܾ��>$%�]/C{��@V�@���.�V���[|'��+ˉ$���f��N}����g��Nx$�ŏܲ+/�nmf�'�@]B.HvxʳN�O�v鴴�3U���rk����[�(
I��m�(PAA�?H-	`���	�n�o��4�e� l������u.��v[���Nl���)�^��E>X����^{5����	sl�i�ȷS'��Q�G6��.�L�qc}�9.�~ɗFʸ�NPZZ�@N�{�Z�o�h�������@��Z��4_ ����|
/k��1:�uE�r�醴~\n�;��:L���+X�������oq�u�K��XA�[u�<J��WDw�2�N+��䷨�������B� -�b]�<TVO6�m,pCI�҅<<����T��-SA�Z\�#3�k0cV���Pnanڐ1񇝴�ʒa��s@~�D�G��/|s}�&�����D��_�}��_y��8Z������= Q��p2��>c�aX�Eշ�Ꮃ"��U���1�b����^+�ܪ���n� -'��]��RK�T�G��Ѯ�~�o6�m�M�&��z��^�Vz�EI���=��:��廭�X �m�!ܧ�:�2���x��[�Rꆦ� �5�1��º���Z����K�@*6I��F?�DN��}�}�17,�he�զdO��/l�	�r,m�?���yRZ�����vPH=s�Q.��s����[s4;_C��% ����0������/�� ��#
N�*��l���-����.����^p������o��J+��l�ψ��(�8�K��r�A�n���y�=,;OE|� �->>�'$d�^oݵ�EÈb6���/S>'d�B�x�^�)s�MOYI:E�:�c��<_�q�P��'/f~5���*/�ϜS�OoRY�e����N|��^(AG��˯n/zx�F޲�U�w��I��dh��k]R� sT�)�(�|�4�J!�M�ǵ�n�s�us�<��5g�6���k[�8��c�
�Xroh��*"�Ԛ�&�R�2܋���USK?����-qT�Q�aĄ�9��'ma$q�WP0̮�	B7��a�2�J�I�,��y6v׶b4�3�+g1A
V��|53�Xݡ*��A�%��$<�F�GGЬX#��m�c7�!�� I��&q3��c!�%�=�U�G�l�@š��ե�1++��q��\��J��$ʘ��.�J>�[�x���FM_U�	b�f�����'c���N���W�"�)�=���
�!�x�Ȗ�\�.?(��!�E�w�*/+Vu�#�$޶��o�Ų���A�ˁ��l�Y��M�6ϡĨ���i�*]+SZ���C��Z����o?�X#���
�-A�X�[���J�s֗a
���I*�~}�����_sÄ<��@�H���T��H���\R����[ �s��FC��T�l)�˕L�T��	s,[��f���j ��/M��i�\t�ޣ4X;a�2���R�f6I�������˨ �O	I��X����!SK9R-���	c�I͉�H�TC��vfC�ia�I�-h8_F�I{���4K��/�+C��v�I f9��3"�s!�c`��g��,��� �h�(��~��X���G1�/Q� KY�4}G� @��]�t��/���*�h�lم�XKy�Ո�ΪW�R1Н9�4�]�BZ!����:͉��т�@\�N�F��d:�
�3s!�R�ݲS�L����w��5DAo��e6sY$,����ni,�~Xh1�T�Vq���x�H���*��W�P=��2�;�Gâ��lg���5|�ռ�fBSv[�B���S�}L{Q�
��8B�V���(�_�����-EޕQ���s4é��=�^W��,A���%G�hw4�eJ^�a�Z�7��"�	w�u��� h�}	�A�鷯s`�������J�N@(�.j\����|�y
yn��'��.�$�.����� �|E�	,�>!n�Rp����c3N@&�CU��� `�z�>�w�4���� ���,Bd�JȶU���I3G��!)F3�Vsv�7 �['TTi���I���cc�qk�/�!�J"o�f�O��7�c��l�+԰uÝP�5��U1��\[�d��T(5��~ē3Ք� ��飪�� K�8�/=U�;��x'��[`�'}W�V^��,ЧEh�dC8$*i��^C�p���_�E����b��R���df���>qRK{4#�X���0��70�/���Yi��ˢ@�P�\���Ơ��U'�b��pu,�V�25�F���mDڝ�<��k�җ��(���U͐οLy	j��	�C�tS@1�0�|��T����N!�J9Ea�~��)յH��+�N��=,���H��۳���q��W��Ƒ�ZO���!t�&�`UVa�"�ld���[m�M|l��r�]��jWWn�TβL�@�S�28�ME�ït�h]L�ؓ���vDe�`���0`���:�$�ښ]g�,��u~�^	�U>�䓡�"A�')T�gW�s�.1�;l9p�h�U���/����X�`)�a��Q@�ҹ8t!�-�\��
pk��|A�ZB��̴A��+9���z{�E�Sg{�M��R�x�pD��Iɖ�2�P|�M-SY)���u�7����8_%�,B`[���T(��3/�`l>��{���}T֢��{0�FкJ9�Z2�:.5 ��a���Js��:�i@f�^�Now(i��e���*'@�kZ������*A|�"ٷ�A��*!��Ie2_|�<�3N�ݖ0G��w3�nb!�xgU�!옣���bw�מ8�b8�%���B�	F��tS�~��_��6D㨱�l��y"{��D،��ۂ�0��o�lkn�d�ߔqw�秝��S$ظpo���́���˾4g��о\��#��a�Z�\��87Aĺ��զ9O^S����&�e{|�@�l~/G)�CM�̘��0�Qu���W ��)��Yx_<:�S+,"FJ�`���:�~L(�
a&�\�>#{�^��LԊ�K{�e�u!�JA�C��v��!v�9���2�A=,�k60n���;/
�AC&��0���V�i��'t�_�n	6���C��v�+�	�vR���rF��#�xۊ-R���	��M/���
����y�[�)|Ѭ��-���ag��m1�/LޖL��;�%��=\b�7)U��n�O��j��y=��6;�$���5n#Y9��e<�Z�g;`w�k�8aD�����CUyc˫qZv��1�[��>��(Z�<�2.pD�m��cO�S7'��Ҿ^w�Ҽ`ew�_�]w8ϛ����9��꓊���T��VÉ�Sj���������mS�/��E��+6BV�`#�ZO��-��'$��d]q�q~^d^�2!Qq���m�P�,��4����_	U��=��#�X��:�8ؓ�b�?���N���!�)*�e
I�D��`��F��k�9��)�����ڝ$ٚ�,�<1���.��q �z��J���	#V��u**�CZcNc�ѫ͜���we�^;����Ϛ�$�*�����+8p��ֺA��Dd����^ͫ;^�*���9z���J�U��bl�x�`�M��YWM,t�:v}��C�EXR_��{�CT�*ɖ�z? c��r�*�;�� *��{�P�9�Q	k��ӫs��)�+wD/X�.$�P,�$�G��%�R���Y�.Q����9�Cz���x(�8~KuQ��@������'5#�Y3��v��5�v��^=E!���k��:(���L��Y͹����F�F�`�kU�a,,&�����ld�(���B���Hc���N����v�R����{&�ב�V4Oҵ*�̙$5iK���͔�y8� �#l�`lː"�p�2�$!��9b|��ѓn����� �l#l��qPV_���x�fF/kK���̭h]�Fl������Go�12_B$w��*�/���qT����b�B�k���YTN5���EQZ-KS?XE��X�du�E��(u���g�ܙ��z�T �V���'� �\�%�;d�8�gn���#��}����f�8�(I�)�S!
f����+sN��5%�UP�L�M0mG��U�P�e\�O�mr�fܔ@�FTOQWG�����?���댬��FrWD,�V���9��%� ��53����1Q4�2;�E&�pH��0�A׌�h�{(��fwQƂ'D¹��K*��'L��tQSdѐr��9J�-a�{w�=�]���?U�/�k��jf�R�;��S��H��������*4%HUٌ��P>FǑZ�[K��_�?iB���1l�/��A�C����Zt�(	
q�;g�֛b����n8MB"��-:��Z`�{eLD�^�k��r���UO��tx%���ZT9e�ǅ�-�0l���a�@za��w�Z] �x�W�q����/}q�`/ۑ�{A��zoz���l|�3}7�0F����%ӿӖ��7��q6����T��fUR�W?'/|�x��@�-ZkN��!���"vIz���:��9�O2�G�'1>�67��Q<͌o����5��p�hp��܎������ =y�^6}J#s�I.YFKS)\��tMɌ��M��v��;�0����7��<����Y#f&���t��aL��A�{�g�
�ތ|��>(:q0=�JAբ?ƊNkrp�\�j�;�Q�<5N�,W����O)lo��"�|�C f��{pʏ�1Y�ƀ{�œ-���p�������3�(8�p�!���j�)mk����Pw��b�<���K�|�tۺ��}=܌#����`��}-ߛ
�Qز>����Gv�ب��E����
*PK�[ꘊHV�#��jv��BG��y�-�˝��V�f�U�-�n�y㚏j��[��8i��<��a!���Z�$o6�fC�)�d"Īl��i`�ҽ%@�a��mJE4�vMxV�wί��������h,�xxr0����SJ�����f�K4�{GmI�O�z��S>�����_��M,n�;������1�1ɨ~K�>�0X}�q�s�+oCB�\���Ρ�{��1�8��a](cRp�����జ0�����<�h���l.)�g f��VΩl�Z��c=Ƿ����%���v�&o��(>��[ xZ��z8/x���ݡ��~��?���K�jY�p����bǉh,�T�q{"�y68����m ���#&{y�s��{�x���k���vXP�rh'�R��N?�!E8
��WNH��H���Pk�;�xѝ ��9��>ɤ��oC4�D�Cn$����x�1?=�ag����)����|(�ur�-�"7��� \ ��苧�PI��R29o�u}��]� �0��h�C��E�6������c?hJ�֑!��=yheR0>��
6��KB�eshV�`�N�]���M��ਊ|tU��5��e�~�IKG�"���s���߈���2 ����Ag�.iXF��"2��c�|���wh7��`�2�f-�H�_sWbja�%h�{4��¯1H�䳶�=6	��I��Z��/hŋ��@����M�Zf�p�?��a,/nė&ՑGP�i�����"�+�m�o�������*�ԛ`��&W͜�1ߩ��^鷍���<�ʿ���(��z����Q��M"�����av&$�ͤ��m��MO|W���*w��Hk+�Si�m���.B��� w:r�����*'a�er(/(�Fs!�*˷cj+%�)���V*���&�^���)UJPqr@v����Ȯ�"��mV6���JW)�^.q���n�hoަ�OϜ�a)���Ԫ��
���d�*sb��ɑo;n�1X��D�h�xU�֖j���I���=�(f��ԩi1`,/��5�㺹BǊ@��1�q��Z�y �E	e�n97`E����K����A���ޯ���]�F��[p��X��D!����Ҝ½z�|��j��컅��sn�<Bf�1mtW�A�n�H�B�Tt;OL��}�5<V�XإA?��Ջ�P�����_�zs�/-A2��<��;��_���k��-�0n��<a�����qJm���^�+�j� �Xa$�1`9![���I�+L�y�ay�l��}98lF� �{H�rIA1GA��4]@�E_{�������Y�2q���f���8���?�w��gF��ܛ�P� �Y��sBx�D�]yM	�*���o�<4s|��̊ y�kF�� �l��g$�>�b�+�&R�K���Թ�/v�dtj܇_��6��fZ���V)��vV������ȟ}�T� .�r[l���}yM����H�C�F9�&��H�5�ߋ=by1"2;�]b f������r�)RS�?v��>8����� Z��B;Sչ�l;ɾt�W�F�E�-?�*��8�,�T<;9�Mg�?@�/Y��MQh�@8	�R��J�k��C{�cL��@旟�aJ�^X�y���H�
�?�Q��m�*k�4B�6c�Pcꮢ��jS�k��`[��Y���N�C�Kb1�jqbk�꛵�C^����9��ٷ�ܶ�]'�	��`��_(`���J�>E�Q8ݵZ��Ƌ������!" e�� �<��56p��2|=2�Z����L�9���EٮAXaVAm�f��,2�׆�c��Z{�U���vڦ���g�l1��#���{�����=^�F��;��RH)ĩ��b�3`3c��&桃^����#�;< �:�E^ՂMA8���PA��+YZ�X�۵��;�����J�p䈿OlR�,pN�+
�Ը����?-�-F�7L ꘞ���t�b ����+Y�ޓ�	��̓v���PG~���u�cx_��}h׌֪�汰֩�aGH3	�Ů��:��lЋ=�ɪ�#"BKW\s`uF?:�q��k�������.��>�np�~��"�]q�7�m�1L"�( 96E�.xNn[����HK䙔�\{f�>y2��[c��}��ܺW�����S��R�MA> �{�����m�(���gW{	�g�Y��fhU���3���X���!M8� �-HCu�2�v0�@�`�֗�gr9ڎ¤,�P}�T��x�_��3�y�z���Tvփ��"y��]li�4�p{��_�-%F"mso��e�1��G_�B�h>��O���d�R
��Sƴ'5�7_ff�!e���C�G�wd��]8��a&6m���H��t�u�� ��8ͻ#������og�Ld�D��vL���,�P��9(m��ٗ�@+��Sֱ�ˇ�ql���Z����a�N/	c�m��GA�^��FW��ءt�����6���/n"�����O�Z��1��PíN,Z��b,!8~q<;+�鑨�-��T_o׹���gЄ��u�C-oZ0{��[W�s,p$�D�|Fv��C��Bӛw�IU�d��q��S��+�q��W��J��l�xX�خ��ԃݬ���V`ў����w�C����[X��їa	��id����&gi`SQ�6��o��z@��J�B`.C�M!ܘXUS	��W�I�`W錔se[mB��<��Ɯ�R��z6��r����x����xΧx��y2m]�fk�����"k$��ƂԌ1�}����U�#����*�]�4��f���Fg��C,&A�>IS��K���e���5!)�\��<c�]����\id�//�k/���&�*#Qg.U��	҈�m�������i�)�=��χ��Ꞃ8N=<�'����IE넨YK 	u��u��0�6��Cޥ�kg�fǤ������]m��oTր�k��Ͷʡ\ԩ��4�)�d:S��v��#��\$c�jM��;Če!��r��?n�^a�/-���br���6�-V�4*���ʌ޾,@��G&�W����ʈ۽ؓ���@��G��J�3�H��j�#<	0��qC:�M=��c��c�h�Y��J*��lPa��&�i�-�H�
��M����D�)��k�NC�{*��*�g��)_G�C�\�km�A�~桤��ߍۑcø���9�O���jp�LX;��{B^I�|*���}p}gI�����������}4t�HD���8z8I��*֡���l�+g.�Ln��l5����z�8G?xX�M�Ch��]Aa`�O,j��B�Op�����K�*���mc�(�%���6����}{���Z�R�������Lw\j�U60������g3��W��}bXgb��l'��`�ߣj:�� ����p��Z�����&M� �@����2�����B���'+׉Q[��K�RK�nT���6������;I�EB���v��z�y�0`:"�H�*>p9=���/���\�ۥ���O[��d�:�pȄ����� ��f6���Ԑ3��~Bt9�W�|��}{�n�j*1u$|A���`UŨ�Iz�V����Gq��ٸyE�B��������V�y����wT_���R�fr�)@��Tb?����lbP�B��GZh���*:+4#T=��.Ki��"��0��J4ArT)�W��"W�3z��Zx.K<*L�k]Ĺ��@�'C��q{9�b��<��.��0�$�p�e[]��q��P�`ų�_C��g����Fg�\S�w�@k��}��g���T����(�[7�}Q�9�[_�\�N�c�O���e�����<Z�s�.���1�x(I7kD(,��S'F}2\s���cu^6RGhz�ng�/���<��v}%Tn�S��u�,�m�pD�yY5�f��5ԡ5p;��HF���\��۰ԉUl��zn����lw��[=ZZ��t�����:L�j
�XI(z�*��*�KH�r�}J52��[0�,T�b*:��HZ�J�c6�Лɪ�Z	���@ �?����|01����Q�h��tF\�C�+mk��wR=��kǢg��}�/rxf,�
.�j��2�}㭐:Z�a�qJ@�gh@�a�X��^ Y�.W1��"Ȝ�C���_cd� U�Q�
���D�� �YE:ި�F�t;�̬��Ȉ�gn��7!��5b!�}���
����?Ct|�ƾ�K�В�2�������^�ml-��xV\XQ=�{�"#�� ��I1g��m��_��n����?{Em�|�:��6��얐y�s�P�I��D��w�r�2> ׁ�]ۥ�W�$�]o�kB�hs�#i�wLQ
{���)X����Dx�i>�à�i74���U\�v���)Y�:��GƩzn�of��Dq��Ƴg!杕�5�5;6(���5ba]�ȗG�#���<�xbS�&�3��"�W��zA$(��٧�2��Ef�.���ƭ�8���J��D�G�nO�P]B�C=	S���O=�X\�`Ex�=[^����v!����&D�q��E6w���F�"��ѨT'K6{?w�.)�I�s�W�D6�p�%i���˙V��"�*�Έ_����Jt�< ��������*����iLB���
*H��$���VE4��&��LrDI����TV�]m��fty�;)(L��ƻ��S���D��ݨ2M�r��ς�/5�x�H�Ո���w/3��kT�g�P�/f���K�.��Hf�E�XƖ��o�1ㄍ�F�M3��
G�8�%L)e�� ���F1*;(�K����^θt,��~�푮�4�'�_���ʢ�a��=B�J�"u��S��A�R'�ڗY�;��ݑG�:��D�g���t"�+�T�$Xa	�i�^2�o�=����m2�o=����]��j�͘��,�e��u2����&���7\ioGBS -&�+��|�x)`;G�;�S[:���v&�Y�>�C��_"{�E�y6��t���#� ��t���4]?�N�
d�����������MwBy]�1`��K�.a,�;E��W���;��s���	���ٝ�`3/7`�I��ά`hn0Ho��Գ#K���pv ��M���2O���,���M���p�Ꜥi��LQ$=~MR%+���u�4����O�þ ^}-�M�/�g#�F�2��Zk{sg���`-�����~ٻ4��I`]u��}M}��+^�n��ɱ(����\˾(��	�/N�.�
�]���LJ���}L,�.�e�%[�5��1h�)�ڝ�M�.�4l�e������E��|k Z�:-� (�MH��2y���[��c?Zb����*���ҷ�����Q˓� �lS�/c�m=�AvA	b�r���8W�K������KZAm�d"����%��i���")���r%��l�=��mH��w5��ZZ���7J��{$�;]�H�mz�Ϗ��v�����Ċ�OOa�dFyʰ�$��wJ{����P+���e%Sr\*"��u�=�g[��0��a�*p����_�$�R�{$�.��/<�`���~����K��e6a:�"ɕ���}��%ʱj�'�B�w�Ȁ�F�;n���jP��$��ʌR��\�֟hm9	���q���JG3��h�O�F�b�2�-����n�a�����q��D2�����WW�~�͚����$����ƿ�n_�yܚX�I]��G��F)��.H;7��ѱhJ@S���X�(!�ڄ���=M-BrCg��8��}'H|�_���F���ataf��9��H4�������r�|�Q�V�%9v��jS��\��,H(��1�a*�#���_���K�R ��F��炅��UzhԸjc{@��3�_n�riv㙙.ͳv�$N��)YE���iO��.�w��Z�X��
e���^�!�
�ٖ=.Ao� 糴����EkH;�S��2T��]�����ro�*5���芎^Oj����?$>g��0k���Y����}���0�[�ܚ7�T�12)V�k W��Q~��\Qx!Wwq�=Z^��G��M�n��p�r+�ۂ3S���sS��o,C;N#��\:��StS6  ���L�]�5�Cz%0F�d�4�������C�ԩ��;��ؼ�2적3iL~�t߼@��&e�x~�C�N�?�����mc�� {8�3�BA�1����G����j�P��1dN�M0�D,1��g�4��w�M
�
�A�����^�d$�p�w^���&g�K������#n��.��^ �'Fu�a=B����Y�ME��/|�s�e=���;*A[wKb)+\?&�����U��p��ғ�7�mr2((4N�'���i_dNP�9a3|�ϖ���3��4&��K��Ѓ�̃�6�dd3C;H:�2���G}U��+"�_���bؕ��/x�����>��0���\��f�O�-��6��ۮ��Y������?��Y=�9�m��c�w7�No��|y��[���vFW���4ۂ�V�ȏ���sqgH8��-B?����-R;���HARZ@��H��k�k����v��df#�=��+�0�G��0���c���7(7}�;sO����,��������>{B/|{��=�7'�:�x�_�ʎČ��,-��8��������iZT`Ø�fj���v$d£��r�@��
�r�Qf��MƟ�b����p\����D�t&Y-e�H'�{��>���Lb�㒲%�K2�Bzr�KTy�;(��b������N�.F�b a$s��x��d�	Q8}�9g��r�2#�e�����";{�� ��=ߋ�|쌾��$��3/�����]� 4��D!�,^��͈o@?��1�� $�s���v�A��M�`�|���:��� ��jģ��c��wU��L������j�v8�4|W�~V��	zj�� �޾<q��V�((;?Q��8w���n�j��:�e���}�]��&�4���u�j툝��	{nT>02��F�H�)^!�(D��G�"pVa�W`�&`��!7�k��6��������*����3����Ɩy��UfM�NuD~�W�[V`�_u2m�&��?�eU�GI٪���|��/^Ð�Tv�6����;��z���ک�f5�oY�ES
��	���W��4��3��+���|�)҈����g#���{,�dn���t�w�5��v�}ˡ��C{U���Kc�^��A0# r�Ph(�p�rhګ�t�3w��"�O]
{bN���+���;;����X��n�>��@����zh�텹_ �ix�<��E�r��o QL6��}����`��mt��X���;a@�ϖ+�%Ծ%4�zZ�1�k�\*�DG�'���;dfP��+��iIC�MSb[��� �w��O<A�H�X@�����K��2�6Fb�Q����ݐ���"}�)y~��`�������.� i�5r-�ӛ�#z�Y6��Z�-2z8��k��A ĉD����X�E�9R�Of��grj	���\L����*������-$	�.8��h�)w�=����
��f�4_�X5y�״��Pue���/\M^(Z�B��B�mL0�y�w�Qր���?u����Ӊ��Ȁ�F��M�:��篦�q�1�W|A�9�����q��G8�~Y =�ֳ�j=��7��~/��a��0M{4a��V�+[qtl�V+���=��n��|��1,X�J���൬���]�ջ�[]<���_��j�Uh��X!͒"R,�����t+2i4�qr���!�˖k��S/���ҏX��U��6x�W�(��hӷz$����'<g
����I��1� c�~��m�H;�LG�^e����Q�k����>�ʗ�EN���R(�4��X2���n1�O���E�g�&-��?d�.�����|�l�^>���r6�iF��7�J��ݳ�G�@������@v�yG��~mѻ�h����E�O��C�@�U�ϸ�]������o-�*$����DEs�a�=�`k�!`>�-Ev�ֿl�i[�*e��--�5|G�~|��G=7l���y��v�6�?����pim9q�G#�if�J.���ڃ,p+�3�H�@c}��]x���&�#���_.��~_�,�e��-�3��a������_�K�U����;�\�H��2_��:c�� >A�B��lG���P���H��Q�L�۱���Vs� 5���އ��z�YEG��^��:2�C�/����%�O|�z�S	��$�>�W��s�t�c����*��<.�K�x��)`&L^p56(���^G�m'�.�m�S�!���Ԏ
n5_���71֘3P���������(��	t�P����T7�����+b�Y_�;6��v��ɛĎ��j�0i�{�,�f���R�~���ϼ�łD�ˁ�Ƿ��h��y�1�nM����[�cxu�z'�����HR,�e0�]���F�����|�3o�`��?��5BG]K8�jOF��f�C�v_rc�C&|M��A�������!�7{����[����|�g�k�%�����xt5n��ȈM�֥�D�Q~�`R����­p��*/�0��!�o{31��t�+��N0bia�៎mu���ދL��#�Ϥ�G&D���S%5%i�������U7�\�<�5I��ok����1c�=zP�̤y1�ViIҞhD�[O?�����Q�FO}D��W(
0��wy�pK؃��q�ǵ�r���F3H��^b?�{_u{s���� s��Z��Ȣ�.)n���j��+��z�0���޹Ԝ�8��,�y�E����������kN�h�EhUp��7.r�9�q�El�.���I�\X�sEͬ���wr\LYa;p�N�S�g�=�XV}�V�ḯ��RN�,�A+�tQ�2z%"-�/�oSJr!�,�hi�pk�jG�����0����$�յ,R���Ǹ�:u^���G
_�PĆ��Go7�j`�L���)���Scm��j؊���n��[�6%`>\/�����+��py'b��×���7��3PN�l
�.oF�k�o��5)SX��~)�Y�
�	nM�D�<,�m��w91�|%�S3��nz��j�!Z��jsw��Q���^7k$�o��$�W��*P]���I���;�*�8@�J����ӥ}��V��!�0Oj��ʾ"E%��a�r���Q}.��6[��~���>�Au* ʛ��D����3�N����F�K&x+�%��0i���uM��!?�A����7��7|8�4�&����n��Kv��ó��a���<sl�gYk�"q@cz��۲�7A��$�iGW�w(�W���@W	Llk�j�8��+�Z�s��#�T�2�KCp��|�:ם��>��n�:3� ������&�VX#�uN�[��;��˹E��%E�%�!�h-�r
3D���\�_mw�7���QR,!��{�=u+|v�����E��"���o�G=�,h�_���L����T�>�k?�b	��0"4mȪ���h��([��*p�+Y��=���q�1)Ք<�ΟF	H�/Ъ]��μ�o�G��2:Y��:ѫ�.΁�n3α^�����9�����E���Z��=�׋�پ�kED�P�7G���$ؑ�����W/R�	Jw��c)�`^4�,�s��y�����|Q��4�&�kҵ�}�0���[�A4AL�A]�,�JC�ZSI��{���[�PoOox�F�������g��\�;�C:}�
u�πw2O�)>W̐���Cc2'��VF��2m���/h���K�.?�´;�V��6>�FI�J�|TI��D��D��78[(J	�S1td��?+Aom�M�ޠ�k������:��N����ts���	Ϲp}�a���˿��Y];�{~N]JT��9�D��t΄ɨ�di4�`"�e�/&��J�o:�0��'QQ�����Sb�?z�Rߗ[����J��_k9[F9�x$�BP�I��!"�t�e�����~9'v�W@7H v��nkѭ.�^��vO��
d���ݖ�j)�q� 
r�pY��s1�O趜�h86�����A�&.�K{�AB*�IE�����	�]]����
�ꥄ�kB��������>�e��#t(U�݃Of���!*�����16t��eA�:=g�P����\�/P�ߣCHd~&<���w�f��7Q�^H�@�c�^
��3�����;���Z��ɀ#ٜdu����G��g\��p��А�gb��J��S!3�\ފfwC^Q�]��X�VN1f�h����6�aũ$�sX�˻Ť�Fd��|ٳ��WR��%^���t?�3�a�c�g�?���JP�u
��}�Ie$����!<��1☎�d���a5'��P�3?H��X���3W��� �Ig�Vu�Zl�2Oh�E��������G�U���M�$a��ꈫ=ɢ���^ ku끐�BE6�M1�� �{�������U_�X�'�e�I� }B{�<ݿ,cbCڍ�?0���Jr��b����ض��Hq��CR�$���8�L@��-�z�
���WzD��l�R&k�4�fzTthM$���k?���2Z���R�fJo���N����X����;�#�� )��/ �RE!a䞪���r��h������-���K�5
k���t��h�u��$���� ��e�F�z�ȇr�*j��S��IQ��$"���U�8˅�B���E��~�߾�)$E��#��픩�X�S�a���7){��r0��b���B�0T8>B��s�Y�̣f���ǃ٣��i��"�*�<�iE���+��e��f��)ۻ��^k���:����r<���'#&#Ay���ҙ�o�t��P���w��ݐ��g9$7�MD̸E����*�k��"�Ĝ�ܼ��%%CA�K��UX�O����xӍdU�O��o�Uྀ�8�2��ݑ�ٺR�rq��Q��b}��J1'������u�Q[V`,��F��ˎ��ި�bO(:����x��ޥA���9�]!�;��)4��u o��}���Jy�aLw�Z*�Y�H�bp��K₤���?�T�Ն�5ڌpXw}K��J��+p1�vq$�v\<��o��E����W��Yʕ��&9A�����~%�|O���%��18�T��W'J�X���sE��M�Y��(<ZNj�Ǔ��˺�15��Y|	ȁ�6��vD�����44�޵��޹�c�Y�jT��u�H���>M�jr�e�U`�KEkT)"�a�r�_e���2`QWD(��z\Tz�#UM���Y�Az����������`3]g�S!��B8|�qe�֡���LA�F[��jbl��&{�@�r�*A�\Һ�M�xޏ���s�ʹ~DS:�!����w�T� O%}Ұ!���@8\u��q|���2d�2�S�v俛Puπ ^l��Q�t��x�c�v�{W��������ӷ{�bN
� �����K�1���O�z)�h<���8�i9��;R��u�z��uo/��3(+�)�Z�$�V^bU����_5���	w�M��Jn�=��� +���6Y��?�u_�_qY��f�I	ㅬ�L�/_�,1������rl7ϊ�[�1���s��F���M���:0���nE�1Y�B�[����b�P
��Uy������;^�p�`�Y?W
?|Fm{���۾ٽ�&F��)K���>S��낽�dP�JM�iB���,Q깓�L���"�k��:�Q	���#��ip]��C��x�N��|�E]��BX�է���,��J*I�c���� (H4s�T,�I^7.u�.�rJ���N�g���dx���]�tG�K��T�rt����澨�z=f��V�������i�uC�K�g��Ԫ p��
�[� ����vHU�2ћPRT�����UK��5�nQ�*���ݝ�ceD��%�荩(XY�'�2�)����ic��ө�틍l�bG@��+�G�y0=��%|��$mKA��F~��5/[�:\�蓯=7��V�-������)p���B�r��� �!g#j_�\��� 	�&��[�͸��عd���z�S�@�<��F�Y��`R��$ݒ��|��FĤ�� ��l�R��/��	.�ܿǵ�u�<d:d�K&#��֔ �l��<߿$�,� �	c)��\�^��v�*LmXвV�߁�yA b�B�?H�4!5�{v�n���Yr15�w���A@�=�;v/����wtʧ�q���HO@*�uһ�)��U���B-��x�u�����	U�POIM2e�T�y�xΞ�ɕ�w;!������A��;+d��?��P��byR�h-3;��wlL�������9$���n�u�༄���<��P	���z���˜Kpi���V�ޓ�aT���1���YD2���98Z!�U%�I".���뾚3%p�VxR��/��i#�C��`e׈���w�e���|b����q���(Z�v$�c#�r�Xn^�m�Ϙi��R�ԟy`ܻ��F�ܔǺ����c�Ql������W%�w.7�Q֒R�y�75�<�K(	{��}� PV�>�6[4��T�5��4�`��>�-�=����Akt��}��4�"�Y����.ßk_�!�n'G�Q���`S�a@c�'U���2���9�R� �{�����8�L�ԣFz8�R�H�?��*%��-m*0u5'��� b�����M`@�b�.f�{�r�-ӗgjƍ�|?��s��]�+�Z�?����5]þCN,:�-��&3�@��0�����$��$�4!f�lP����yVvJ� �r_�<�V��I���?z��Q�!��s9I��� �p��x�~F�q>�S�ް�8?I^^`N�]�p��i�%��Κ΁�̐��]�T�[&�/a�Wg�6��['$0@J�P�e;�;�M����ٕ��EJ����Bq_�:�����8�8��������o�梍g/����þ��yP	&{��{9��g�fm��㷄�nJ!oN���ن6�Lz�d�SBܗ�����EX�5�kN����EO�.���Ύ��E93�J����ۗ�k?�M�lM�؃}]-#t��7���l�/z���1#�8<�g��&(t1,�����Vi�>�}K�j�����8��u�i����?�F�ۤ���h��Z��0ȓ��7��cɝ>M�*������V>|W��a�:�����ko��jq��b{���w�'�Ly�z��G���F���Wu�t!���F�1���0]�/@��Fk�����׭b
��߈a�_ѩ�	[A�P�8V62���$����ݻe���'5��`�2Q�e������u(��[4�2��l�;��V�����d�i�ףZ�2&J���^cf��OCݳ�R�G5$,D=��KG0�D���k_�u��HO�
�dƟ ��Vv�� tAAV�5�D���t��r`���%���PǿJ�h������udN��#�->U	5rw�l@�?MP��(��m���n�a��#�Լ/��!��_g3�"q��0��G�,x�;LN�s{IX��N�\��&�%�.'�y�QEw�ʸ���g_�H����RSm��Mt��yE$4HS�h��xJ�:�b����n[���_Sk{r��V�/kARԲL��3�Ue��OTu"��W���"!�Q�CU��(vT~eۺ��J$�0�-`��l�5�»6�8�c?��(4��$N �@�����1lLz<��)�yL�Om�[%45��҅.5���ÀLG�T�m�?������э�u�eC�e�K���������D��0��"������[{IVʭ������h�ΗI<�S��sG�C,;���!����i#}|q���dUȐ�OP�*4�|�Jk�4�G��Tj�8����n
�UU��?���n}�%*�]�t�%�̽{.�D�ue \�!���F��zp|�s5@������C���kV��n%c4�?��>�&`�#���N������ƅ����@~[���0�#�v��������KXK�$��T��;��&tM��O�l�1e����^h�����Ӟ����E�&8u\�V�.��a�jRT����A���� �O	Q#)�����h*2�s��m�H���?����S;L[��/��_��;�2���`G%�<,�5]B	�S^;�g��G���7���|�Z�AϞ�z���_��{?bR���T���N��b��J]B��1�B��!�%yJ������v=#W�
7k��B4��ʎJ��"R�֙�=�8E_@�it��.���Vò)��Y2K�N(��Oµ�F����3ԗ������?ȓ�}��!��;���ꌄ����΃�(��>�%n�`)��.w�
�D��	�G���R�.�*�����EC�e7O����=�����g^,�7�̳��g��T������4�҃��;���<�A����^pr@��3E���P�,h�Ց1u���=3��Ժ��	(�*'��b���(�d��� O\ZH{���T\����|��pV�=�N����~�*���hD�Jr��G�1��0��m�/��WY��x�n�y��b����e��B�!���h�#��h<q��`�E�n�����S�aE1��βY�1�oZ����-�[�P�1z���;f&��n�/�X�B5��'�۝�?��zca�'\�&g��X	�,J�
}6$�(�F���'	efp��	I����6�wY3��wt膮tz� .��1u.�����ী��`�|-&q��e�X�b���4��-��3ա��c�x-Ti�-�iwV����^���Hb�i#<���8� :^���a&id��Q���ƾ��	�%�_�&��UV�f� l�4�Z����o���8?�~ra�>.�y��O٣��-
��;�J��f0k��؎����E���V=�m���H�6H�:��X���b)��C0a�wL]�H���V�ąIO���̅��V
�,β�j��7���	}9�D�42���{��Y/*o�U�gp��0��.˨���{�@"t3���ʟ����b�@Q�A�s3qɃ~6���tݰ@����懫[����>�T|5�?�Q\Ŝ�S�^rqD��eK=�9Z���#:l�|�ax�}o��1ԃ.����uߊ-XMh�d���!���>��B\�AՑs����x�vą/�U�5)�Ϗ]C���J�ߞq��c��;�snx�bXP�g��?��? ��[K�]%�M��,m+b��:���K �+�;3��?���&&����ĳ@�&rҥa�_�q�'l5���f�E�`sM�����z���
�#E	JF��
�
�� -eX���!��{�Z�l�>.���AR}]O�M���yݡ��2�>�wuh,6Rcu&F��h��ŏ��4����P��������f���,�<?zC��o_U��jOz�B07��P�����$TG&`��!mJ����gМ�{O�����E��	���3�y�����J2�����c_��y�W���<4��h 6`�Hy	F���+�X���8�a��� '�uߐ��s��I���pV���s�o��;��cy��&0�㨐H�& :���"[� ��{�="�]3 
kk��1M]Թ���i��eaz�g�:�f6�"� ���b���,�u	�%�L�����\�.i!-���?ؙߩ�vtՕ��.(���.�Z�9<�/���ɱ�\���N���7L��I��x��\�Dtk���`|�ks�*/�
2�/�����T2�h��yO*�8�����S�)�$yY�.��0v���Nu�/�*������ E~>b��,�ct�I�L-tKђs
����4������T��1p���H\������#c	���`�$ѺTG��
N�/ѽo�|��q��>�<>g���͜���uf�G����7��Lz�`���  �l��{-Yl)�E�U5;
�z
�]�h �^���3}$�@����
B��;���.��2�({���@��'�"6�u�p���yK1�b��$����.p�����5�		U��P�kj��v�%u�P��d^��.���l��͛��{5<�q^xb�tR��JQً~	#�\S�r/��`�ѧ�z��� �#bt��R���O�~b�ѣ&��d��g��WI�[H��y�x�K�;����a�Q�)�D聻ӫ[�I|`a�Yש�W�J��>����l�O*׋'&w{&Rߍw�Ӡ�=pf�.�Fv~2�s�͏�ź��z���dI��V287�&��m����G�$�Ҝ�7뚚����mv�g��dd���M��-u2�O�e���W�a��yr4R��ڠlSU��Ş��~!.SeU��u)���C8zM|��]&4iqK��4`��=q%jQN��K{�&�(I8n5�4�����o-��������sy˕��Q�ٟ���IL�w@���$8�w:����W�6��Q���?���l�����ډE�F���{5�����Zlw�\��/5*��?�R�g�L �Pˊ?�Q9��Ě���Kj��DRtO)�I�"a@�f��s0����|�D�k�Wz�4+�q�;h����i�`kY<�A?�]�5|V����5�ܺ��5��������B�4Vҗ}�h_�#�}�}�Qt�D/�*�/�H�6�,Q�شZI,_�0�C���>���$j9�3Vڶ�I�|���%�	Q� ��� �0,��1(�xC�<Ǌ-4�$��!Zs�-�e6���w_ۥ��=����%�^��0]{Y��9Z8�oڕ|d���R�����F��o���i���Tp���w;����h@��ߊE#�m-/��cQ�k�N7Ip*���ghOӈ���1nMï��GN�џ#/�Z��"�uS�P"b�{!��1