��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���FF8ZW�@�Q~o�G������ذ.|_Y(��ߘSaq�q�Ƕ���f�x���^o���q�Tq1�z���f���**D��-@�L�9g�iľ�<;i����+����j�R�5g!�%�M��q�� �œ�$l�Tș��%MμG�G0ܞ���`�]�\��Cͣ����Z�e{��2 ��R%�Z�bf
��;=SY{�kE��0�	̫%U�#}���E��d��5�@�� -H�s~�J^LcT� b+���:�X��`�0i����Jh��	��J�Mt9h��[�!I��W��9�u�:��҈��6��*�$Q�|���7\�2*��\���]��[�Ys�; ���c0�?c���4����x���؞��,H#F�R�'L������(ؙIsǤ��|�h2�;#ap5��$�K\�G��a�(���)6 �LzZa�x��:Z �(�FJ~g��Q�P1)���߃@س������Ĉ/��Pt�<r�Jw}�V�<�xE~�΢����8Q2�_Q�!�/��R������18Y�7TV_ea�j]ޘ��21���mȓ�`��r	Gm,��=b��d��5�����TA�zN�gEg�����ze:�������� �R��z��ڙ�9[����U�x0����e�S+�TA���|���Z:�᝟7 ��2R��`�EG~�ak��o�۹��C\[�fකa%,n���s������8tS�����A�N��4+��u�y���,�|�W��p�?U��s�H�����0߯�4y����a���g��xᲨ�J��5-��"��C�l`h�����%���~<ݽ7��.�%C��jK���Te{,G��?�}�	a���hM�����R2��܂^4?32�62�0YF��Nλ��PM��ހU���I����:���q������I�_�V(Vv�ޫ^��j�T�r6��"p�ܾ:��Q���x:U��Dl �?�t�	�0B�s�~�|{���
�-��%�|��U/���R���|9	�� ����%�W����\�:�6��OMb2�G�E^��K�=H��A�k�4VKi��, ��O�t�S�_ݵo��P${�uAPY��2D�w*�L����G""��5$N2I:�m��Q�ߒ�3���Nk���j(�L:*����XT���?�)$��qS�@,Ig�/f��+�#�� ���oD���[rq�X��nʨti���vG�|�ɳQ����x��n�ʙ_��DZ�)D���}�Ȥ��]��������nE� j�9͢��.�
�|V�m�p�_����:o���T
�����yS. Hl�B'̹`�>bwodhܚt�.�Np��֐��夃�Q����Y:�'Yb�C���0a^ܛ��SJ�+po�y��Q'���qkh�Z��JG�Y���}I/�����c.�M+�4� ��9�1�o���G�s���T�x�ĥ�eƯ]����$(�
kI^�5��( ��[x��@�V� h~bP�׷��`��8_O�!|c�SK�U_5k�\s4ߣ/��D��s��OdH�"�@� �Q�{r��~V1���jǷ�PB��՚�#d��1?4�i"�~e�>!��@�u"��� I��A�o���;ϻIE+�I���ꢥ�+�y�>�(��#^�R-�i��X�;�8�*YliG�_<3�ΤΛ32SJ��ߕ�B��q�LelJ> '��6h/+��a/l�x?C��u��xIa�A܉~�f=�իK�[ k�ۃ��]��S�l�M�1ڜ����A�s�m��nH�]0�Y�4,�R�G$��$gzܻ7s�lJ���-��5I�Z�u������s�Y���TK��|/�:G�6�ș�`Fg�1��5ϡ���, ��sv�h��eg������18��r�:k�d�6q�5�􂬽�X�^r�������֌1"a�J�*�����@�v��[S���!�1�.�-���/��X8f�s��0�Z%�/��%�$ŉﺻW��7�
K�`��a�A"���g��K䵻}LPx5��O	�%�)5��vgw�E���ٹ��^u�kp1uao
�,��;>+PP��nU��}X�&�:>�����'���vTF!��M�0�Cǣ��>akP��}�\�r����\��%�fA+���E�nid���h����=k�G֎��c ��l.,<PH���T���55	8�u�#�-��4�P��}6N����MTN�q�&ק�/)ܸe�(�|�K�r�LnQ w;�_9R��zݦ������C���ĺ�c��h�V	��|N5pґ醒��0�(9�,��g��n���ST<W�PL����C������[.Ǉ CEA�,������u�$}�h�������{�\����<]�M�H�֪��A�T����U�i�}�sµ 2�2�|�(t����-=�0ØƮ	o'�]��\�a�ݜ�m�]��Ʉy�>jT���<����5^�"�N`s?eQ��i���s�E��{����۷�Z%��]Z��o8�_GvZ埆]�5�ok]�|&<��U�WL����s��!�]��?\�o�*�Y.�SR���@�H4��UV�7o<p5���V�ғ&&�A��
��:I-���Y���)��>m��{:����%�3��e�X���kb��i5�=)�dt���O�Ps��񤾋��~7U��J3 �-2�@�`T76*(�T���:9s��u��h�G���5�Bz�Wi*�8i���c�����j7}���cv��&���]��\�},�^����*>!�Y�<��)�����AT5��;R�[�����!�@_�:����=ĝBx,�UTS�]�v@�>cV(D/�#���Hw��&���6�mQ�hj0	���Oj\�b͎�q�ܪ0�F2�<kuZ�Gt�9H�{)��j�E�ˉ�z��ջЃ����_�e��t�ơ>s]2D�}ذ=���t�om;XS4����
%�[UM4L�W@�f!l�+�xC@����;�~��e&d?��t�UXԊ@��XV��jbKht	e�:�Pɽ�8ng�
=�2�n���R,�⃐�C�T�R���h@Q<Ǥᛠ�jf&>�N��j���!��ռ���{R��^���ԐR�%{��~F��S �o�-F�x��	y�͜��e�����+W�<��Ǭ��R����B趭J��u���W\�'��� ���I���r� {�0pE"����
��h���lN�AN	�&_�J��u�'��i��X��w��۵7�ܜsU��rB@� ~���e�M�Ea�H�p'T��v�kzNLPԝT
b��'��]�tGz�}'37�6ҩ\w����~��馱n7�^T3HC�be�Z�Q�Vİ�9։gg#��lOG�Hw�ƙz<�CE��'�b��ԫk� �^ϜIK:ee��]��"�e�/�N�N����V�.YQz*A�דu�vJ	M�����T!�{	�g����R���S?4�o�7Q�C�̔>�	/�)�8Gw3�G
H����N�"��V<�=����{p6֧�WI���������oo�AfZAv��]�Z��(�>:����#s/G�_=�T�5΋!�T#��3ķ�wɔ�ɣ���/��]ru���ԗ�B�s�B��]F� K�\}��y*G8n��c��������~���=e��CQ۟�
8����S����9�mi�	Fܲ���(<�*�hApIn=LɘT<zW�GA��G��y�pHo��F�)s�
�}6rj�G! �Ak��X;��NCi(�q���Q:/�V%�?e8%0��	1˰V���:�lfC?��Mq�$?hJ������t�\C͸���'�㣜��f�֪|�2
�cd�KX���M�IY�]�%�U_
�'�hq����T�8러4gǵt�RV7�.�.��0\}Gܱ!��"/ևU6��#?��YUڙ҂�eeYB�j@].�pk*t1�������(_��
�n ��&%\(ۋ�����n�f6��6 ؆?��`p��r/�C��n��`QQ[�U�@�[�U@Q*b�Ц���CН�f��ʐ٩����5%���T�5z|�SJȧ��Ad�l��ӑ��~�~�;q���6[�(&Xk>��n�4��xw����+�i��lЃSw�����(�;I����������Kq�j5�����*Y�o̺ �g=C�%�?TOV����:^C�ޛ���|���gV�8K�a�c��ʒ�h�۴�5D>�L�� �eך���	@�ڿLg����	S߼"�������E9��}bY6'��z|"���4&0�NO,ٲ��=EcN�p�_��'n�9��B�sݝ'��7R7��J#����~6]��M��OR3ab�0��u�&[&�L�L��g���"7l����  ��xW$��h%h�!u
� S��r7��齍C��~]��(���1���,@��%4r:o�WfWf�
�:���:�$u�C������4�c`�R��vw)�A{��� ��
4Lߣ3�/�Q?=��uX�8;�(���N��&�̷��1�=7ɓ���+7�1�p���N!�FI�;�^��������Rb'	�]t֚y�v�qde�nˬ�Ŭ#����	��=�`�'��5X��4Ћ@�w_�j�y>=4�3.�h&l|q�����fo�k�Z2U<�,�'S��O+��b�xgm7M���V����Y}˛���vt_dj6���qUi� ,+�i�C�A�R�6�paH�~]F�v2�2��ӎz��(��Ӕ�������c�8�����jh~y-)fe,s��5���^�������<�'u)�r�*:��p��3�_�J��J���g�M�q�J]���;���d(��T������E�F���^Z{����]cfl=�s~妙xˊ��o��|RY46��Ke�����鲆<��
�����Ɛv���Ba\��H��t��}�Ey'���4YFI�|Ac:�B�x�/�h��T��T�9p�{�F�zMK���@��2lD�0R�i�P�ծ��)���z��8:���g��}�-Y1C�[Mi̼�܊�ڧd2To�4L��^Q��)�Xs��V���i/TH˅R��Õ&�������QfPler��a!�[�}'!�%׋<�$�g�-n��[rG����l�C^��7�+q�b��O��t�e�Ȱ�lH��~�T���x��I�v:��9џ6
6�����I���1�3;�f�ǐQ� Ǧ�_��~�c2�����-~��Z�����υ�f���_E!Q�нg@��)�}=����+羾�H��<��4EόR��	��f�R �)��"JO>xk�~�<w�BRC��X+�l�G���z�^}��ɐ$�^-б�`�&q�������y(B�	���ߥ���'��m���O�� �P侐,�b�㉁����U��Ԁ����>�yV!1K���������_j7X��G���<�Ҧ����^�X�����p
![%�Җ�"��7	��C��6j?���c�8�#IW.��Yt�	:-F_���y���5��W�.Ѵv�fC�a��/(���"'��Jg�o�+'O�62p1���\��|e_k��*2��
5Ƌ��擭ݘ�D8�4�
�� �jt���L1{�kķbeF�E��]���W�;�A��7*%ϸM�Hi�n<�a��W�� ����B��hE%dĚ�Or�ܸt�6���
&I�J�D�:hfW�!�w/����R��4  u��;j�'�����"����xE	<hՇ+���5�!�8R�J���������b+���$XK�����OM'���O��\�aH����QV�*��~ݢ�܀w�%������P,	҉����q����S\�͐uw[�%�KW����0`N��n��*b���O?=��;�^��Q��c�0^C9�)ul-C-*�8#(�Ͼ��f�(?| db/�/��S�IE�Ӧ}�j��!�A|�O��>�p�{B��7Q�W��$��y5<�� �j��ݵϓF.C��1��O��]z������A����R(�~��qA�9���8D&�/y~BD����ON\�!a扉����l�j�,�柱gj����<Mw1<U��:�)�ݽ6^��_��~LӀ=r�L�K���N:���U�����xc�]�Z�^�;�0��\o�\����WvZ�J��|
N���Ch����K|x'��+a�\眿�N��7���Df��m�|_V�k�y�b���A�
ۀȮ��RFUP`�l�zM�d��P��K7��j�<y�0�Q�dr~�%_�#'q;Y�Ҏ����~ؓUg�3L�@j���,>�#�%;7ŔS"��:`T��_��|�b�����;l��T���ڭ��a`��q��O���H��8{-�-���,�tn�s�J��DRYF�&�!�h�۳s0 M�������mzD�|��d~��J蟫���4
�W�f�^*I�
�(�1��)�Ў��t5v#�5��������b����%�\�OY�g��V\��?���D:#�@:D�l�$����H�QL�by����8��B�=˶�%yk�A�����Q�(�Dn8�A�/�͑��'s5I�;sS8}������T�̊�m�2���1��5�PhEY;Rp��?0�����7	�r?#�c��(7,g� b��=<�3�lMu(-�xu�:�@o�%�ȺW�m}���g�6�^@�Xe�L�C�H=J���⊀���{��/X�Q��h�u��8�s��Ӊ��nX,lk�%C����?�*H:���g�E���fFq�)G��V�6djsI��)��;۷Ϗ���T��x�!���L�x������nMk�D�i^M\(�!�����~����r���Yg|\V�ۘ1��)U�@4�+N�U��T��YT��Kn]Y�6� !�i�`�`�������)e�-R�@�9Z���]^���ɪ`��4Yqf���S��*�
����:L�)�w�'���zhY��	Ҥ��N��[{�֮$�ƚ<>��E��іT���2�%�W��ʫ�[���9�ؼ0�V9�%hd�Է�|����6�A��Ѡ� �*�>Լ����WP�u&�Z�P����E�j�*VR�U�.���&p7^�}Zs�#)j01�g����Ӳh@�h�Jm�#6�Y����Yls�ll6ݮ�Q�
���Ue��~�8��Rϒ�G���>���0��x�%�!H{e����od����GO���{���	��˶Du36��PV�l� �"�n	�R�P��z��й�Tߎ=K�@"-j�B[���&q۶g���V�»+�4�0�i'im�
��A�v�t#�릉�c6��xj@�B�ci�)�P������G��/-�G��m�)����.9E��.7c႕̠H�k'm��\N�x�^�����=�K�ǁ����:�u��3��L�ͫ�;��\Uy�3�pV�vTlE%�9ﭕ}Q�m��B�-����D�%3����Pd��o���zR�;��S�w2&f0rj��[2~]�W�ו�æPTK?[dB����(#H��٧�zWmI���������d62��OLn���R�%��u9P;�X�=�x�b��ĦL_��c�t%��)�r+�DH� ��ɇI��M�mR>b"=��4�����|�������X�2�?e/�&�8%ӌ�	��B���f	{!���5w�asP��'�ro�-�vd`05���-�Ѯ�ڠک�v�40�G��,���<u����򑫧=�:�����\���;���+����ݴi�,sI�M���?�G�p��ǿ
/\%j�'���0�A�sw�ȕG͜I:�q��3
p��:����C��l�$�#b�)�V�Μ��+Yy�C^/��������o����m�VJs��{���6���L%�|��f�f����t�?��Z�