��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t�ĴH!�7FA�$��b�����y"�T��d��_ق�f�,!��f#/��x����&G�[�Ʋ9���{��5 ����"�y�{]ݫ �ed`�1&��X���1\���v]O���8����d�3�=���l�ӽ4�*�Ԥ���dţ�vV"q�'���lWVE�{�7ۇ����b?$�_��J����F�)C�FH�rN#�����(�ř-�������#!��,w�~���{W���V��v��!��25�J�}���ǂ�u��j[��ws�5��_�c�2�Wa�&���!'IM�fт��S���⋖��]Q�{���l?y�Q����
��o)�b���u>��*��j��8�L�c������`���+E������,<���M�>�
ʵ�F&i6��o�_V+�Ks+s�z�e�pY��o�sy��Q�F���h�'qb�Z�(���g���0�Q�9u-�տ��Q)$��1�cCV��ɰ���6�A��V�T�X5{��Si�?͇�V�{c�݂s��{&����VR!�������I?-���_�wS����²U�>^�*=�ԅEa��א}�`��3 �GH�Ș|��n~���w�Q���*�ȷ�IazL=6بgz���m���[b֟��Ju{F����4tʡ̞�{���N]�_UG]�b���n��PEdJN��N�4J;�w�`��Ѱ{�IMX���V;U��`)1M���_q��dj@�5��^��n��?{rt���|etܯʮuH#1*b}��&g�ɡȂ�?�Q8Z�o��m(-\"k�f\d��������p;#rn�ʺ��	%?��t��@hQo��r��l���
M|�`'����L�ZÆ*��g&u@,Y�a�&����[�>�f�Ӕ��7:Ŕ�#]��'j�H騫�1�U�ذc9i�dT%2�TB~N���*{�&��{�e�k)"�(K[5d'��Sx��R0����d�	�K5	��NIJܺ����9��=�,G�J�����Q�����'H�P(>Py��ⁱ�1���?3s����<�^�0�2�Ja�X��,�!���D����q�E�[g^)�3�/��9uY�S��yQ����1�����gF���sZ��f@u&g�M���W������-���(&d>�_O�kI���M��uZ��H��?.�Q̟w�z��G/�u��nj��3��g[鴪`�\0��shTa�����͘vQp�% �"�v�Q-�?N�˻pd�~���.&x��"顷����<P�h����(D�$���Ii9˝�K�^�XJ��q�z��VL	����/e[�L^d�ۉ���ʴ�.�Ff��OkЅ<��!y;��֎�*K'�*���OniE�0��R��ܕ��N���J��N��)Iv\�"�ښ��eZ�3�o�}� F!��/���G�Y���	�%�>��N6�E{�E����7�uu���*��΃��
Z(I�V�4^����$�#iʋ�w��]V�8Y7���e9�9�����0閄�C��y\�3툏�y��w�&~�b�B� #pR�9m�,~�F��ѭ���X�"�ԲoV�扻�����)�35�ו����+8/j~���$�HJ���_�N�~���S	8���~_<-�:�&Ϳ0�����W�H0zUﴔ�Eg�Hgb��S���g��TA��W����)E�+��u�g� (�ӻU&�0�bN�>0��Μl�_�oT�%5���W�NO��X�[J�E����*�h�>J�w�b��vF$�>Q�2te��'Ӥ贅M%)>��u�i���@p
�@=Ȋ���&��Q'�-pƫj8u�=|�>D�'8�o�n�|���m�B(0ڞ=:����"8#���@r��9�?>�F����D��r�6ZjJG�
3�(Ƙ-)x�>�����@�"��T�&Y�ue�֓�h^p�+զ���1�I6�m������Y��ٺ��]�����"�d5��CW���o_��8�U�U?lM�l@��ɜ�g�¾�$� *�{����+��v�Rw�`H�V)�]��e	�B��$��i�ጿ�eH�<I��"�-a���D�Vt�i4��2�R��Ⱦ�n�)���"��ǚ�2^p�)iv�>x���/s��!�N�)��!�Ӟ�\���'��ӫ��������;���^��7Mn�3��bwK����tn4@��� ��G����0˽1���}����y��;��8Q>�l���A ���%�$A�P�ŷ�ƕ����>�٤"�����;���/~�nXY��)����Э��IZKH��Û8-��kɨ(Ι�?��q��O$�8u�� N�������rI���lt�ϙ�N�_ @�	_�6�	�E�"V�n��#'��&���B�H{Tq�"?���O� Խ֔���X�/W�� �I{�_tbc��ה\�xQ���og��Q|A�! ��)�������m�iA����2S�au�������rX��"F?����D�
G{g���$����''����,��`��w���,G̘Th+[�#�*8����6/�ѭ�fS!=����8?��ȝ����!:(H�X}+��kV,KU
�t!�5�e#1�y�������M��%�%�R�u]�H$.�AzBM���3<N��P���3��c��S}(��ф��9�$�z�u�z��ǈ�/�ŞN��uc��+���i'3��(�es.B�CY��8�����M�s4�i�f]Y%� R���>��ݔWǚ�<<����`��&������������O���6u��v��y����Y�č�eC]���������?�-DUϦze�6�kd���e�5A��ȃ�)6��q�NB@NjU>��ꘞIQ���
L�2��9�\/[����L�\ �M֊o5h
N䄭��&=�O�DS�ch�|�t20������{�Jz��"���%��;ԫ	���F�����)��ʋ��zLtW:��0󷏔�Ïr�?i0r`#X���R�ŕ;���1H������0uk�ܣ�%��)�9R��WzM	�*�K�ur�w-ˠs��B��t��Z����l��83	�l�Q��ҷKЩ	��){� �� W�Gc�wn���ݠ�j�8>��F#��ԟ߈