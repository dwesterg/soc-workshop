��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D�N�A(��ގ{(� ��ul�l��i ��џNr�:O��'�k�>l���.ɋ�O죕Y��9z���%��Z����7 ꝎI,��Ȕ����w����5��&�q=�����#
������@��=���b��#������||̓��i��9��=��h;m��6P�?h�O�{����}�>����� �?,foM�5��O S{�1US�+E�3[���a��Diy���ƒ�W��5 ����e���&X�1��%�#������i!��K��|��Y�lV���ݐz����#j`��wέw����C4���?(�R�̈́�ׄ�i���H$y�������	j:���{��d6��
t�|Bۘ��D�Q��y~��ES�lr۰��#��Y��z�I��hHN����EB:=! ���$H�r�窮7����������\B��g�`""0�\�S�d�\n���/n��6���k���ϴ�4.�u�>Q�̭�8�y��b�T�_TQ�T����Xz�ۯB�U���Ѧ��
��W����i�l>���{	9� �x��3��nv+glt�_�p;����-��]��(��C���vͲw��?���^����r��y\�B�Q�e	��Bؔt�]����7dŕw�m�˞4�L+7Q�L�����H��q\�ALCDy�lW}�{�nx�j1oI�O*�C=Aȡ�W0�*�n#K�=3P@��UdI��<T<r8]�#{�eQXj�/1�!����rη�z���v���T�� )�	Ӟb�%j�\Gv->����dNآ�q��kD7��>�:��B�0��\�3ٸoi�91��r@���^��8t<��d%v�60�o�� ��x�7�Q�V�k6,:Λ�*wOo��a��QA )������5��WD�������:S�Q�i$�ː%L���ѡ0��<���5ݗ�*)XR�_]w�44H��tĤ|_�`��US����}����V�Z�T���w6�bBH���9����z����P
W������P379����#�V�p;n��P��8-�uB�.E���S���Mv�%D�e=�2]A�E��kPs0А���"��-i�n9�v#�9^�����F#׹:���G���K��J��͛S�N���#A������;�r��>F�%�{�R++� #�/=������N��ȩ�T����`c�#-�E���7�=@p(����u@�����]t�ȷ}��#��P�̅�I�˘>�� å�,�`ߝC%�}=V3�3iR��c���F�����탴�o��2&jx�'*{�=yi(p]��u�8?�pb΂�3	�c� _F���Caqw]��ʻ�`�W:	`<}��b�m����~�g��$<��vYh��ǫUMi�k:�im�	K!��A�m&���F�q9���1Y�:�V���u(���4r��F�����ćE�c1�h��-������D��N�-��×ɍw��!�Bp� J\SJ?4�=Fts�w��ux HT��"�5�i���3#�4�y���Q�Ne|�����'U��B�J�i�JzI,�g���)�hv�'��J&���/�,aQG��>�� ĩ�F���a�+�l�5��BFHz�sjq|;�`9�
ǖ�����wS]SH���I$9����9Dor����"�r���=�������5�~6g^h�����ڄfz�A�= ��)�4+I�7eږ��)��wu-�K��ȕUP6��4-���%2�%k��H��W� ���Ǌ�gĿ���OI�a��4�x8��c��d�8����5�?$��:W	�������HZ ��G/H�� Yժ��0��,��$xh��UNFI�I�n����)s%�r���R���'��(J��X���L)��$�4:�A�%����F�v�20��>>泝b� VN�ǋ�ErU����4���YΥ��X����O.�tQ����+��ϖ��]��l2�m�s-IW�ډm"n��Uy0��S0��Y���(7����/a����{��0���ͦyI���JT:_�S��L#�c���� mlG����6�q�E�����J�x$���p��E�{è��tG ����,e�Y����|��q�\��N�����FJ���(K�l�Yk*
S+�~�<�R����:\����r�Y�Û*
�y]��ܨX-�B;�.8��@��`H#kuV�F!�M�m�G�K�}:�>U봮�6��	��tX�|_4���l,�l��j����J�QJ�f�S'�Ң��vT�1��x�J�� L����A�'���y��=��@t|ԃ6���cM���CtƖI�\
ԱC�%SȪ�n]4�c&ܢ�d4��콩ܓB���8�09�x��f�H��K U��!��@j�t�)����K��+q�`�տ8`@�x��)��-A�ϯ@Β&@�+���^��s�4/\Z��G�}�8�,�)n��B�!������5]HY�BE��mF8��"_?�� %�Ru�$vg��o�~�4h��Fo�]���L������_9�m�=�1C\�A�$�^�S��,i��v��1*ͰY�L���R�]VK��Y\�a����	�Xߐ�+��"Oq؛�}��)훾l�@S�n�3��Ѯ�݈ZI�4?��l���p��.�#f�9�55J�*��RTS'o����㏊u'�*v��MP$ԗ���Y�E����%t���!�g���pOst���g�}� s�����r	V��4t��J��u M��]wF�����.˲��wK����u���4L]f�;�|?�(g(,+��5�n@�}�Ή\a���R��uAF�ol���(H�A�
�b��&>Z�{��Q,*�t�W*��"THoӘ�t\��-�5��4����yBp1Zِ��-�DI")Л��F��f��5��m�o�/�S�cɉ~&jy7���C&�	����%�ͺ�8Z5����S�\�L'L)T����=��!����Uh4pD�(�|�h詣tnNڢ��o���dA%��+�R��&ZX^�n��B�Ӣ!k�Ub!����G5kc��*����c���>�l^uz��M#����M�y�O]o���'Q��<`�Ů.T]�����`�ô��9������Ԕ��qI�Nk���R"?m���`y�h�
D��o�~�r���i���_��`=ġ�)��PVx�!#{�[L�T�.�	56�Ȇ���o�ӎ��v��6����<o�Bl	�����)���n�y7=�	�W�z�o[Ń$A՜�n��$�e�)i�u���ĝ<ebU�`�T �}cd�����/���{P���$FOS�K�9Lq=Z���Pm��P�ѣ={��R�ܶ��:�t�pN��5*xMʏ��Q��ON_�k�K�8������'��� �"pW�J�1v�)ԝU	��K���6��M���Y�O�nK���X��F��1�/척}��$L��z�/atM�I(�r�Uy�Z㛜�	����j�j���r���fˠa�����{�Q��#��&����������[�C��g	C&@�v�E���1��ԥ�v�C��c��q$������	(�c{�ob�<$ +��Mjqt9l-�$�b�Cr��|��EM�BhG#υ'��W�
��K٬��sY�r�̽��'��w�饥rʖ���?���s����a�p$� IM]����w�t����w�W��O�h��^��@���	~)��d�� B��㬂ASf,*��Oq�d� �v����6o@�������{��Cf�Hڷ�Ì:�0-�m|1bJ�������T,C`(ÎK"Ӧ�k�8���(�����}�6��5@�d�5�M`� T�m�R%܌���oiT>2%�p礽O����LS�ƿbSa]Ln u!S���I�l�˟^XU�[�3!��H���@Aղ�+�5v���7���&�sB<��ގj���� �\<�#��P�6dt~��|��R��A��G