��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0�H�0q|x�F�Z,2�6���̘7ш�)�7{<j/){��]o��C���ػ���y��?��ȃCb1�UB� Zv�/}r䈜��p95q;}�l/!�<FuNF�tr\�\:��/�i�$c���'X�D����;��V����sc�sۀ�K��6�1�{�citW�RjQ�mݧJ�K VV��D߸8ЬJ�q�}:z�X�k���]�K[���L��7�T)	:����n�b6��c��Z�?Z4�=��X�����\` ���U����Q������|�dSDks,#���6���5q�l���AQ;�JA�(�eoP����)a�m���2���'��[�!����*b��W����$ QO}�������O�Y|�D
�N��<�8�B;8�"Ksc�Eb%[��Xi��
."/�u�4l����������3v��ӎPuom� xA �x��猃���b�q2ٹ�,�wt��ܷ0'�j݅�	״�l��y��)�r,3aq�����ކ���M�Ns����$���n��F΁iq�xi��}jeH�4��ÊREO�J&�;%�%�aOȋ?�.�k�E
U���kh�ZB4�$S����zv_<�{�X[h5=�͓�,�,t��P5�/�%v�� ��0��L~�� L��0sX�_��7BN�a%�p�T�%��x�_g��'0��^_�X�1�������1���o	NU��_��f�z�B8�z"���t�C����TArof�z`[����h���Al�/>�/j�br-e���P��D-�.�P���b���ӧ�d�HN)�#5�=5���x���ta4N�ch�ãr_�zJ�n%9gW�}>)�(V�A4��v���>��l�Ɠ�X���}w���ԕ�^�,�����:�7/PN���"ڞ}�'`| ���ݝ������ ��PA,�<�8��y-�=H�٢
^-�bt��꠭\:��(��v��B�e�F	����̹�2+��u�O�B�Bd،���Gv���֥�<A��Ed��&pu��ߎJ�F~�d�a���E��*���ީյB
&�V`�]11ԄD��zH>Q���^w;k�x:k=���[�?x�3G��$�u��P�s�&D���X�a��DiW��E���)�tJ�w�nL��7rN�����������`/��,Jm�5�uG1g��$��,��>(Z�\[8���ZS��}�k6;C�J�7�����g���@��K�'� U���	���!�m�D����ԫf�d�;[&�r�j�6ݶ>wJ4����Ӳ�N�b(#N�՗�<�?�%�ޞ^��.]�~Z���Q��$��i����B�����'iv����Kid&��uSzV���?���MGK8j@1�z5�N[@TV���I���~�[�&�j�j�Fq*'��ͣ&�)��V2�-��Kϟ��b�Q��e���JU����	�U�����
���X��m�=jR�q{M<Ն1�g�O���%���U���B�e�P�`}�� �#4���_o�Z-qU��[���=n#�J���$F8 �f�bQ��>�j�R�E~�����a�,<��ͩ�Rత�
(�(��E�
i1�70̆O������e�'g�N�� =u] �S;���^�n�꿩^����c�>�^��F���sA`�4aX��G�M�^������[�u�0<R��6���l���2iQV�2�}v |_� �Io7e�_�Q�jk��j���At��k����b���$��9\�>�}�����^#�݂_��.��3̦���%��M������Sy2$	І���>Bul�>1N1���yh�V�_ފZ	�E�S����I#���T�f�;	X󍒣[ȹk�x}����>P�OP��O�nMf�=��އs0��6eQ�d� �2i��o  f��� ]k��1�Kˌ,%T���&��g���  Rg�B�.Q^�;��a\� 4,�pR�@(Y�ڕĻ0�p=7��]�p[t(u�(.;t�-g�fP��)T��:�����6�zČ(�(f�ߖ'�d�I��DZ����p�Wr�!�K:=��v�){��2��|E'�/����7�l�dN
2O,9f�WFG��9l�*���N�����L�4�s�����,�X�A������"y�hZ����Y���</�\�b�Rs�~@rG�}#K%���Rd���im/�1�?5p���I'��fCޕ��j�V��2�K�N����}�}�¾��nQ3�1O`1�;�uzW�2����!���e�̤z���ʥ)�[�s���۫lg��Dy��W�nb����Dl�#ƻ��(0�Ң�)Gܩ�?2��x���ٽ�l��(15zK	����:	q��Ȣ���e#CU1b�i��={^,�R�]H8s�KC�xʏ����t`�I��+[v���ӯ��s-K���ٵ.4��ð�sM9�z���O�:�"��q��W��B���NO�(,=�5ޛ/ sg�4����]��<7�T�,��p����t�+I!�Q��!���Z�!�U(�"1�^t�5�5
�ʇ'�;����DȐ�/-|#C��d
0��'*87��H��xy�7?��%����h��`�_�V�b�蟲���)��S����Y�M��y����^����b��V�Z��9�L��=)!o��w�	�r�]QŻ��5ʮ�����v�����|�;Y	y��s1s�
������!�%(0J욱Q��&��hBj\:wN:����q��Xk��Q#��XPm���Wb)=��U��"q{�X̲�<���lw�I(�r��ͤ��H�:��%��b�Q�}Ǳ> ��f/��t�F�}%"�r�Aʀ�� d���NnI �>v�X����Y3hC` �0�#6z�i���CYq�ܪ��а�f�C���BIP��e���,��Oo�oV�f4u��J2�B�x��X����7BH�����޳��3�!^�ka���4ܩ�zR��lq�P;	P�s�����͗O�V;�A�RI�^�7���5s��K��,�
k����l�+m5S��yUO5K^@�$^�ּ��g�.�
���F��4Y%6���VQ�pn�'����T��%���H�U�r�����$,������\X
&��f����L7~��p�j<��M^�9*����?t�\Ň�Z��J<����c̃foz������@7���ze.p�������?�w�U��w͓�
�Q��N� �S�t������Ų ���������_��o��ۺ�Z���Vߵ�?{o\��
���@-�߃�	��"W��Ē���Y���=�����`�.��F:� ��ᝌ�h�1KHӳ^��E�r}߳��Y��}�m��>�/(��w !MIu��RN��tc0��Z��2���sY�u騥�t����������YJ�ae�w��*PC�����5~f'�����!�
Y���GI9��$6d��^�z1��kpAX��社[�ۡ+������*���n�|ԓ���@|0�h^�	��X,jbv��Г��6�y�i�¿�dg|%��S>��6}t�� �ZZ:��4/���L��:����{�:È}%w��Z؉��cDI9�=P^��֘ M(}�8��B�e�@`°����A��j9�U��1����r����fuY��ᔓ�C�:�w��
����6��/߽ƃ'����Zs�#�������y.^�!�E ��)�g��PkZO���m�8�Ą7'I�y��Sk�`�/>T$n�P�JԜ�\{f3E�o�����[��sv}h�ǅ�;2���`w1�%su���w�q�#�����~��u���&�ϪHsK����ш�� �+}�k�v!�ٍ��#gP` W�&�rP�K#�n�!h>�v.��O@���%�RR�-��'�'8�4n���-�/�QDdM@��g��0��8v��;�}���zy�xQU��9��I P��͖�Q���`��]�f�!����s�N��	���,/~�T���SI���,1���QT��X��ޗ�Es�w��;~x�PP��뷐�H��5G
���dm�X�<ޡ:�0���=ڮ�rʉ��YV|� �A[c��{��2}�7��b��_�h�&�4Lg��r�ށ���]��g4M.{nIy�N��@4l7���s�u_K����`
�A�x+��h|w��%��s� z�{�l.៵�x�9E-���	EʑJ{���q�(2򪵨��;O��9���%��TS�v�����rW1$	��x�@�����AS��Xܮ�hf�n�f�3ao$��i��C�7�r<�$8JÏnJ�v�Ԟ^��/�CO����ʺ��=�S�/(���s��������kz�#�׷�%d�8�8��	���Cނ%��?R�v�;��@%g�w�{+)x{M����"˼��Q��ܘf�Z
^�
�}����Pf�XN��}�x�+����(����%��R�J���f��2���{3%��q��~��+�$����R���7�Fp��B�2	�4xd nyƘӺ4V�]��ʋI;���Q'X^`P���e8�FQ2A���Z�$T�E�f�[~) ��W�$�F�x�� ���ٖy.���z�e�ʜ�8����a��4�Z8�3����z\h����'ޞ?T����,�^��?"�7c֮A��IƄ��<T��=�,4��g�v�J��/	�����B���#6�eϭ/��ʅ��f"d���v蟟�Ci����[�& ��*�Ҳ��2|��rֹ͉S	]w����z)���?~�%(=�0Ku{����s��`���eeK��hsa��vO�&"Ǒ;u�>7�H(� �������1�Y���������
�����&�%pY~x2��+��%���[�
s�Q��������C��V��N�L�R_�$�˚��A�ȑe[���tY$�=���m����%�ҧϺ�g�̎�VҞ��^8ڴ�s�Vb� ���~��a�qw�=�lU�<�E�rf��2�,˝�-j7IX�I+�CQQ���ՉկD�A�����7Һ���:Ta_:[[.�R�FI?q$�4Z\�\���tT�����B[�5;��BS�~��E��ݕ�Ψ5'���fN�G�@�V�R��~ �l�?�&�?T��)��'Q4fv��7I�k�;���3�YAahK���پi�� G"#ڟU���F���_�wC�r��7��h	�o¼�A6�dNy��D���H��Z�$
��nVp�_��ZSnΫ	@Z�W�״�Ĵ��Pǁ�Q��Le7X�W&s�����N�U*��3�E��(���Md���t($�)^��W�)�8�������&"4�[�d��ɰu�#���$���b'���}�Al�On2冽4�'�>�'�&�}�Y�\�#�)9.�]r�đ�V=0�O(������ޕ?���*j�q�K��=s!���ѰW����A���Y.6<�-��6��2�/ ��7�s����b���L_*�����ZD�8~�*��=���"����#�oS��t�*!�0���Ss�W9�����)"g���	����X�J�.�i��`?]i���&�𑒫����φ>�X���gU;Z�S�=y��7,��JT�S�GՄ��g��-m��s+,��59�gڼlӟ8����i��t5��Ѿ8�;��{љ�׈�x�9�KA�/�9����i'�#m�M0��'-{������R7{}goJ����a�qN�}͘q1�����핽,�fB�gZ4�Xj��mT6W���9\PxE��Cǲ�öb�Z�&iZB�n��#l3���3|h����:;��Ǵ�뻲��^[s�oΦ��[/�ny��:��a�D]��S"��2�J�J]�ۖ�C� k�^��1��pr(g���N���6�v�;	a�͒'Fq��_H�>��OÊ	�/:��v�-U��F�b���/%���C��y��M|�wK�������Q"�i���A^4�����G�T�m{��BG�\����˫J��c\YmV�@A-�:q��X#��!�p��:��l�3��Ī�V7|�_�����d�º�g>�5F��f ���Y� ��s�V��g�H�Ʀ��AT�ΐ<T�]�w�)�s����ɺ���s����3Tn/���=n���67�{�BT7�r:�𜆞��˵����au�L!�Of��ȨLVӛ��>wY�����6ǵ,���v�Y`�|`L���Dh�H�l��w.�Ez]w�D^�B��z�j�[�"e�r�	�d��z�W�������Z
!�������u�U�eV����Hh[^����g]��$�s�u�7>�13��K�����z��֋��J�`�!�����؞?r<Ť`�E?�����	2R�j��#���lk1U��t��v)��ܝ��S���ym��?�3.'M�
���%\3���I\%��m�Vi_��R�ҋ�4����n��+?ADi
��À1���772�|�i�U+����{��h�/Ѩ�=�)���/�ԣ�.�_���TԹ^n��v����SM7��	��07P�匟g��x�"HBbNm�Va�g��?'ldI���f���i�X		JX'Ay�GD�n
�������/��mvH.�np#��v�:|�`��<S?��C���B���dI�bcUP����HxDY��<{�s+M�O�zkP�����w HbF%�'��˕�66
V;�r	o��g��ܵ��`��Ő��+R?��F�5�jG:��o�G��Ii�џpCQ\�~51u:{�����m|m����L��frK�=J�!G�f�o �d�Le�N���*��o�G#��3�!�W�K�J)���qy#M�����H+U7�7���p������N�����(R�?Ҡs��8���7U訮�s���`��R�.������ѧ��3p�T�`����R��^��>1���pBtzC�A�?��X{� �r
x2���	�@��q�G7nY�M��^9������ad(��q���� �Y�㗏t�L3��q�/����S�a�ٟ{S,9t��,M�#�q��M"Js�P��ɷ�kaf����o�Ʊ׌P��w�*M_��7����ov��@d�8�z2����9�3[)7�[cի(�~A��0�]I�w���\��	.�զ���ع�>LT�feIz+���Þ����`_. �_��5�kR����2ѡ�_(�	��w׬"����B����!>�֯Mg��$�L�6����Pў�]m�o������ԝ>`�Y��"�\��|�WH�s���+ͦ�����*���m������[B'���y�1z��CX�+��kS����>߻������A�v���`!_���{��֒[��.6���.y�I�8FM����jc�� /9Ƞ�uȘ�X���k3�U��b����;��%�ڗZl���k�{�~���tC��i���w
f
���nA����v���5��	yw(?5p�7V�q�$l[�c&���HLT_]����\mU��{�|)v�؄m�w���3<�C�M�#'��Q-�`V���d+��1vX�W�ny����=Q��;�ta��(^W���y�ד~�o��O1}���1��<?�����x0hE���T�)֠�FV�9�wĖx���6l����l	F����ڋ�s�f�w�7��x��	�����Z�����P��I�׎ �X8t��A����_���_B/�N��)�a`��ɶ�뺺;����Q�������̐Xny� H�2۶j�h����,3�X�aUN��v��ظ����(q�nK�R���W<(�ҕ2��u�ʈR[>�1@J	r���?Ԝ�M�z\.���x�z$��P�u��Y��<Cq��ޢ�����2T�R�V0�{�M˴u�vy��0�Iq߲Qۗ�f�=:�����xN
9G$����4��*m�_(���Jx��ְ/+Z[��3)��e|��0b�\8�zZ�TL��m���O�D�d�&��}�9�lP|y�E�>���ޮ��Snb�e�k"r�LE��)�6��W��_m_*%�Ԧ�~c��7��F�M��S��� ���"L.?6G�âv�x�5��L�a3��It�f�������~�m�Ŝt@4�gNx�k5>���P��L$�)���ER}��sHUt��X����6_��
ζ����0+���?F^5�4[=vg̙D$M(@c������x���1��P݁�t���U2�����:�u�{���tܴ}�}}�ɔ���%À0r�����w/u&��b��Tê��/9��T�G�!(�n"XD�_ñ}�k�Lyɰ�&Q\�@����b~g�A1h���jH�e�+amň=+텏��I2�Ck8��,�;�tLUWl�!U��0�������$���+�@�kGl��$�?��Ǖ�]q�a� cU��]�)����5������L]Q����2��g��o������t}�%�������O�[Z�_����u����|o�:L�� �� 6� ~��i�>g}�!m�5�,߭:�KE�id>sBH����O�o�_�/���F����p�r�i�Q