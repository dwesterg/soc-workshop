��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��/E���3Vʅ�����v���p��A�̠m}������"�|7g�f 9�����9y�ކ�������M�罘O�{j[_Qg>�1�89Q��v4ac�ʋ�Ȍ�b\8����W������K����R����s��i�vrr���ܴ�<%5�s'Y�G�ӣ>�$s����
�נ��{�%&����d����m�kB8^9�ҏ��R�nL'qn4N_�����l�C��l����l�J�>�Qv���|V y�e��݇�ъ%�=!; $K�/Q�]w��{�<�r�$fC�=&	��@DKd� ̮wu:�o��4��w1���/�}*f����W��c^�
�����.�Su�;��
e�V�8�ַx���	&���t5��a����܈)�e%ˬ�F+�G��O��"|W1X/=Xt؁����x;(k��+r����r�9/n=��i��=,�9��0q��f��V�,�ң��x��YY���@��(b�@���'��G`�>�#�o�.&S��E#�2B����ad�-X�@�Z�Z*���?u���_@�gv!�����K��(k%��znDs:3�4��rll�Ng�����T;�����ls��a��I����c� �����E�`�y�Y^�^��i7IsTF"H���:��E)b�VR���'ݍ�l�e{��Ѕ)N)>�Z� ȥ�����K����ypʫ06�Z��	� �������Bss=m�[[KB4H�dAY��;��C�J�Cf'	@�<�刻� 5n��ۅ��	j��H���L.W�OI��rv�)w���Iٸ2���>>W�\�{�O|��8l�D�"�i��Ȥf�J%���9%DBF��0���{�][�ܩ�]�s� H�r��G{�/�]:��:�艩�zH����'��
C�7h>�K������J0uv����.��GS��RHOJoQ���$�R���>^G� P%/�Π,��Xu�$��Q�ͫ��G�̂��Ow
Ƚ�ـ.��Ta��Ng�x���W}7�Tp����F[bM��ӇƓ�K�����k���R������!���L�u�hB����q^b?#�X$���u��X�#{��^h��\9h ],zd��Py��u�#z�v�(q�@C¤5>�Fܳ��Q� T3�jcM�� #̕�%HQ�o�Yݵ]TA�����plvUl}FH������Tի�J��ij���h;\��`Oɵ�N`܂�Dx��SZ�����y�!�tP�,�由p��s��6�G�z3�;Z��3���$�%�,�n��3�R���O�fp-ڱ�b,=Aos��r��v�Ƞ�z����R�����h9_��0�9�Ş��1�eTM_�9ξV��TC��Ko5�Q�lN**!}���k�^q�l�Y�UXU0����Nq��Z��'�U�>�"�do�ލQ����`p�]9]ьKNi����JlF�������k�� <�&B�� �4�ǠLkp��݋ٖS��3��q0���*��9|o��a&���ۨ���QJ��Shl�H�X�z5Fl�!'�x�P���p�bĢQ,ȸ��d��*T?
���1Hc~w���Y�EԽ�ONNOV�����x(��N�����JUl�>�_�}rRD�J�m��Vq�m��T�lGE[I!L��0���g!�Φ������Ċ�N��Ż��Y~�]�(���9��2+�q�F�V�	
s+ ��܋�~�a�����þ�P������ִ(=�0-=CEd#�AƧ>�4���^�`^�uh������*DWd^�ݫX�������۵]�i��e���P�v��j� h��?���c$,MG�?�h�%�M��Mޥ��IAa�*�Y�7������
a�d#@'�f�=-�d�#n~Ny���Z���#�Ã�Fo��5C�}n6��~n�2��z��lM;�͇���5G�n�I9!i	����B��YZYd@u�N�f*D��q�i%$�Ƴ4�LZMr�wL�����h� !s�u�vH���ɔ��o.1b+e���jY!B��a��/�U�uz�V���&
[t�DHd���i y�Q	��_�0?�g�w_,�«G{Cl�c���[��y����	��Z��X�]����!4��a|�5���OH
���4���b�|�"����X�ȍ�=�ͥu����r��}�v�b[�����S��9뻦Ӛ��������^�X��C��N��CH��#\���W9D�o�d2�6�0����5v�C��a�z��ro�qaY���^�������-�Q)�m����]N�e&͈�����Η��t�*I#[�p..�P��*u4S�d����a(�Ӑ�Pŕ�����0��i^��"��tJSľ�'ExψB������P��*��s�֎�Jҡ�����0�v;�v�^�Ig��aߺ�������<���v5��E����y�֫&��Bu	uBc��]#@f��
2$��}��a��	�s��}ö���e��!���=�R�v-� �_+�C��р5,�����~����S��{�E��%�m���R����V�y~��_d4ٺq��h��z��j�=��d�P#���^�z�I�<���VT�q���#���+F�x�2��$�i=�0m�:�H@��W�}h��O>���P�;+3�J�.�/Hn>�6�'kɄ,���*�ԋ�l��������&����_�J��i��UաH*�J��zh�v-�Biޏ��Fr]	��?�=��K2f:ـ�М��������t�CP���J�w�ͧ]�*����+�d4��SW���6u/������ƾ��uȒ�s�2�0sb�0ߏ�
ώ*����2�s��)|N/D�L�!i�P"N��Cm���2�|roZ�}��k�n#���1�5ɐ Y���(�0Y����RL�tE�9�K�k�"A�q66��j�>�4�"�z�{�t6�_��T�s���Q��t@?POз;!E�+[<ʇ�d^�$b���A	�u�}��P�^~�.-�pT+�%c�V��>�Y�\������$d�����ye�}�B�����=�$��?Nlj�+`"��{�_�f�Q<z�hD�����UPiKeaӵY�2̮��.7ݲDV&���1��h�h�Xx�w4�zv$H	!Wr��ܫҷ5>�#cıUy,����8���L<(��]7�|;�̞�!Vѿж��Sjs[�<v�����6��C�xV� ��5��Ľ����I�j�
.��2����k�2�[d��2{���l������`�gqQs��OL���XN���1�mw����t~��>I���~�� �j2;&���9���o� Gy^�����M��ގ
��&8��KW�`"?�D--:��u�ᤳ�Ol݈kV`��Nwu)�u��������]�B��r��_�����f��O�*��nBg�ft�@uY������u5h~@�yy��B�?�Np�m�f20�i�c�׋ ��U:j��8VB� =PŁ��9�Y2���`]{���~����q�����I��߀
S�E�;�r�C��������l���J�0�)��n�w�+b9��mY��A�i�J�J��"�v�A��G����W�������,�%0�O��V��2V��U�*ܦZ8~Rpu8,c�λ�j�k��+�ĕ��#��f{�v>�}�G�q�3�L�ʗuV��٭�4�L:�i7�Rڷ.O�e�kO/ߦa
�'#ހ*x~�<�`�Ʌλ$�I �AN��t���2�ܶ�S����a��r����kwɓ�E����C��p:�'�]+9�J�U<�U^��wwr��\�g"��y���R��:XȤ�O��5��i�xaw�	 ×3o_8�H��U��������\e�J��N�V���@nٹs�B���L��W_ʔ�ܒ��2'�Vp�u=E�\�Pe~k��Ij�d.�c�#�	��5 �����3"���ܤ�P���,�}�v?�$��̡@I</���_�&��#~ʴA�~o���h�����n"��U�!�Y���&�>����������/Jt�$�*�@<m�! �`IHD"���}|��}X�Jy]�ʩ�w��\�4�?�0 ��!����_������r`~�Ju��7���V}��Py}�Qm^������L���k��@O�` "~��5�6cD/]�P m���`�ڜ������R��1�pH�����Ʋ�r�����e厡�>��Q �өI��B7'(�혵,ڏnO�,0US�e����$��Ck�z=���vSޏe�Y�� W�E�6=�naF<��߈��oEAQ��jw�p�āk4µF�{f�L��HW�Զ�9�$~hdJ"�h�x�?�c�j�����$��{W�',�*����=9�< �����8*�^�B��쐧�.�)b��ƈ��ʃ���W��ظ���n�{�SœN!t[��IA�H�K���
`<x@�A��~�I���Ժd�@6Q�x�>C��G���W��K�}{�[:�ǶK|�����b�y��1i0V�1�x&;(�yT�K��Qi�r���޸V���7�7 7�ɪ.�z�S�{hձ�>]���7�>��c����]w��
E���e�)��eZ�;���&!����4D3ޥ�+^o"߿���~��7�)RF5���׵Ds���V8���E�?$��]�&���\Ҹd���[Է>:�e��ؐ��hu�	l\���"�/����u	·&|����*�Q�������[��y{2?�}�����v%��ihs�6�rT�/��^�`�жۮ���,�%QF6�A�q.��Zu��r�yЧ�0�K�qZ��xd��PT�� 0Z�ٗ�^�y��Ыݬo|�b|�؋H��(���aA-����Wt	�U�����7�w�0�X�o4��H���X�N�h���@סIc�L���3B�^^Sn�>`���]hG�!U�K��WM���Z�9k��k�&T��ՀN©�JyCQ�lY3����u�<�#�ƥ����^�\��Ð��l��,��B�'e��O��r��5���*+߰6��nZ��6ܸ�m`��@�������pk �`�S�:1��>�����x�Y$�1I�
��:�*�?:_����P8C�/X��]�-,)��L�H�r��<u�0�w�1�����mh�L��g���
�}'\�X{��$��2�Lۭ�����Oz�[�t��9Tn�}�W��Ni@��fl�_b�"���S�\VE�⋏�p<r���䂕���;�v@�|��jtǲ��'k��(fG���&f����ļ�డ�g���z�~^��m�L�'m9f�v&iuJ�'��sm�Z�y]"g���e�?_Wl��EȈxsqBy�	0��s�V��Q��A[p��8�
~��(ڄ��>VG�t	6�:b��-���:����'Ԥ�{>�@u+k�|�Ę��2���d)BX�`�&!
��߶�P)[@]|�dњ��i�i�n�Q��
�U��lN�^1��ߛR��Y߉�U����{��Mָ�K��K`�����|XdPõ��� �-<�/:w�Ұ��-e .�h�NhJ������1W�_�fK>��ܑ	Q��F!~��L���6A-�4�4z�Z��E��00��Ю}��}�0{A��MDD���!��~��'�R�
{ɀ�����0X�w��}��W&� e�̀*9�C�y��ͥ����$���ia)�~���(�e��j[�X��ŵ���G�E�	I
��η�쯓\�l�\��5�w>G��T�&�H�x>Js�;��v���<���G|�<�R�.�Tz��&��7��}Mk�ykxj-%�9_���J"�ǘ�**�Դ��=�I��L��V$�(�M{E�Л�e�H�0�����w��kg�\�w��~6������Mϟ�+��_@�[�~Okz	��'�d�}bE��	y��a����U���w#�	Lӳ0��rC������p�/�����#�b�v!}�_�u��=V��AT����J��=��F����-��^�4ě�;�Ӌs���#\}����KJ\^�j=��s�x킢>T�.c�2<[���rZ7�W�NX�Ty���J�B�"H�$p׿t�f̶b�]�[�ߵ��{xh7f��'X �h�'�( B׃v6��OOii��]J4�����z�s1��a@y|�^yX�D߂m<p�6�f؏&��K��I}|Ѣ~Т�Gf�^Y���^wm��w���2\9|M�^��B�8;%�*������6j��\����P�3�4Vp�cQ	z��2E���ٟ���&,�8��V+V���:C�-����ɧ,_J)��:��)2No�����]����F+Z��Eh�SrxT2��B2�%�;������Z�CY��W�"�Ç��5+� ��+�����}�$�#�e��^'��	�Y��;�5%@_e���n8ɟ�`▀�Ŋ�[�(ɳ>ǁ�J3A��l�#$Jk!����n��x�Pc���Uee\��7~|Ey0p��L�!�*���y����~������UZL�Z�%��;������8sI�W�}rq+��k��������pC�;�8Gk�#mL�q:�d�f�[P�)�x�V_�] ]lQ���ѡr��f9;B0Z���9�������=L���hp�����S��^L�Z���/��4>9F3Gp"P��"���O��*K0�3-q��	�	��/�ѥ=9s7p�`¢�-�g�G�i�ImH�Q�V3P�5Qȃ�x	�Q���I�T��H|y��~�$�˞ �G2� ���p
���y�z��O�Kk�c��p�O�Z�\��G?F�l�@c�8xJ,#h��{&f���&=ҙ��r'�|�mf�W�{�zay��	m��/�P�O�[��(1�nc�j!IYF�d�$��1����q�p��H0-M�P8��;�+�jZ�T 6�_���}����;/ܭ$���v$��fc<�-S-��3���N9w��sJD:�/������W�x� ���)���
R��k�a��T��HV�?��v���~S6m
:jgz�hͣ�FR����t	7n�^�<�O8"���J��SYl�f\����r[�G;)���ш�ӿ���~RYB�Ǘ���_�ks0@M�8u����+�R��^/�0-���}Ą�ϵ�D�"Q�'e�	�������1 Pyl7b��IX��2�/��	���R�_�G>�ޔO�J��0�L��U?�q��]V)�s�͊m�n����R|���h�^��ؔ�
&ɂZX\��w��1Mi��3i��]������N��yScnE�DΎ[@��UZ���&���-�ie5��R�h޻s������݈c�R~�b\�	U��vI�7:��Ⱥ��X����v��d9�P�7��
��� �ޱF�3Z��z���D\�b\�cM��#���b�H.��$��)u���������zM���u�9�x�
�
���u�p%�}4hm��8:�.�vG�Q?}�L%�"0.i�t/���	�KX/P�N�i��{���e��-h���m�l��+#h*�?�E�M0��q"ͩ�3�r��[�z���9�2����C����w��Z�ux|+�.�����ChS�n ��}ZTg`��JR�4Rd �����J�͐<D0�u�;��}V����no���FC�~F.(�5���t���3Ɨx�_�� ���y��)�W�/�y�s��8�I�
�_���a|k�zW�e\)y�-���_�H��F�%�����6�
�k�����$�Z�]���0:1�+*e��p ��1Gn�s���n���y�K�#U�/4��o��b���0?��x�]�C�q�^�� �����9Ւ��	
a�a�Ɛ�"��dƹ�;_c�ո�����]��(���U#�u��F1T�K�^��P�y��?2�lmﾰ��>��;b��Ѓ�2so�=�6zC��-�p.4OJ,�	d1�Ԃy8-]�
�~^t��O�w����sN����揋�Mfx����(�g��c��ɴ1�?7�_ �Ֆ�.��?O�I��A��fD������@G��#4oH��`�.`���NhKg�+�+:��d��1T6������6�{�����B�S�k����C��dw��ۡ�����PK��{-U�vokQ�τ���`R�J�`gl��yl$�PI�)��\�^���5��<0����p�m�z��F9G��e�%�����P�Sb3��gQHD��(D����l��H����;��f����dm,�ڣ��pI4V�i �~(���>��=�:<!��´�f߷�pg��@V<�I��Bʛ	�s5��_�k�m U��;:��=
�U����^������5F��G�������Z�����1Bc� ���~�R��l����i��6)4ȕ�"�d�P�E�z:i�^����٠ۍ#��x��K}^ꃺ	�z5�S�c��r�u ��:��썪�g���t��&�1%�~��$�	��������㊻��a�fbk᬴�9�-?"!�t���p��[ܯ��E��R���%W&�4Xi`�W�_Z���Kה��"4�X���9����$u�Ts�7iI�1�G@�Sҭ�Md_���� g
C��:���� �!��w���l��A�������L_��������x�������h���P
�J�{?��$u>��&i�҈lI��	��Eg��1�;�(#j�v�&��v=ȗ�W��%���w"�O�*�{��I_�� X���t�Ej�F�q�]P��@x���e:����x����	tơ��0B��~:�6 ��AK�`�۶J J�kc8(�/ ��&��l�r���e+����B"�=S:1_����>����)DyQ��|:T��UlZ�����P�بIb��ssMN�e&��O�J�����:����A��s��%Q�dg�y�I�Q�%VA�����h�+"D+�!���!Rw��atM��	�5��y�/ �fb��V|�f�@��$�>e�I�1�P�@�
k��Y*aQ����c8��OC��F[�5����)����� �ɜ�K@/a��8'���^D���uR}v"3G�Fcƕ�ǿ���e�a��o�Ϲ�ڽ�:�ӥ�)f�Ə�;S��b�Zy��̴���o�w�S>��oDg6��f�����aG{Lφy�e��mf�؅9d~��F�4RR�e`8	�z.����[���E�����c�6���(�Cb7X�jg�x��iVv7���݇�S�r���Q��-9�F�D�;h��#d�ɉGsE���~P�.�n��#�^mל
@G��W��w(A�*IU3sm�^��L�,�'n��B4n�CP�����Y��Ӊ�J�����'e(�ܩ�wI	B�ơ�aH�Qd�f�0�˚]���ޮn;����0@�4zi��
gC?��:�2X<a{�z��p�lǰz�����" X��|8����Qw _^�N�	:�w϶�E�}��${��;2���1_�~����H;p��6o5�i��=�I���k�������4�W^ol��W�B�yE	[�G��*��!iΈ�_ G�"�j���ex);1���+�k�x{�0�ת���=`8�w.�����m�6�U�����~*0%\��vr���z$�N0ЬXo�$�N(�)�mZ֚�G������嶓��� �fu�6���:ҡ��G�k�^����x7�u�&Kk"�Wr��P�K�m�{��g�t{�a�����_��j�طk�x�:�`����� ������/Y�&-���!�z��]�P��(��W���R���=1�����>1�>g$���pUE�^`���qgn���.�y��-$cHN�[\Vnc�C��yK���*�e�X*e}��X
�Y�+/cX��xG�b�Y�z%^���׃��=X%��o�M��VQSG�ԏ��j���C�j������D�Z��������$�c��w\�b�Axt�j�xV��.���H�����܋ghr	 �?)[)��:���j#���^�6�t�����Vi���I2�_�B?6,уNQS��gl%��!ɷ��p�H@�Ϸ�#�;�R�3��u �}_!ˢ���e��|��5+.۳�S�N�����w^n��VA�����~\�I�=�7U#��+ir���t���%Ć��K2��+Do:���}f����^A��ŝ*4� X+�����i_0oBѸV�Xo�]V�K|��ru:���C�n���%g�#�ջ�\��x��*
���.�{��!l��t�_�6|���ba��G��N\$S��N����y����	��A@bS{9�%�����?��m��]y�laRt����7y<�NZ�����G��& ��{��6�
��"��Z��_xڙM�A���2��-�ӜtJ�����F�ܕ2Q*���{����O��
B]�f�K����z@T�.�?����'�O�Vn4��o����S(O�T��4k֗���?��8��vGR>[yf�mנ�!���x���rĐ��*g�Mqb+;��dV(��d=�t�wz�2���;l�&����܀ɭ^�@�����d��mA�3 ܩIC�um�h�β�����Uឣ]���(T��ې	c��$�SG�*X ��x_�̵'ƴd� m�4a4�Q��ut�x�6��B*��h8O����Ug����a#��]5JQ07��ݛ؅��"$�R�R�y�Q� �q�Y��n$�R���V՜�}�*������;&C�v�,���[iCziz�S� �v+���ך�A��u��!����!buW�e���(��1����>��O���g #���P�)�8r=Wv�Ε&8l��LG�]""�^D�h�~)YF��x��q*Q;�@*�@@As�q�ߌ��0���2��y����Qޔ�F=�ª��[���d����\�|�T���SD�0K�,O����k۩���� 	e�?��a�\}vKT���}W��މ�3d@�;-��d#t�Oe�Ԍ�oz����)H���L���; ��+t$%hEy*�`熧Pʫ�2�q� ����~|�kE�Q���<��䩶.��[0�L���վD�L�P+� �;�?�����.N�T��,+$�I_��p���2�*y��B;���
S�D=)0�M,���̑��+i�?B�.U#O)�ݠKgx6Zzf��h��R�qH�AY�V.�=L�9#��`z~Oyn/|'ɣ)�7M|��u����ѽ��
ʾy���2�>?HnY)�hu� p�O6��Q'�>��-��Z��������nsϒ�-6{B�����C��*%�_7��Ћ�V�,����PC��[�/�Z� �0��g�$V	�� ,�������*� գ���[��׵��{aYl�6��l�=B'�?���0���-�A
���U�FzN���8+)Rl����B{a��}�ț����?���*���xgf��3Ś�]K�q��S�h�@a3�C���sX��i|wɾ���(xÒ��ݱ�~��h�@|��F���D�6�/��XDƊi?8R�6T���Yu�����q�E;c�:/̫�F%������#�����/H؜i�����1�\e�,Mw�_ �Q|��Z:��yYT���s�"��s�S!.S� % ��;�"h
�^��vZz���|@�zs�1�$�Y��IL�����R^��$}s�#���ۇ9a:S� ./�8��트&�/�ޤ�Kס�B�t�2����we��d���/���]F0G�Ea�3��L������
�ڨ:�g[� >]�2�y(�kB�^�Q�h���f�PM�&��Q͕��[T�*8�@��ǧ��-��x�(�ff��g��ź����=�X�&ّ'd	��
)������)΄���Jt>�.F���E���Oԝ�U[����T��N�6T��O$r���:Q��c��3*F��X}�����W�bQ��GP5�yJ���a�8{�f�6��8R:E��JΊ���Nc.��zS��͌�pہ�!�):΁"�;ÄC�w��t��)&�"C��I?ֱV�7�(;��Ȯ��	�-MQ�$V�/�Iԟv���:iZ�W��	���Ȫ@e1��sO�"�4л ���@�_�!v@R�o��<��5�qf�]\>�n@���^n�L��=0��c�T���z�y<�/���|����8�t�^f����Q�Ô�~�"?�o8I��j\�ٻy[y�4A[��7�5�Z�~�۾�=�r#�Ĕ�T9�Oj