��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd\R�̾s(��MI���C�X\ņ�Z��'U�������(��@d�	��3��o���]�$f����ܹIͮx'_�w���2���������S�9�VV��s�W�4i/J�!{Bɦ�ܘ�Z-����u�ys�}m�)D(|��R�=��G�E���	�+9��y�Δ7��f��w'�M&|�9K��ʑ�}mB����33��!C���t򹼛���Y��f�!ST���OwU�����8>7�9�({R+�M��qS�{�k����E�ӷ�c�j��yg���cRq�j�v���0�;n�' �N�%w>	�޲%�"��,�������@
�敡�
��ao�8KG�qE�| ؉ O(q^8}q�W��C�]�.�y ��;��:LG��%����x�xcTʝt��S+t������]�A��dP�}�-����r�{���U5��n��`���ù��r���\|H)άv���0Tz��y�DOŹ`�&�Tݿ��G� �ͮ���(�� D�LW�N��B`����LZ��@�ζd/br�Pe��0`$���rX�U��7r�� �!J�ɋ���#�U�ڕ�G�i�ik6�`�e��m�Q[y�v��,;�C
[ޠ;�Mt��rT���B���cy0j3�9T�Ely���P�E�3�41�ͳG���?���&Δj`��̗��i�O;���HE8q���ʣ?U�K�rD&I��`�[0@Y�͔�=F�/��/#�D���֥Fڊ��KE���_Đr��0�-��ztKR-3ˏ�ɩ�F<x~�-?-L%����(+�^}䱾>�v8\�bX�#��b�@l8��2�ff�Jn��hB63N�U,��7x�MR-<���^���]>�E�<�2�N���n$oD�)o�FC����,	�v�"�r�\b��x��z�R�/�S��I��|�x]3������x-�kL��,�$��J9TZ�@p��w��'�c�G;Q"V��*J�w���PD�m��r����z�I����`8%���6��X�n/`a��
�t���gg'x�DӾ�����M0D|~�'�1
�p�.����^m��)]r�|�仢]�L?�Ř^�?�ΐf���3�c��u��5�|���""?y�Z�y~��yI�q��|l-2�5Ўt�~� ;��R�j�h�!��3+��l�+aޛ��B�oQ�F&���AZw�Ftv�fgEִ��T�q�#eM�I�y#����ӒʇC�����v~�ݞ����z�7A~�,�i���$�L �����w���c���vE�� K�G��er���,�r�όX��p����RΌ�3��	�cyLp�� �Me;kn�I��NԊ��yN�:}+�o��,�BF�	����\��`���]$/�h�+�<����D�\`�G��B�Sb3�Y��0~L��-�m����h�O� YJ��8p��0��u7	���?bҪ@��-Ǽ��ɰ��~��1��{��:��i�s��T�t4�	
�)���V,H-�����rγ��$�c�2���(�gv�D��gAhNiJ�hN�N�E����$
0��Cc���|zj7���y�,,;�/a���,X�&��}�\��bv?,�p��#��@�y�{4Mړ*��Ҋ�)ШҷsRJG٧9y�d�@�4T
)g��`���AGLiw"?+f�J�-#�8�WYz����W8��T�z��t��Ig��&�U�a��3	ҙ¡>B,��/�-H4�O=�R�hg	6�8���U��B�R�^��Ԯ a�ڗQ��Ƚϕ���	|A��q�_�i�v��N"��p�o.r� t���Z���� �kR}��cok:-ckRC������f[�=P�I?�w�����>�-N,�]6�aÂy�ɾ|�G�
=J�P>��n��=?aޓ�=�������]��W����n8��S%n��4I3��{�T�J�V{��z$K"pG���Iъ!OJ�Hx�����1���nK���A.d���5sT��ٻs?Uܤ&ôr�����W?OT��@���[4{M;��m�ܤC,������ܱ� x"v]�����&���z��@�=7��x�#[�=�7��d����e�ԍ^��8�xuß(�c��3�<�6���l�vSE�> �o]c吤��{�]>��VЍ��5G���HvY�ɱL��X�(5oڬd=�l=P��!L����%X{!䂢��9�u��[���X�ʆ СvR��j�,a�,�J�m�� y�����燄��`},SKy�*,U~��@�'��-a+�OQ-J"�w	�E��_t2h�'�n�b	Sc7��N<e��ǔa��%�۩G_� �SX4���S���F| ���f�Rj6$$]�D{g]���ƒT�x<ksZ��jYi�d8����N�P8~ܜ4:5:Ȇ )�fU6@���Q�����9F�-��M{�voy�Ц}M)�r�N���}xi�d�S$�k<�p������C�s�9�ü)�����aG18�U�nA�39�Ho��ٷ9���<�����6z
�w_9� 8.�@�
B�)c/�O6���d�*xP�K�ɿ���7�@<����{k���o�v�?@AǍ�}�lУ�y�r���1����=�]V_'H��mU��0��@��:~��*G����b��ӈ�w����&�迌�m�,�WIf�8S;S?�G�+�0��׈1���[GSh{��q
c+�<��o�KE�y��)�ڨR=�lI��t{G1��O��㪝��iz��b$���`�52zo]��g���|�Iv���NO��d�K��	<D��d�k����R?�H���Ato_� ���T�]�k��c�T�{b�IH&ٴq�d_�j�DJSܗ+H����0�{_�Ga8�\TU�5٦�65���.I��1;���	�!U�z?QB��s�DJ"~�n]x�;��`�PW�*�Sz��iT��Rj��P5��[93�+��y����^��_��Yd�z�4"�B���ޤ"<�E?��'gfN�W6��%-�͖;3�Lн��0���s��f�O��{=͹�Q5A=KrR��k��9����d�y�Á�~�F��6�ʫ��&�}�� ��i��zc��(7x�S���_u�l�ډ�D��ϝ��:b��ݑΑ��\��D�^����ςb�Z8�]$���������j'���X��	��6��8���Rh�2N�a"�L/�væ�j�q�(�8���Ojoi�9b��K���1�!�N�ӹeZE\a�e�$�}�X��=��&�I�,h��ܴs8Ǘ������g�\�5Z�	0:*z���7�Y���Nj/�5s�&��{RC�#L��̔xzY������ޟF���E�u/����^lӤ�4l"K���6��~12�r.�f�>+�!^�����Ftp�����;��!��D٪��)?�^ԣk�5�^y�{�S���:���&��f��\���)Hz��p�������+�.n������!%ot�@�q��0��:O�x>R��~�Eަ6���œ�5�1��P�T���6��V�`a�X��o�"��,!�>����n�2a*C1"��A����1��Z~��+l�𓡽����Y��g�*�"HX3��ڨ�K5u��9M����s��
������j<;����|W	[��|4(�?My��YH��y��"o�t�-����Ʒ!=���z���.�D���1�9h��39=zFD��\���t��������
>QF�y�NKl�w	���cN����,08nf�q��c�.u�]Q�4�ƣ �D̫�%�zGW7*)��g��^IT]+����{���n	��$X�L-آ_�c��� ��L�k�_�򤄴��F�F�+䰿d�ߛ�PVQv,50�Q0<D�2@�3~5�n��P�5L֮Ҳ&�\~�t5	 ��~5-�ôd����؞�.9?������W��_���7���b���6y�8�p蜘c�_+\ăt�A�sA��C�9�<�ya�֙?6okr�"?��_���yO2o��S�}��z�iy���y,1��c+�0N����	���iG����kL��}ZI�I��uo֤a�?�߲�~��/��� �ş��>���Îӛ�-��$L�9�V'ț�ݼ����ʚ��6Q 3�d�q��m�ݠ�֮��uYX��OZ��kl@��ŏ�t�BF�J����A�3##��'�!�p2��L�a����e��]4y1*�a<�
���$��^�2�>/��N�Úv.�}EU�0X����L��>��jY�)�BNO�ZD��Ԧ�c��*�@7�\��u1`*�S$�H�|y�m�vg�+����:N�X��Rs"Bdۄw���44�3n��x�~v�h����*�z걍D�R�Pv�zf�}�ݦR�D�x���m��&�َ������f�kt�S爿��0x�GE �N�s�������Q��MZV q��si�ׯ�b��6`!���m��bu��uA�jԬ�W� ���*��|�(��tqd��!�@�a5��-2s��x��̏�3Z����
D_��M<��A�� �ׄѢ�����ܵ��iD�[E�8����`�,���ƪ�֙�R�(�ya�vl��l���L��.g�'�S��w���O�"2�iĩ��I�K��'����B�b�����n7^�yP� ��2�^�T�&<¨'�?*� =a�հ����t���{X��CM�.�
�V���gP�԰�5~^�v(���=^=H{J{���1Kqt���M�:����;�=�`Px�����A�fZ�+�v���0,�Sܥ��g�i�/���{�x)�-�غ�xȰՑ�4����Q���G�/�/���]hrN]U��+��ܟ�#{9�_{޵�"gf�H��,�v�ݛJdgv�J�"�Z�#V����پ����O�D�4���5	��q+���l�bZj}e~_���,�M����������5%�rB���7���ňXpW?~]�w�-��W*����m�����14L��k,�>���]���������[�u���2���AG&D�"I�Q���V��Db�ea�UOl �٣�}�e�J;�Sp����k�e���F�&#���TB/7&>)��_�-]CN�'��W�j�|�P%9�@#���-�YK}�;�	\��!,C�[NAb�����W�����We�$�@R�W���'#��J0G�O\�H ���@���\��DM�zA[pZ7�S)�gEO��/��:��#`���9p'�
�+�n�n�v�<����Q
�V�0�4	������2R��������'�_|�Z(���l�f� D���������K�-tܩ�r8��o<	#�~IU�KBt���f(r�ZX��I�)���A_�8�*�ƙ�9����jC04�V����o����w{|z��3O��Tz�x�B�R�k��e��L1le�dv��zbu��J��1Oz"�3���-3xzt �.����Z�R����Y�H��$��~��6aɄd#0�<��Z.K��(�N���⪕���P�fU0���	in�<f��L��xq���D/��v�3���1SX�V�j���D�q�V#���G��U�i+�l|���3br��'���H90ו�C2*�|�eO�7��
�]�2{�ut!��<�I��)�׫�аnu�E�K�ui��z�;�>n���I5�6�q���8��'⎥|�7[�:e��'ʸ�E"6"��?�Jr�ݿF��%�B�da���ı�̒���Y�z��8�>�u�Jbh��4N�tHU�1)���^fhʂ�]ˮ֘g�T��hj�&���@=T��
2*]�}�:&��_�6v��8;(��]x��\^����-�D�E��	�Ue.�ӊ����,�,g0hgȄ]��)(�=�Q�Ǘ�A1�Z%�i�ˍ_ͭ�OEV�4��)��U]c��L&t�O���q/��v��Ժb��=�{ȉtv")�,��C�W<�Hˆs�Lj1>y�~&�i/�K���jZ!ӉG���湢-����K�MQv�L���t��o��3'�A�w���z������$c�㱑H�/�C>?�Z���l�?U�!>�4-�_�S��*!�	@fV,p��p��0b-�����!�k"�@ 4�aE[u���W����9j�\���q����H.�1F�_g0f�A��x�����]{M��	Y6��/�`(�ǘ��j@��K<p�����@���en�+�9��\�s�e��~ŧ�f���x�9X�S�tt����(�P��ԧ���<�����E�	Sjk�D�i7����MA4'���U]A��?bR�NFT�����;���^:��>⊄c�^�����oy{h�����8�e�[M%��.X���<آv��no�<�3h��ߒG�biOV׫�=���"�k�~\��L��(!X�t4ˋ.5��Q\���Ì�W���tu����D|�"`��� !�?�������!6P �8i�`�0�]��jޯp�_Le��䧢4��b�����iն� G_�!��:�'c
+!������DTB5a�o�������r=���'O��B��Kix�򸔾��I �,�MŅ����������(��b�5���Zk��J<�x`��<�%jw�  ���sB�x��$���'�Tt�(���k�[��9e���!g�d���$�Ĕ`帅eOK���Z�A��1m<��r���pƴ�-��U�d �Kӽ�
 q�#±�9F$�P��筱7,U@��:ժd�Ӑ�ik�Gr�ݣ[��Z,-�.�}-���G�D|���+L�ш�MSV�d �X��:6(���ۄ[{��s�+�Kyk]3��A؏[�~J�+u�,��*�/$3�[1^d�}k �d�V������_��}�(�7]��W�܇�'�Ri�!�5�mt����cj��|�C<�Y��,��;�J8��$bo؏VԈ7l���mG�bx�+n��F��)b�/��S:��,��,�B�ι�rJ|����#�qP�k���'�YFw���&�	��Y�ﲊg�кë�o>�C���sr�Y��.?�Y�A�]�݀� \I�E��� S�O8͝�!-�=ť�ŕ7�H���ާ)v3x����)t�����|P>��Y���*80�ꀱ}]A��Z�g�ҏ��<&��?a�ׅ|-�ƫ�.JK��L"�U�u�풩^I�݌'{����t�L� ��wn�a
���&�a�L����׫V�U9���yA�C�9t��A7�#z �
�����&[����(�P�t��d�\Ц �8�Pz�e�~�v��D�^���R�Ĩޖ�	|<:7�R��P��F(#�` �� ^�gTQ<�)3�v�b�[c�^>�-�.gAo/��^W'0�a�r�73��Uc�>�r��x׎���Z��ĽiZ�c�w�-�a>?־��*����#m�m���C�8j8w�
���O�L*!�_��M�U�ǈ%3wa���q6M�dEH�M�I�(�	�͊d�({�j�\���6c�|��w>�6[S4:[-$�d�E���1@w��@�Ԋ���� �	6
 *�r��D:<��7�F�U��	�!^�-4�};L[�G���L �@�BB�8�~|SFy���{�7^��}��)1����\>O�� gA�N�8����j����<��](E�S-��j�Z��𻦿^�����wc�Q>��n<f�Jz��H���[A��Sgn����4��˚.YA�v���������ja �{	���6W�f3�X��f�<�50���DW��ޚ<bb�ᣣ�Z���"��7�<�g����뫰;>*��/6q؍P�a�����7n�Sn|�'�r�������IU*(X'�Ѕ=�S�!f�������T`�Ft�PHW�.m{!9�2���}$��ρ)�8}��P�pu�IS���'u̏�.a�4R3�2p��ؽ��-�Q�K����!=.�h&s��/���V��w��׸��\z�>F�6�+����fu{���%ؑ[2�c��s�p �P�r��S��M��}v�n�d_U��^?`X(d����O4�<̇T���$��V�b �H2bWtA'���^���v�dh��`����m�6xiWk���U$:�{�<�s�@�1�j���hN:�����A��z�?�hB��s��c�yyТ%�{ ~�ږӄ-xł�\���ܤ��z���-�/�S��XX��VnyU�'��q��~���Yg���Ng�Kg����=�κ�6��;!���̽�&�:Y��9�? �7}�^u�Y޿b��<�����0ˢ<q���S�7/rř�6~lI -�y��z`��<�*��#L��{Ѩ�w%���1��S��_2�O��*�H�K�����c��߾DȵjE9w�R����آ��q0����-��5��g��&�k��z������cN6�x���.1c�����N3�����Pc a��fï���]����'Z��y�\rZœ��ű��{�f3���l��ҴHk)�ib���m���Җ�k^S7j��	��C17O�[0�-E�C�rkW�S�	�)4�IBz���Z�����)%��	��Wݙ{(�_K�'�~ܛ���ªU?��{j\b�ߪ$�ޙ��q|p��L����H���O��w��Fa�B�j��P�E=�=I݅�h.��{�D��bW_}	%~˜B�:N&卍�����TsB�&��]J���YG#��q��EoMAB�_�T0!��}��@qt��"�ýM@�ݭlTC� ��ʺ&:��ͬݖf���x�ܗ��,dS�X�y%�7�Y�!ٶ����գJ�ݲ�u
������i,�_}��Nb�Iib�$o��������3W���p���=�����A�y�0r��|���x�f*�9Y�ڙO�M�u��B	�A�)��%R�ŀ�P	���+��m���*x�X�RO�����EJ;���� ݏPk�=\��O7@N�0=�\�ר�oY�Yq�`*���"� [���/1'�r߭[�ݳ�Qf�S",&NՁ�]���4�(+�Ț$��?����W1���0W�L�{=ZzI��\�;��n�rfT�:(