��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�G�'��"w�$���9X:pe�Q�e?��K��Gh���C�"?Xk�A�'�����*��oO	�3F6?����gK�U���)f��J޿�΃����y>E(��-?Ha�T�s��T���Q�.[Ѫ��;�����˳��5~ߛ�/��`	Ā�^��qsR�(�_49��%�(�{)�GM.�L��'�i��MQ6�v/�����HB��PS�2�d��������Q�,쀬,����]*��F)ē�:���C�s���0OWK�j(;%t�~�ӥ�U�Q���DҔ[w{���W�r� <�)	�H���L��1�:ڕ����g�/��uS��6���u��W~�o fa|��9�(��k���O�%M�ӂ#����[aT�ŵ�6��jr���O�}*��݄�n�Ƞ\�Ő6�X�.��4�[Fj�XF�A����.�����r5���0�(XZ�|O$Zޱl�M�Nm�qh�8�������Ѷl���j��iaqn�P��k���t�d�7��ϕ@@1�3�g1��<�r���%uǜ"�8>�Nv�D�u�Qq��Ԃej$�֞�X�ª*h�w�wϏ����mM�A��OA�>�@���{RsU��uJ�E��K=Pj2]xΏC��6�e�-*� V�c�PrT"̖.����j8�*�(�I	{����~�m���PO��XH�+=����~�l�	-�}�fay�<Һ�#B\������G�Z
ꀊJ��+`�2�X��/�|8^����һ��������a����K���	�h���w t&"HO�:����Λ8EzL(���R�܊o]0�MW��~<�/����oS3�Os//f��į����n� ��w��4��(x����[�NS ��]&Pj��vK4Y�9wD�@���5Ow��a�xN���|`��R �7Ք��0)|1��m;��G�H-^Хڵ��a�*M�?5J�%s����}��gW�bb�c�r��|
'N�r�A�tg���65+�-�(�������N�2�Π�$�r��p�K>JK���#k�Y���������EW�[��(A�M�����mrp���/R�`Ցˑ��`�0��Ꞛ̥&����<�`u���n%MHv��ܟ{�q��9[��͂�w`��Ȉ4?Gt�p#����3+59�������2`��!��l�0(o����N�q��sB�*��4gϹ�o(p��x`���;\��� �Hh�-k�f�gt�6[��t�z~����q)��,�l�fMF �L���,�ChloT���q<Fc���wd��y�P> :y]`Gm�3ۊ�U��x�ޟ?6q/U/얔^�$x6�*�\=�V�άY=�J�q�l��x;
A���zI���L�(�1ԙ�/KT�R=O���*����cV'�ͩycc;��8�#�=���t��`F�|�#�����WGx-�������*����ֶ߁��Y8E���L�(K>�d 8�@b�A�������X
��T"�!�����U�A:�����Bb�h�>w�ކ˃E�92��fs��� �U�1!��X�Q|�����O��
�|cw��,:0�Ւz|�?v�``c�w�n�,j>�aV�wq�!Z����ζ��T�]�JA*���m��ܸzq{D���uD���ռ�L{Ƞ��X�$֩�JM��Eû{���u��2���s��`��mp]	̆�!0�s���H�|����.�S1�����]��~E*+���N2�.��!�:K`��썑�<>������w��0Ý/����-*V�<@&����"C�c�hdණ�sN�-�S28�)�"; p���	��'(ȣkp
�Y=�I�8��J��`�tM�߂��<�� ��o�������Dgn�n������ ��V,����������LU��a��%o�a�5��^�,K�]�\�P*WB��h�<	e��Z��-w�[�+E��%��4�����KE�A�$���1�Lͻj�� '�
�/��Cq�������x]($ƨ�J���]�ʮ�,�e)����1u�_7e�Y�Zw!p��B��$E�(Z"O�aF�]`�\f��{�{x�%���F�Q���js,��t��{s&C��D.�u�#�����y���^�	�nw�oۊ8k1D�
Z�K�ԨF��=�	Ұ��(�vL6�����H�i����F'�^���E�ц�p>�7���T�p�L�ۧAe���Zw��:#�I�:����ʓ)1�.Dq�e�^�)0j�D�mh.�6z���}�:�Ό�qe�/��$�bI#�#���+�	��ҚѮ��\Ⱥ�m,xEr�#�/v�`�O�6Q����im�H7��$Y^)��|V��{)��������s"� /+$�L*@"�a�p�W�#~�P&�.\�Ͽ���C�2��8�fʺ᤭.�Si� 2�U��M���=��"��$j,��OS�|�1�K1�i h��l����������qɟ/Ų�(^Q���m�R�"���ְ��"�0�'μ��QQf�*����c���ׅ��X���I��J4\��͘����q\�NH�"�Rw~ߛ��e�@���ù�+(�����e�Cj���m���W\xZO9d�O�U�Y?��8�]'n��}�����@J��8k�9A�Z
¾~����畳���Ƌ\�}�à��h�
=�*xq���Z�p�Z�Lo?D�z�x�=>}f"�3��������l�� ��+�'K@���_:�����%�Ϫ�S��y���u���f�`�Fx~cn��zsY���&���kq �X������+c��8��H�^LY�k�O�P\���־f�#!�M����1J~� �����@��#�68�P���X]��LW��d!�̺~�h�����GH�p�z
e�*��b�����*����ȣƳN�b�S�����u��3?��WM5��`���ϙ�"�;��[	Auh�ˡVn��}�)!�:�ݯ����=�7�7��˃���%������\��}Iy��O���'x��f�w��0ÍE����6_ج���}���Z��]�;�q�[�q<A�UW\@��w�K_}�[�
�G?Z���@�ޞ��̵��@q1���?�%��V&�X�����M���;FX�q桮��zG�k]hFU����8|ٍj��i{[��Y8�_;v|�X=���;��E�#�:r8�2-f~�,
���eP*ۇ����׉04[�Ȩ���c;�|����_��ٹ�;w�9E��ƫ�#4UICe��vi��:��ʔ�^�<ҭ�%Y(����i1|���Z)�߫K���\�7;���	m�)ISc-�@��4m��!/-h..ՕV��޺7�o�8��%������Տ��\L���XmWbC��-I��}㙷"�x+��� �;)�"��	"��k�[��r��o��#���*x{di��ĳ��7*��˩���k�4�k��a
G��]}+��-T���t~[�C���� ��%�TY�Z&�Q�-Q�!Κ�=pC����^��4�ke0�X#5�E�H�r�ba�����{�`ԇ h� ��[l��t3�a�+d@a��]�|?�1G��W U3c��i�t����L9��A��/>�[�k^,�9�'ϵ+xq���I7{��e�ZV�ZA��j�+_�'z���R�4���kxN6p�#IHL��*��HL��~2�̬��%��ɀ+��7VG�Y���[uQa��T�ۣuИD�k�tLD�*������g��}wɼ�a�@����)�֖�iq��'�!Q);�B�o�d*p�#nϱ�����f��{���o��b`F�b)}Y�%^4�`����k��PltN� ;lO\��p1���]љ��uۅ��o��`��>�Y�R.⩋��2�y�|!�$�W�m���d��ɄQ$^����im��A%н+�G�P���?����z䶃�@�e��Rw�"�n
�֯�%� /YJ��Ye2��ݛ�XhgNI�m�t�d
x��pi~5�H8�BeK����Z��H���]�ߩW��KSROX1�ok� M�c6E�\��&��l�އe�>f]�@�T�u�tgG_+�.0e_�X����0<��\{5���z��L�-�
��i&���$�,hw2E�Y�g�R�e|�㭪�D:?A08���曎j@���Kxb7�5U���Q�i� yt|�74�X�a�_Z=��\� ���Ƕ(w{>D#p��j�K��P3s"/3>zʓ�s`�L2$8Oӷ��~�껟�]��o�n)&!Nڭ��Ԥ���m_����~�bm�Ew���b�޷o������<#�\GT��SI֦�-�-6���������ʩ�L�4�sD����8"H�|�S���2I��wr�x��<�yK�2�J��_�c�uz�ךH�@���^�����tO�1���Эny=���`�o�m���~jR[s#w�䖁\��t��5-+��%�4�?���Au��)�	�J��,"/Z1���+KC���J���%-��9���,���}N�>s��'����h����x�
��J/$ɐ�NrNK9J0�Wc�z�6\�L�W�еFU&-�(�"�gUI��V���G�V-u"ٛ7�0�p��"v7�[����"����ET�cg/��עxx7�E�-��B� ��Ҭ'�/�����[��o]��: 8L6=	bGp��Q�տKn"���*m�Sz��
}?p�Q�?VJ��dYȬ���ՋYg�R�UT$��Ө>��$�%Æ}�3]�MB�*�cb��������cMk��:�z~�X�I3�%�Zdپ�O�=c��g<oC���K�_��ua�ٹ�ƒͿ�J��"�����{#��P�+�l,D�����%R�9�JD+�UlB|���������9�����9���1�I��)���&�[�V�{��[�*.�������(���e���(���l��`�H#:1> �-�p�)��Hl��a��Ҩ���r ՃCzU֓#��rm��R�V��]v;���>�F.Y!�)8:�CrM5���Pk֤oI�,2!X�*5s��)��"��bw����Z�@?�sQ�#�a��o	�ͷ�^�9��sI�@�2���7�i�k G��% y�:~qP���������,i�dR��a����n|�OQ�c��}֌ֹSC�*f�i���!���1+�P��M���Rpp��Z��`X�	��41G��&�5<T����d�i�}f�?�"�@�$��.Q������[�5�W�]p �·۔����^�:�@=��g��#�o�?>�:R��&�|(��Y�6��yң�v�G��bR}���-����nIA],]��k�3⤂.�6�y,�+���_��O���*����P�Rȑ���`rn�ɚ��aq� ��f�춦���I��:��M��kL����3竻k�癗���e�S�$�ߏX	o���S^�4�Q��&�z�6ϦY+���)^W��A���at|Kj�鰴�3��J+���t�`{$������/#ω��^��uR�瑞X �%��:�q&�R�U(rٍ�FHӛ,�9Z���[ @좗S��Ͻ�MbH�Ӕ�� ~+ؿF��P}�s�.�MH�Wҩn���\Q�x�]�N���}������q�>�(twR@�2�S�R��7��řf;��_D,_���D�B�SD{��Z��8���:*�ѨAz"=��IJ�N~P/�rl�kEc���L�T�X |/'n��Q���MLaϱ�0=�7ƵO\
�����7#j:�X���hP-g�uv|�F����ů�5�8>�ꁵ>���D����I����I���f-�T~C�2�;��nT�\��!I��1��vM%��Ea����K�è���W�v4U�Sa��0F���U×h?��������ڃ�>��DU�_4�-<ℕ#��½���h��h��d��9��uBj�fB?��t���6��@d�t��ָ�r�0�IU]���Wa�Zh��Sm�DW\���m��>����9�S풇��2�:�������I�}o�w(�@j�0]���B�ca��P:`��MB�HD�\ױ�#=z�)l�i	��U lyv�ط�K{�a���R��|V��'��D�&����o���$7��M��-O���k��t��������,����5X�@��4������#͵����D|=�oI�5q]l�j��u:��!������t�Q����_����F� 4�1I�ɚ&(�˂�\��U³|Z�<w���L�E��I�B���ٶZ%�R�w������*��WO/���l?�20��iU墳��wҰ3���7h�g���������N_�tƉ')x�|� >��4u "�Ό�����c %�Gt f�@��i�nl�&�����F��srFkQA�^ݢY�C��p����R-����If<�b�ۜ�%�-����ۚ���8ef�����x���	
�M���g1���
����.nz���j�Bv���gz�_�&�/
�" ܴ/v;��Is������l�Ŕ� �Q{�S�c��<N�PPND��U��멆��o��.7,'�.EU�KW�v֢�'�dq.��$���H��2�^@��wk苒�����ƂG��+��!�t?��/��'��9Q�朧D��ű�-�9��~��S~�&��zYĖek?�*�T�j0��'�Z��[��S���G�d�A2�p�8)XW�6���c���R
t�ZpC��l���_9�i��4$؆��|���#|?�L`�C�p���}����o�8s�];���Md����p/�)F�?O^H��>�?�t�fIu����#ִBͨ�)7�[/�yh��ޣQ�5<C��q����a�q�o�O��n�3coHֈK@Y���vi|�	�S��n��è�� 9�r�l�!�7���k��~�,!k/��^����g&���jp��&��/�[��0gϱ2� �ݎ[�R�|�/�^h|����MSʼ$��M;�M��Z�eQ#F��gmD����M*>W�u��oPHED�����ýEf��c �[kV�(�B>֚��F����o_�(G�ԫ��4�v��k_�et6`���ŗ��5p,z|K~4�;�g0�k]ww�����x>s�R�2Υ��>��m�]�2B��o�W}�^�T5�J�.��,Sj��e�\׏�@u_u_����뉱\rH`��T�p]S���Yb~��Z�UH�=~iL,Ц~:�O$��J?+��v�qr���C���E�&g��[ۄ�uoªҮ8��q��d��Wc���� �
����T�Z1͘O���u:H1y��B^  ��s��XG�pŭ��6hƒ����hH�9H�%��oV�%���dOS�M��o����in�Ӣ�/�vR�>��.*T!�7��N����7#	��e�܄w��K�H���H�ܴ=XB 5!��7�_!/���s��CHDC����!9,�~�S:��~͂=�N\qƄ?�m�R��`���.ЦJ�;����8k�4���$)m��u��p
���)�O\�M m�NX�b!����.�@��t��V�����S����V�
���G�\~[�./Ϫ�5�d��_�?\	H�4�%�*?E lHo"�A�f���8𶻔��ѽ~�&�5��{��DHM߅-_�\�N���H�H��Yk�)�9�|�~2���ŕ�NAj�d���a�$���Au7����<�/�ۢ���".F��l^��J��m! 	���z�̨��2$8y��N��z=}/I������*j�<�{�*n*�&�m�+86�]�΀d��	�p�y��h�J�<����?D#�}G0K���k�x��T�>%�\��oQ%��J��
��>�zY�)*ނ5,C�ڢ��6g9����B��ϔf����c!�0�(m�k'�=���K�P�ǁ�`M��'h�p���_&��M��C�o�u_�"�h�� Y��<-�4е���*g쁪�(m��Mv������ɓ�4>
#{��`�`n\;l����XNg4NB1�@�G��m!�")�=٥��vs�J��y��C��*%r�g�Ӧ�I��/d#��h��C�'�c��LV.Tt����j��21FYG+�z�>�m��E��-�y�Z::�\�ث0;�Xb
�Ag��]�y݅|l�z��jAE@�,|Hz��l�/e `7���J�����"i�i~v��tE3@bi�!V �
�����T��j�ư�_|T���r7},%�D�����^p|T��Y.�M#m� ]h�*>�]`V�>���;���H��P_�2z�]��\�2��HN���Ԁ&�\�������\ξ�tlAҸ���H���Tq��Q�r�hTu�J�+�cwgӎX_L&�7/��\b,����qWق��r�3�Rs��Ѻ�\��������tO3��Z`���1��s(G�:��ǉ�zC�Dw����ҵ�|���d�O$+^������G�ѵa%�o㺕g9��l5)����k��jȖ�.�4H�?�k�Jp�/o���iﳂ��4�*p�Gj���w� �TGt�Y���f���-����AT�����o�i)�
��^��@�F�H:)?�s�|�%�lO������˺��ʃf�C�[_qQRٍ���|� �HQ��a�6�����㔶˘�ҫ�mQ�}��S�Й��K�,�oz���_�}�8ID�Q�x��rz<�Q�W�H�{��<�0�Q��?����w���c�V�m�#�B1��FʜrHV	�`��+{t�n���έ)FؘVD�d�g�d/J�r47�"���MI+�
Ɉ!P�T�Xb�7�:�u�1H�tƻ*D�� ��!����Z��q%SH~�v��#TbE��.����Z>v���4�7R@MR�
������s��^��ۖ��.�d�Z
XE��6"N)���ʬ�������V���r	j��16m�ە%(��G�O0/9�7��XY)����9�oץ��^��_;���9��2�����:�<�o68j�(�[Dy^�^{�dd��c�����Pf}#��7�2�g�w��3b�+��U 5�3,ҫC)�K�BX���{���1K�x�q W6��K����B�8�rԚ�~���%p_���]E� ��M��U���%b�����T�u7)q.�^�S��5\��Pۛ�嵦v�h�Ïh�/� ��#�Gg��j��$:�k�4"	4�7�r��g��3��TsF���{����[k��GѺs����8�G[�saY�5-z��Sd�a�<��RJB?}�d���#�|_î��_zz����j>|t޽���T���G�؅�W�3|�T����e����8�Ÿ|^G}�+��F��JZ�����3�c����D�̔ф]���+�K�?��S؉=nK<V�p`�j�f�P�l��M(D�&�/8]_��.g
���34���$d��7��j�4O��e��Nݘ0.�1,�T(k�8�1Hz�,�Z��M��([ �b�E�\O��閌��:��d���� ���jL�uԉ�&�*��阛�P�q�a��i1�3V�SJj��\e��ヅ{�� �S���q����Ӆ�w��=��d��H�*���f��D�b�� �A�� �#LO���2F�]�ո)�h�{�y`��F�w�`bND��vZ^�{Yf��K[h����?�5�#c�+f-LQ�z�l=e�&��꧌�+X͝��m�E��*�\+�h]>�Bq&��]ա+�ا�d�'*�c�8Ҥ�䗶'�E*�ZGR�#�@�)���
0p�6�l��3���ʝo��w���O���zϙ�]�8e��՚�;�Ԃ�Գ"��Ț��V��|���6q �\*�Rx;	��~�a�X߸PA���e"x���v. s�~���������:���BR�u"��Ge�
D6n�c�]��X��w�5�B#����|��`����jR���+��: ��f��
-����^h{�ž��������W)�Z�u(5���V�N.�MY����}�q�g��Ya=���p
%t�H>��g�����}��7v[���ϰ��t\�[��6�/n��'ށ�&:c��j�~^5W�p��&�<�Hi*�(t���/�Ɛ�9U<���w����-�=��O,�p�h���1��Ƶ�]NT������ܗ��_��U0K�|_���T��ԅ��y�남Q�w0;l`�޲6��Bd����Z'.E�9����l�=q�Q��8��0bJr��M(&�o�΍�͛�c8��ǻ����k�ǫ!C��4��z�pҞ��`�R����pEF���fu���V_k�������A��6�-�W�m���v��z��1KG����|�C��֩���M�<<j������$�:s_���HL�B-N#5v����[:˩&�.�M��1�\^v{r�$����k����+>�	�O��$��k �hg��j�P}��,�(yF ٷu��A���fT���z5����FdB=*?U߱�����3)�NE�B����U���l8Z�Hj��� ��o�7*Yw�ɨ=H��Y���MjdR��|S�3tW�p��JP�`$ˏt��� (N��d���ڴ�F�+�ѽ��������͊`�<���B�g�ʒ�6�&�Jq�?|�.J���v$��r|��*��/_��9�{j&�p`1,������8�7���4L�SDh+��+��/�3K�/[���*W�=bQ��Ζ�h�pm�t��-.�-�<Uq9�O�
�c$�\<�j�K����=!���x�2�R��BQ"�t+FoK܎��e��6O��C�:�6w	5�-�;��U�<���:�@�����:����ܓ�N�!di-�t�ejR%"��UVX�����n�Y�������esS�&���ڑ�������r����ޤ!��	ptA;�e舚r j�����My�T��1?�ﭕi�����~C��d��v�T��*�ތ�z���ɶ�j��Z��c�yk��U�O��hʰ��I��O��Y��(Ip6.���X�o��r�Zs��L�,46��Wңx�uK,~[#e�b�k�������&��,��#���9|������GĤ� ,��"��g<˔�+�Aב�TEq=G2Hcu<fб'��"6!�=�L��b��4����X�ʘ�=Hƻ�ӱ TVd{�����	����ş	�r�WņA�ڣA�	q⃝cH:!��ZD�z����Ko_)�����I���.�mD]�+<�dU-�8�zJ���5�F��^g�w=�=�*f��O�<�[4ǀgw?��y@��|�?�˜f��)�oC0���]�rr�cځ?n�\�7�<r+�@��~�P_�$�o:l�����_��X���N�$MA�P��O�pi��X���4��Pu��x�O�y�lNϯ��$��_N�"r��KfJ�[X�g�K�"=�G� ��T�=��r�r^�4���񼍱'!k�wu����쥫�b���0Qdˇq�O�'ٿ܉�b��?��)豟�,�S�_�� lwv�!%���?h��ъCXr�<kz ���ԁR�K�`gՖ�*(�8l)6� V���Pc?�P����c|�q?���Ϥ,���XϒFn�[+���)qb��{��Ra�ѡ�(���y��*! �\-m��J"�.ň�_F���!k���Ƅ�1�ry�^4.[�g�o��_���ϰ��N����7*�o�V���t����lJ���;&��fok��%�9�d��o>�˥чڈ����-�i:�1;H�.�{�� x�ՀR�Y�g���� L9�k�lz�����'��rj) �"�����T���GU��خ���,���eB놎�tj$-/�����jS]~6x���Ҙ��twu?�-焇��_R�i���ȯ���>'�g�xmjX1i\WY�;�u�g���M���^��MQ�<�-��q���1���o�lSp�r[y�?�{=��Q/k/��m��ε���G=V7�9�җ>��⺛J�>0�GT�[���#���lV�1�p_��Ģ�we��7@����~ؕ�!ߔ1����2��X�ڳ�̆r ��������e7��W&4b�x�k��vR���̡��Ca~x�,˽'t?g��7ϣ��t^�{/=(�G���n�vbOrH���7Y��������Q��w� ��G譗��j�3���J�`�����e��$2����V�0�X���x��?ZU�%2ͣ+�b����"!#h%����	�%ꋰz*�Ս�.������d����mPx'u�@���Ep�YsTC���:dm7�*5`�v�]�k�0	k`NX���OD2V�|�۱�pǛ��xH=s %���f�-�ף�ra�B		�~�U �SFS/:�����e��l��P ��`@�e;!DiI��ZT����ze�H<���d�#Ԙ>�Whۗr�t0
>�'Z��Dtӏ+�Q�J}�k�#�)��P��h���W�7�́�-S��b:s:+)�Y�۷���v"�&�5zA
)%�l8�bm/L�>B*��M��\1�GZH�]l�]@�;����>@�
W7Eլ�����d`��VB�l�G7!�Z�
�pb�-�3`�࿿J��ot@?oL1��S�:N66��jg��̑�Ó��[�5!�I���