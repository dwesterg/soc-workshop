��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��P6��%s��Ʌ�6�x� ȡ@4�L�;E�*����f�įs��mg'�iV���0�j,R����j&ت��׋�a�y�6% ~،ii`��-��t���*�R��`������U�q�ɭ��#�O����>�V.*N�2��pT��Q?8�'�%#�D,�����*���m��1�WU�����Ȼ�/�S��Z0����V���rnN,K�=g���u��Զm/x{�]1r�9:w��Ky@�2��E9�	� �X��M��6jMC�?K ��7����,#�9x�M>&8���V���y������T��|e2�B׈hf�lH�ٖ
�`����8��
i}M7��n�$ZČ0]�ݓ�d�E$���腡�_g������%��-��*)բ�̚�sP��S��Ae������7��M���8�����ǜ?�J�F,���&��~� T����GORf���_r�L`O���闌5��r.����I�����0^
y!�Y����!�˦\��M��h6u_����8�M�4����.��+�o�گ�w9~����x��yk�ck�B���>���OB'/��jN�h]L��7�uqm��F��_���F	�t ��N��j?֎i�&�й�B��GY������ d�x*���%���R�+V�"�֊�/!�Fi0�H����k�X��+���Y�2{X!��ե�"�Ȭ B͗�3F_&�@�����]'P��������V��g�I���^OoP��M|%m)e���x��51�vBC���GmFA
��B��b-J� ��NL�l�0�<��:�6�V�<'m�1�����p䰷"� Y�7�.��f�K#*Y�v
���,(�8�z�0:���k�-�"jw�DC�2T�*/�Q�9� �M�5ۚ-���Y�����S�3_��ڳM�EZ͛s�j��SL�d�ވs�-(N���^�	��oυIR�E����MsB�����9��Gր2��c,�=6A��O���Iռo��?^�N}�S�����>U$s��,rWX��w�2n���yr����'�X�@�ڼ�D�_�A6�E�v�5ӣy>�Ѯ�L������'#8���O���鈰P7>w��Q�Ь1���(��7����<�3�5��������X��;����J�β�d�'�Vﯷ��Co�h�$�4����v�Z��m��U�]�ȁ��X҃�7���Vy�Hd;��)
{��-�4���k�2�ޜ^���Ϲ!�Kp��l&Y��]KNf�����]���4�)6�Y���a�,#޼�v�uwr"��s��� p3lO�f-�%n�W��Y�0'������N��T�!����aO�2��wɑ+yn���C�Jhfi�>7�J#�g6�I�D����I#�)l�+Ѐh8���U%/��/ϊ�֧'m[����t�#�)MYֻD� �Y��ح2��"%�B041љ�i6B���u£%�,�8��~W��f{�^��י~D��eo�6�k�R�`�~������$&�v�4��Z}@3.�$>���7��