��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�TOg�S�(�U�3#���ɉu�{+�k��
�w[2G�W<.hS�b��A�X��$H�7.���D79��-o0�W��)�6��O�us�A��\\�D���ҙ��v�:�P�q̍;-��4�M_�/,Ь��h
�l���!�V����(�bS[]".�RUM�.�7�m�6-V�T�H �lRώ>~���/#�Wm��������� ����Bq��2t�J�Y��i�����H��NU�lL#>������F��m�2��ex}ͧB�#[Q��������q� �g,R�b����@�1��S�����Ȩ'&�y��L��֎ ��gP=�m.S� m���P>/ڄ��I.��.���Z�I��͋-��#8c2��ݫ��\�ӡ��2b�,�������u���2�a1F��ܣx��M@9��W� F�
���ifF�G���w�_f)0x��+����f���I�U��~�d�
I������%�������*��MN��T8v��cW+��7��9�;�G�i��翳��	jEgE��p���6L;�����.�����HD�C�o��a$��k{�F���J ���<l���52E�	�u$�>��Pi�?��w��^�a��
0~���!����iα/ץy9������5&ܢ��j(^~�>��l����v���
O	��?����z��`�>��4ޭz�5�;v�=#��4&D""<Y|�P1E�|�ֲ����,����h$	���}�ႀ�ᦔ�
 %�]Bon�BPh�ʻ�V�E��R��f4Z)�f
��7���cui���a2�l
V�^ڰ��4�(�����@��O5�McF<(�`��"��w�0%�3�?���æR��Ůd+�6iM��",�388�,pp�3��~_Nç�� ���P��|�M���5pƱ5�)��e��'2����|�<�`��f�k0뗓O�e��%�,�;�-�ߓCNS�W�Q��Y;�+���)S���3���5g!�Vp�&������^�/+�͈;D�0� ��4������~e��d��g>��pv�Z�~����16�V,�ٽ���֔Ŵ�]��vY�3�̌��b�kT������p��bi����ԟ���2����ۤ&"�ng����J@�2�ݒ���L�.��v+z���5��{Õ�����W�ׄ0�gpD�B���bȟ��) �� �o�g)��m��0�����b �틣�v�R&����Y�=��ڃp�^���64X��`v>"Ɖ���;�����>��Tq8�^.��8������5&:�0A� ���l�ܠ���U�̍v<I����������A���A�wKG]�W%؜m�ޜ.����t�|��	�#���i��@s <�h�X����T������$�M D@D��f�ˀ���t~s/".&��� w[1}8�y6?���^��yn=u%�3�<t���\�x�'iHā�����)�����&ybi��G���*(s��n2PM1+��Z��O�*=�\�m�.�-'�l���:o�z5 5q��|�IJ^�՟1�c"���r��i3�O�d!�3/r��yn%LR���Ԋ���2P�M~#ȪMbs��3Č���IV~��c�ܥ�-{�S��]89j���aԫ�<�=7��{�+1����g|��5���4��^zR�X�S>M�6����l*ق�����	>9suE����{��@�w�t*��*��	���/�|b��� ɰ�()(�:MWփ�o�Cqa�G�ź�����f�78]�"T_t��L�J����M���Z���m`p��N�
{�	,D�<T���_���x��E2�l.6Ĥr���he��� ��f���x{h���s�Y���DX��F�z�Է�n.`?<J�Ef)H��d�im��ݷ�����h�%$���=}53�X�2�|�wM��qh��&D������83�qR|�M�HF�r�eI�jv����碤�#J����ϾR��j627�E��~�C2"���"�κ�A@��@�ya����Zx�<X\��Q9|-��9��j�w����e���R�í��S��
<DOT������:Dѝ��y%/I%�	x���崙ӵ��%�Si�1k�}�Z3Ζ�23�Л����]h��^:��n�7�/Ɲ76�EGh�+z���S=�2�r#|Y=X3T���N�uu0-�������,��<Z��O��&����"`{��A�-R��a��{�H!���%�B|k��!ۼ����W���Z�WR��U!���MT7�ĘHZx�����ن�b1�{TEn ���`#�=���t�<#�]~�]��p�t�Qa>h^� )S�..����|��K�k�BMK��x�mb�I��l�5�T�v���XXQ�����B��)h�Pp���`�3m���(K�@�8d��츴f�kM�a ������;T�F�
�N����ԩqZ��S�]]�>���'��rK��"D ��hP�ks�ֶO�<Jl�d��>�V�J{}z�B��t��ҙ���cݤ��Q��d����2��+^֧@M=+���G�jƺ�ҵ�������G��Ӵ�$���-�c�BI<���[�hlg&���y���dʸs���#� �;mWx��L���\~��>�u�K�^y���Т�_�K��He4�c�E����60zE�`����.R�,�\ֈ�=H��H��,����뚅I��D"�k3j�ˣ鴹e�֌Uy~��T��)T�j��æ��,Sq�].xT���3e]N�`�$9�ۿ'�X):�0|@��WF]U�Q;@8�x{
�a��x��-��;˙L���D��a��G����{q�F��f�W��z��F�>(���>�t�v�9]�چ~�r�K\��U��0L�Aҟ��I�M*0��]��ly�7��W����g������'�=j�E���!� �l���`�x��U�_��;��B��F�C3��+<@��4�ډ�@�`�B�k�������4�Z��ۙ%�@�s�*��!�b0Y�X�f��W*���f��5�kq ����d���[�U`Jk�ɛ��-5�%@��t-3�5��_�C xN��?C�z�s��P�pz{��I�y?�{���5tP�� F���
��xT�\7g�U��cޘ�{W�h���t�i<GV��\���e>��j^�_�	T����Dl����wxlFo${��r^&�����B��e'>t��EĄi���7��R�DK��K*K
��1 �!)����-2;�*�����*_,�:fx��a�f>�����A��� ��i.+���^)&"Z��ErZ�1��ٟRmXv��O��v��a8M/��g��H.��	��}>٢�%�?�LwyMx+�<��?�X�*Z�m�8�zBE$�ĝͮ삕�ykH��d:�d4����y�K���v�#/>�^=]��=����f��L8 >A�b���C �9�5�&{Í�&;8,� �n��+�6�Hg@t�P��gǀ�"�C�
뢂��l�3��h
�}�����:�O ������RA�7Ś��4�d\� ~P;�X��8��5	Ζ��ڷ��g�J$�S�/7�+��1�#&��VR�aF���XH#�ķ{.;�����YoF��L��C���J���2��	�s���է��KuW����͉Ӣ޳v�܎�X��49�����~rI�zZѯX���}��Iۂq
����3˛.�,�~�֋�����Y�WLb[%�`� ��k'����b�0z���c	O�6B�J#/x�')��'$d�U˘u(C�3^�6_�j��+,�:&M��|j��Rt(�)�|%��c������uX�0'�GF���F� ���~6�����MY��u���)����<5�y
��&:�K�3Id$���oӿ�je��;O��ւ������NE=i�7��x0��UJ~��V ��m�\3\���m����x�#�C�n�hA8���U6��&��H ��7Z �F�}�j��م�(����R䷼f��t�0A��Г �l�sII�dň
j3�3��j>7�{��4�8�U/� ]םGj��U�@�SFEdN�L]�ķ��X?�>��Z(.�%���m-���	�}��d�Gd�	�d���Hh�J�TvQ�*-f9��P�H��:�o@>��3#�o��7N��@����<�ݞ�I�W�<*0��H�y�;p�*�*�s�s��0������ڜ\5�҂Ig�_���g� ��:��E0��U�\-�F�υ��1A��I"	;���ܳ߻#�z?4�7z���ގ�%�:�DZC�xGh���50��>q�ډ�3lF
�������-]����X3�\�HQ� 0�.:���q-]k�3���Ur�޴c���vl[kHPٯ	�F�"|O)�3�DYkY@�2�k�x�-z�#F5ֹ@h��cy��b%朷�Tj�|�2#H�ri����5��n�'�z�5�S�F��@��)��/_b���[}m��td,�Z�D;��M҅I�����D}��Bz�Ns�u�{��qڅƏ ojp�ϗ������V׃�h�	�=�Sxu���ADm�jI��$�����rTCR�Ɲ�߉0z�J���xH����X�a���xR�:i�gV�,=��U�g}3���P=���҉b�w�5��Wc��.y�r%���)?Ł�%�j�[!!�v�$c�*�E�������0��Dm'"�)��5m�'7����dѷ�p�J*	؞9���͠�5-��D^�)�����|�v��˱��g����8i_���)a�Bp�;O�0&�`�w������~��5�|3�<g'e�N�
Z�B	&�.�țY�Ç����2�x��B}���#���g��Ƨ��>x�d��T����X$B��I�9��MLY���ۢo���L�Ui U�a)�D�ie�1Í$�P?���ВߺyK^jC�S%�7O�8�� k���Z3;G���1jy��Pd�1"B'}�|�}OW�Q�"4-��Ǭd�_����`�(}�� C���q(��F�#\{͍��[�K��(��y H;�d�'��f��Ww������,�= ������gUQ��蒒��!$Ar���}�`�y�������y��aQ��z�|�h��9" �Ec ~��r'y9�7�K����)����8��H�&���hT5BFK��V�F�N����Ԩq1m�T��T�7��K�����=�DܤUz#]f�fC�m?�x����1���	�@O��i�W�NC�Qd9�2d����-6r����jj�C=&���������N�HKҰ��N�O'������sB�l#��ٸ^'�����d���sf����/�2S7��L}!���HLYmxǍ ����u H!�� ��o�����:=���ǁۍH���ؗ���b�Z?��Լv�@�!����#�����\��@(���CL �tgl�=b5f�e,&����(�Z������Z+��W���
H�'w*�:�S�x�;JY��_���c$: \\���=q|��%��� ���x�ЧY���ӷ��-�
��q'�F����ȧ�W RlP��&u�?`4.'j���r���fF��6�{�ն�_̞�#,N�z�60�2G�L��~���5K�"iW���$qh�����5��z=ۦczk6����O�_lyyI�6���S����%��;-\�f�I_4�Dْtm��W�������9��u�K�:�z��V�m[ g� ڙ~�����\d=�_�*ޠ_s2��̒�E�"T�3g��l�_��h/�nJ*D:�����-P�;5~�a������}Q㓓�G�pK;4wޏ�a�bX�����-�}6�w��Ƌ�AN��@Qc��V���*�^���F�N6P�	��f������k�/�vC7w�ތ�JC��_P����XXJ�e�e� z�tB�]���;��7���M���pv��'�$V{!���}K5���v=j<״fd+=K���'ѥ�|�\���	+Q��"Z�?��3"zN(���8i
�X"^�ڡZ�����^��;&���`������ˈQ�#����]�)�:(�)B�.U�>��,8e�o��;b�ܢ<N�!9b�sP�6�	�qlJ����	���'�¼-�p�P:��F{a�g��X�sz�Z��6B��U�"^�жP�|D)�?Vǳ�* �������1�������*��'�B"`#7J�|]���+薫��I���,r�U[.o?�my�'�>C+�.o�D��WȏP�2K�ۍ��DQ���9�ػ��G�v�;��J�6�΃H�h�Cm���|'ũA3X��4m�%�Y���xޫ_��y��̃�� ���f�ַ��5Y���1�b}p��t��Rq�i��SW�=3�˕�]� �t��Q�gY�D(�ܗ��*���JiTx+H��\�����8��y4FvX��&&J�l8Q��Õ�$�GI�����ʣ�ٮӰޓ���y��Y]��ޢ���g���6�V��`���!��T�{ԕ?��8߈5��C�V@+#y�{{K���ʿ�P&�\�W���H����l��B�L��F�y(r�
�k%�p�+boQ°��)5�ף�\o?.�9v�A!)�z���.�z�9����z��xX�+����xՆt��1 �m�O>��#ryԩ#i�前?fiO~�ET_���)��X^���-w�s���'hy��'ͨ��$s��Ө���0DyǆIJ)�%�p _0�ť\|��;B|��p�Eާ �����r0�J�#>r�E!��p��'5fA93���Aذ:�DqvE�q�Eu4�b��"
aY�k�=��M?�����:�o���3@$<�y <��)����=�h?�1ggG�&'�%b�kl�.����j��бmsMC�Gn>d��r�8>$��'��ba+�E�%lY������\3���P���Pf)b9�&n��}�P���v����օ��� �c����G�l�g���v�c�PfC���bE��G�*��F�ZI�H��pU����
<���'i�,!_�w `��C�9/��w�Z���w��GP����.��[�t"���gCjG#�E��;�1�3�̍���xG��ӗ��8�o�g.@��oϿ��X^�}���\"*��6d�_� �U����~"�y���Ō<�~L'c�Ȑ�)�>|�c��u��,!��C�jb:k���Ы�W��/UNr�Q]�
�G뛔��)I9�}�F*7�mA�E��2!�p����7N�J{D�)S�y���L��:s�����ٲ<�δ'=O�؟Zr�'S�%. ֐$���gؕN�n����H5T����5z\߹x�E@�*�;���-�XC�"�4��j�B17��'��8!�5�+��RX#�a��
#��"tUi�r���6���)�iS��ډ5�ɘ"���T�I'�vH'�޴3J<I�{9K-�UfZI{l<[�Zj��#6�.I������-��ZѾ�6���6�Yy[
���Ҷ��d�'cC�i��7��:N��^�ܻ�l�'.��$��	L
;��*�M��ϧH:!�H+�����' ��8ڡ�f��
��um#��W��N��>B�z>u�Å��aN�h2��"�Fȫ�ⴕvSk%-�5Q��nэ`����ɽ_W4k�ʋ}"GU7��8�Jv�t��SF��!�`�N�k���͠��K�~�;˧J�l+�
���7�q�&laΖ�@cǔ,@`�T���;u�SJ��d�2p�\�}B� ?'Λ�T=`ف��gl���o�$ �7���ܕ8k�~��R��K��;�j%
���rp��O,eo���(���n�!i��3G�@7�)� �j�8��,EL�Q�ҍ���0�&�s���o��;S�t�||��k�v���?��	�9s ��2^���wEnhh�r�a�0�0<�A:���fD�Oh���^z�ٙV���g#"���8v(�p1,t�G�oX��w�@��/�w߫��z��������j&U/kZ����2+�la��V�m�2�=lsSS[Pf�W�^�� p�,r's]�o�GL[��jy�QFo�x7f��w��j}�|��	�fm�2O�l_c�r9)��@�q<c� w_�U���o2�1��?�E5-���E�~�WA.^��WGXT�r�w����s�<׽�l`d��p��*��6�.��T�&��-+2�Xg@c�u�Ǎ��A�tq4\�2�R�?�R8�aٷJ���2	O����4�M��<�����������K�qp�%��y0n�
(<�aw����(}ȫ���I�t�z����^Ù�v� <�&�P�4?�ܗ�MPTj?����Q�'8��?K,�[���������I�F$��S�|URQ;��֟�EՍK �;LF�蛯�c�7A6�`��\�V��{b '�!�Ӆ��F>�.�4�F�A�t�v��b�qoer��-Ќ�L��WwJ��ª�(��4E0��P�h�r�'*Ȧ	k%נS��P|5a4+A��7��w3�ߑ�۹�uh��l}�q!{i�R�:yQ^��S�G�ų�"MB��'+*X:C�W4�~p�`_n�π����80A����C==u�)	ĞNs�v�p�����m����}-0�)Xش�C����R�͇��E_Z��ohy�_=R�m7v�_є��5�+��eN���g�]���h�������� �W퍃QH�'Qͫۤ�����@5�d�F �{���6ԛ�S�Ϲ���KEg���9g�I�Jf�,	���W���=�V�����,�a	ou'�j�����%ߋ��kBU򉪃7fm�F[ _Ɓ|��癬��mF-�����<߰d�]	����9�D��ԍ珽�Nw	/ŭ&��꾯e�$'I17���.�7�a�7�,~o�s-�y9g��5��w�s�4΂�8i"�����œʰrM�>�J9�p���=S�hu��9R��^��Al���Iۇ:��*<[V�JPe٤���*	�aX�?=�7�Ǭ�������X��?�>��CO��
��c����(z8���*pyu��҃$z.	��Ζ�bF0�;E5K ��p�C&ۥGTԑ�q��M?Mp�)��n��H��A��.������[e��	p�cR~q!��͖�'0����Χ���������r�(l��ϻ׍}z/�+�"��mp��(cI7�'@{��1�Z$��!�� 69;������5�Lj3�L�O^ZڠP%��H'��9�}:����z�����<z/Rd���g�l����B2�1��:��.�����{p�uՃ:hE���I|�$��{)����
��}ϟ��`m�'����(aT�\��'��E�+m��F�Ϗ4��(L;�^��n<��P�_�������=�����d7�{��	���l�Z��e!U+���	�O�H��W�R�=�Y�;�#� �'G�1��{�~��9���ߙڡ��a�%^�k����u�p��R+L�ª	���%󌠒�w��1�f���
�6��O�D�UͬM�����!�tE��Rp�Tb��sQ�W�ꆷ&��?���`K\�$����M�-y5w���X-�	ftd;J�qޮ���U�>.�I�;�Q�����G4�f����R	9�Hki�,zfN�l���0�!��L��g�y���,�j��$�~�����0�s�VAQ~P�#*h��4ht�'n�Zˁd��)��(�dtn6b�Y�zW�@����Q��"����.�2K�3�ͷ� ��9�q��+o�vn��N`l�bt���܄���-Dݭ\�ҲR�Ov2�i�~SUGE���%��)RFCmDac)���E�O�Ƥih�˴	ٿ����)�qE5�����A&����0D����QD���!���je��;�I�s�8q�ҝ�en��h��:���qY�>d>�D��K��|)��lNvG8H�F��N練����5�E��H��0 8�0nǅpgLz�(���dw�����.G�����w��^��l�S�s�����?n_��F
��M�wWΑX�'%1�х�uX�-�[�&��Q�W�����]"�)Ti�j蔞1jv�o��,p�L�,n;�U�^���>J]����Oh�Ey	>ŉ�t��{��� �
k|:	�ׇƾ����)�Gu��jw&*�u�>����ZX�7nC�%�p������P�m��R1�.�}�.��B�CE�t.^�Ui��`�goũ5y@�:��_�%	��E�ϡ�F���&@m���F��9'��WЖ��w��(�����}'�7 '?��� R�wX�n}��\����~����.�M9%�j�a!y\pR�F":�P���� ��@ː^R��y���f�k��1S�䮝e��`ǎ�C�;���2U���~�~g�����/��R'N�X�"��wdo�'?�%y�u��ea ���������2,�AGGȢ���s���5@f�Pq�G��K.�AF��_�U��D��'g Fئϩ��˺�z�7 �5+�$�N��m��~W�H}�
L1���lDnG�{{��%� `��ĩ�RN�(%���o���)��W���{�tMu��Nz�̃9$�-`�&��Lr�+�R����9��q�K׻��'�?��FWev˲��F9�(�����ji�o*>CM�K���dNڽ�֢����W)�Z��^�&��%�ԒsbL�T�"��{��3�"��(�Yf��,�Ě1�b��.�r�Gt�B� eD�o�hXS"�+����r;n��2�$�T=r��8s���l��i���Bh3�~�� l�z=�up,���!���(!@�&��8�����B�8���#b�PH�b�kiJ«g�N��m�y�N*�$_���P /�A�w���b]1^�G3|�Щx��t�����x�Mx>������3�a�*0H�ٶ�zZ���B9Bg�bp�"A�<H�}��؅G��=n^I��jIӖk.��X\*���
�%S�]�&���aC i�q��E?b����7
��W�E�Qa���n>2�1���h��=6�{�X��v;�CG�ɯ{�N�Ma�U���:u�ÿ�����6�sm��m�V�:j����,���:tu�jx��x6-��gl�.�Ҩ����¸������P3^��/YI��3�����:�a�g�=����4%�q��gr��KOQ����2��x��v���E/R=���BW�m]0�/Tb��BB�5n��Ng�e)}K��_˩�V�h�eb( ��f��u�ɥ�>l̶��'�v���^�^�L��V����g�D��-�8߼�������_��a"璼_�'��X�I�f8t�_>̉q����l�"���u�?83�߷o>:Ί���a�i�f�|��h�y[oːjiH��A������ZLoe̾�t�g��j
99'��*�����Stْp��ue��V���d�y�a\�r5Q<ײ2Yx��#�.z&Ȝw��n�V�&G�rT�y\[9�<ǘk�|m�ڐ�)�\�ˣCCä)�	����L�4֍DФ����;���)��CIHzm�V��7$eYZ��0�|��~�gfP�yW]������2ɏ��%�{^�L���=����ɷ<=���?���Qo��}S�v\Gcb~sX�B�̲���`nIG.<��Vi�ٽ8��B��MV�0���6H��x�����ᜀ�'��%]�ɿ�WJ�Ú���,�Օ�$?r=�����8=���tQ�=g�_��;Ոs�c�w
�J<��
�;ߢ�Da�l��m���
s!<B��'��`�L����Rd�=�n�Ё�̽�M���Z��a�Vw�e�d�>���g�s;�pp�]>Й'�j�?Ej3њ�c�ZV���:�k$+]{��1SPf7�����h��1.8.tV�BD�޽�����
�գG���J�28�a�,ތ�D.t1w�OKF��	u���W�O�ة�$��톊m�z�r��W��:�QS(��r���*G1�ʎ���֭W����|�f,ӌ?B����i2�����t�V�s6����[��=��P��Mʈˡt���5�?����Ї�4�Aa�G��؄Na�p�s�P@HKI"�*<e�'�� �tՉ�BvH����ロ�k��t&$�~����:��uj�Bt��/���}X�^��M�7�l�J�U]ucU�J*�i�Q`I(�O95qU���n��^��|���c�y���%y�%ch��QtbA�v�G��6�1�k���� &j���6^���w:�>�ا�|4�����~]_�IeZ�-����7�˄���e`��^0r� ă��L�g�� ��*��y�y�]�n��M a�SR��L�&��¹��~�_����`��z�J;So�$N��/��E�#-�����2W7ĕte]�(R8��?��	�HTa��W�^ƺ�U�ؚ1��"�P���	p��n]]���H� �>�|��=��po:ڹ�r��f'�+\*t��6a�TaU��/6RlI*���}n�����C䷿z�a��	����,/[�?y�ۑEm\f#�񙙡��4jtY�� ���ުn��>�鸻T�8M�vy��1��æ�U�
^��y��$G;sI�-~�!���<���}���	�aR� Wes�S~��`�L܍�З�\c��)�WVa���z��]"D�H�]Х�U���k\�79��=hSQ��L�`�70oQzI�;�u1��Y
��%1��yY��a�RX΁����6L�]��^E� �hǛ;�\-��� ε�	�5�����f�	~_�u$U�O��lܸ��՘oʨ<
��M�GMz��1�o.������p�h�0�m�+��x`�eX�֡]5�7\��_7<�5��_�����&TO~�g#�[�a=�r��+i�Jd�5E�M��HN�'W]o�s��#��Q6����]�g��!eI�"�ȇ����-�T�U����AN?1�-`�.�O�=�䵷(4�������WƪRz�l|/��	W�d�'af�7���Z7K���Q�}C%�vؾ���~e��wlz��X�][>�� ��%�����´T$C�T��aPi�����ģ�WL���}��6�7���/ˏ
��I�h��讪�A��q�g���-yp���Lu�{k�q�H��Sm��݌=�r�/:��kk`�',�=x�8�.%=�)PAuNh	U	'?��<g�$%���_��w�s��F�����>F!����gS�6I�݀��ܓ������:�%���߅�)<<B�����\��K$�H��{���w�sހ�n������bD_��geQ�
�Jĸ>J<A.3�U�_��e���J�B��T�#&����@��
�|���\Ԭ��.i��75�1��o�V/@B�Q��D��,ۢ����i	
�� U�����.|�{|�
���a)�I���x�5\\�Ru�m�w]$�6��w�F��;���2$��s��kv!&����|5(�`�'fx�[mb�~?��
f4��g(�/�tm��w�o��+rK�B���K6�V<ٜ�����@j(�8У��gN�IA�~���u�F�SU�(��vm�PȔm�n�A�&D��B��r��c�xZ~���Zw�{���O|�@f���^��������)�b`��� 2�s���m��!(�弲"��s�Y���B���w�������J��OLH�x����jK9UUl�WG><z��k2 ��|_i�p���J�5V�\�|�������U�ս_�1�E�s�����.�\�/J�>b�y*��}Te���F1���J�jϩ���-�ͲS��m]�#1k���|�"�}�$��@�o0\��VT+]�5�:�m�y����hi�ܖM�D;_0"�]��3�������^���|h���c��)b���P,���a���7�JeR&��V�b݁%4�ΐ{Toq�����
�����I�L��w<�f����e}`k�*��_����;��D�Xd�A+h�",���E{"��7l�C��y\�'l�ju��/�@|���*5<�l����ՉB���T�e�ȯ}�7�24�g��g�!��H�G�v�B}�s�e���y���.���} ��.$�IC���Jm��V�T��;q�\�^g�k.r鴎 G��piY�,^"�zh�n��3Y�'E���|c�(�,;��;�o���|��������sNOK/K��og�%�TC���֋�M����kd@!��O��͍�'rZBu3K:z�D��t_k��!d�ݥ��^��A��T�|W��L%TM5(U)��`�͛m�L%@�Ywb�4SpZ��Q��n܃W���"��F���#O?e���g�k�Z73�'3�GU�M'�[� O�;�Ta�߯�e2��-��шf@ˤd�V�$����s3j���}J��ܬ��:��WE���$�	^���,��ךrf=G�ݘD��{�A[�T�=1-���U�.y%@AsS����骲On9Iw�LѨ�Chz��\l��8�q�`K�~r
w��X}0y��ĦeI<Hd�b(lkz�6�Q�:�5�o�E!9U���9�#r�Cl�|���\y	�%�y�6��6d����f�Ǩ���O�qt*N4/��!`@�q���;uy��$��t�e��.��Q&�d����ӱ��N�za�ܞ��H��TL�j�&~����8�Ѓe����%��`MGu��������1�}�����.�OI79&�?r�*��b��RN�U'y�gցx��K��h�З.;D��gj�4Z��,�wz;,���%�l_G����x�RC��ͪ�F��F�j�� o�̨��{�r�f� 6G3����5uۨ!T<},����VV������-pH�
���j�lI�M<�#��@�b�T~�;E����e��-ǈ+��<��a�Vw�N�<����TS�[�
�� �c�#�ް6y����B��s_9�\�ɲ O��w�aHɦr�>�u�]����v��L�9���^�`��/�22J���7�`v�WKsJ.}Gc��yr�0�:z-������UEP�:�#=H	n0��&�K��	4�L[�M4�����2sw>�zf��Q�?<�5b,����:�z�r�'|�u��N��k���|��t�>�Ʋu&D����C�� ����j�\�|�K��7�����#~�M)�c�}�ǫ�s�n��w�!�|�ډ]eΎ�̍?B#�y Ig�N�3�h�<���]o��{# V`�5'��������0��s_ޔ���2��=��/0Ӆn���?��y���j�`-_�=3_��~=������G�b�
;|��k��58LΉ	>>����fGtZd����.6�J��+�sn�&��!�x����j��s\���̙C�/��-���9\=9�(F@d%���x����	y�~(x�gJ%��� ����^wTޜ@7�ԃ��p�n�v� B�
�C�V�t�V�Z:"����S�Dtl3����G(�8h�t4g|<}��;�W�
�F�90-ݠ��eo!ޔ��N�>x�9,P�7��Fmݪ��X������:	B�!N֑�"����,�����$�2o֛����I�l�)>�𝑇�X�~B�E� ��C��]'��������d�:��"�>����ue�����D�S����P��A��ػ2����~���#(���5.�a��<�pY�nRN �j�`�&A�;��[�([��u�'��!-�*�W���F���x��J!=�[����Ca���7:Ȼ+�%g;>��ޖ��]V��F�O���P@���IО�=��Cp�XEQ����lT�
'�Ӕ��RO�̗df_�T��0����ߜ@�]X�����f��!	�3:F�;6k�Ox���W~D.���hF͵H��e��mQ�R���U��kXW�s����G�T^�[�Rp�����j��h�+.�g�Ż�6g���K�'��W��*\ϐ�b���7�^��6��Ί+�X�h2�
"�HjS'E�y�#^�*�˧ǜՂC�(E;%���9?����d��E�����H�.�x�����K�����t9Q0�[�ѶJ[\����2L��,A������XGcO�Ȫ�q��	FP�.5E��}U�o�ǟH|���� k ��[�.��{|�
(��� $��(刷�w}c�����`x��脢��Q�J���i%�늈�|@�R� '!�r�|����鸜��.�E�w�/@<�g|�s��7a�2�������簗]I�i��� ,����K�_ ��G3��?؝$�N9Z,t���ԳR��"s�j_N��uB�"���FG4���69xl�8i�"�ӄԏ��mhCJ|��O��j
��B�����V`�s�Ƞ��W&O�ث�b�g:�e���k;&HȲH��OY�K̿�r��8lźgU��C�*Uv��@9�s��$����;�ˤ!qe��