��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t���8/����K�U�[��\+r�����v.��xb��"J��0�0ID3ֲE3��5�9|�i&�U7 Đ����14�^�_8}����2l3�z�d=�����N��c��M3����-�$10ٸ����s�h����?I����|6�ކ
`eń��E�T�Xh��O�u��<��尤A&K+�4�b8������"�:���&���m}V����@7��V�'!���:�m��U���g\\g?Z�� �֛^��)����>���Ă�d���z<,��^��z��hJ��t}��$� )����w��ʆ����O/����
?��-�b����.��(X؉��e$�O���
3��+��&p��59c��A����,%�9M+JS���9�� O���|�[��4״�(B��o
h�"�Y�>t�~���(�ox(˶�q�3|{������Z�e0`?.o����=��ro>�Zʫ+=�W�i}���0���⩳8B�%�h�7��ـڊu@�fQ	�qQL����j��;����H������nث�b� �cLs9;�F�$d�K[��fڨ�����-o��ED�'�05��\�_+�C�E��t}e�k0*���B��&�[d�~��,���\��
��e4�^��,���o���b��?O�R2L�(���=&����֩+�+�A���J�R^!_k�g!u�5G�\:�L:oU�`Y�-mB��GО<0�l�(*&6mS]�b�[RVe�4+�7*�Q��>P�l��Tn^�U�I�.�s!P�*;c���p����s�(�L�@����{����0*g�
(r�����b�R2���,��ȏ	ŷ �,�J�,�g:j�<� �£)�����P�f���WN�O�&DM+;0r�6[D�j�j��h��I�����?�s >կ:[��O����;��=��5I�E�L]P��*Ҳ��o#���l��'��#���8�p��j��
��5��}���=S��Q�]�=H~9���Vr�9RT�'�T���+��ܖʭ�cbɒK&z���7�(D�ԯ�6���2�צ���8"&���������6�G����o藐���z��,>���(s���L1W3"$}��c�5jU�G�`x�� ��C��*(o�R��Eũ�G����>�v}d����775�\l1 �q����
�pB��#�Gv'I��c�Z=��{�$�P��Q5�F���� �����2u�@7�{���e���n[��8Uwl@�I���hQ�z\���*���(��)��yEl'X?���ǩ�۪��\��I��a�"�b�U�&�G�y�X�Йa(ԯ9$@Ky��*�0�eMHDЕ��S���e�?d-c�C�*|;;��f���;�lݺ_��L(9�����w�����N���5ʥI��<O?ĩ�Z��=0�tlS�}z����*�!ܪ��}���L?���G�y�����t��ת��y���Jă�,Md�3�@,b���s罽pX����"�XD�h~٨�|�k��`�J~��&�a�p�&O�YuJ����e�q*�QZ.ʆ���D�#���m/ �s�&��V~Fj���k�/�ճ�l +��.��-�Ɋ�Z��"E��1��fm�k.��M��?�8y��T�߮�N���&� %��z�^�{4�y-H7G�;ϟ!QMɹ���ޗ�*�C�3�o����3)�(&���$΋v`�ޠ�Xˌ���ܠ�b����^�����\�l5������4M�}W�s`��P�)�Z�#��+V����/oۅ���EϘ�H2	�!)�#�^��P30ew���9��Y�jɺ�5�|{9�D�^�V.��?�������d��~��k�qI��*��G�	:��+nAl9f��/
�|5��y��/[�+uq��X̯�޼�B�3�?ў�̄����Z��;.}b�U�g ��?����<��Wn�7 �[�	�ڄb��{��~�+r�TPd�'�O�����4���_֩����m�����.��20�;�G}P�� ��H[�ۨD.*���]ܓ`��e�_�;v�6c=N����;�K�U��4�FLD�fO�fo6~�&e%o�b�������!���6��8��⽨����RMe*~lȌ�SV1� �($�#Ϫ%�Im�2�C�O-�wAs�jҚ�g�R���S�:�PC��gvK����=W�Tț,X7�t�}����Ix���bd�l�:j��\��.�W��i��Q�u=^��g��2��q��?d�ɫzu�*��"'��J�-�>�c"���1������k/�l%�^�@nfp: �"��ad�`Ծƃ����D!���E]��u��B���8�B�z��E��~����ۈL������g���5������u�.�W�ڱ[����&C����/ʁw�T}�d���S�� �4����r��XY(�"{A�r������H���'��ǐ����lG�J��P$t^�@j�(B����X�,�Ǌ��S��_=�:�*��"��L`N'�]�H�o��댹D�6�X%����S��9{�W��H(�Ͱ-��������������3<���u-�T�\-fo+Ui�����&=0����c�����a��D��ё�J�s���*s�6_:)�K�D���[�I���B^g=�
''D'�|�rmt7����e�_�tm�k����o�t	q#���U��dn�J�3�NN����:X���5Z��0�a�gF�D6��S�j������Xm4r]��J��C�I��Nj0���,��$��k��O��`�dg����)lOn&yʑ��,���ҵ����*�59O$�b�)P�e`�S�C���$M����&�£q��no7B�9fG�; 0���uO��&�?e�;��h9fӏ�t`gY��)ף4�ʹ��=d�u@���s/�Q��nO�+�7UZV\9�)ň��
7���������y�˕��EVA��5�]�[f�ow���%y��- ����OD���/�6Z�r��	`���p�fc<�"�@^��6�ɵ���!
q���D�d�FO�"5;1��7�m� Sc�e��D��`�R�bGH�͓��1՜S�1+�+	�I.�y�����>�|�3B���̍�n�-]\���������1���׫�Cz�2O~ѷ��Z�����ᕨK�k��; ����_7�#R�E�x���s�o��p!����a��8G̳=dKdX������r��2�$�[I{����E����(���
  ϝ��B2��rs�7ӱHɳ.	��Eث''/��-�-K�������5��v��)7훋�	g��f�<ZGu<]嫪ZuN�~�:��%ڜJ�U2"�SW�YmX�Ƀ�<%��4~�ŧM�DS���E�<Lך/^�Z��.;"��!�e�9�2��ٮ�IC���K��j��H�Vi˺VZ�)�Oes˨r"w���B\~B��8��������
֑]A(oa�j�8׏n"��]���ש�H��h5�$z��4-ם�7H$���ɢ%��;�Q-9��bּ��T;Ӑq�ղcSC�9.Er{����a�a�:(�a��f�1��n5��ׇ�n{���!:�)���Xn��x:�`4]v��w�w��S#�H�Q�whÓ�%!��)�]�V�8?);	����� �y�h�³{kml�e�v�L2A��'�Qء&\�:��o�QF��3���;u"i����ߣ��������j*�������3�oP�o`�7Ә��u����1�RBxK[b�O��iӂNU��3\G�{{��f�D��5�~e�QYK�<��Oi`P���ЩZ�� ���B�ke�#������-׌j_�Qk���Z�v�ѳ%{s��q�������R-2�U*o�ߵ����P�_�M�ط��m�Ϸ�,�'?��[ˡ�dw_�H�U�A�{���m6K�\R�L���/��M�E6}	�29���}�K-��p�d��>�X��W�g��N�"���3YUBVU��#Hnٷ�w؅nE�H�/�2�k���D�ʜ�U�����p����1�ԩ�F�{�,�\�%�pѪW��@�2���6�/�}R��hȧ#����N��T�!�8ؑ?]G*o��CM'�Ҷz��+�b0�F��T�	�4 �MG'4=>Y�_�0�$(14��$t���U'�GȈK�ډ�!b���Q,�Ą�qV.в���"�:�[Y����^L�3%����yN�J��ۗ9��ɝ$8�*��1�1�5"<���+����Ȓ2~���G�
⼚���l��n�ϖ#E i>ٰ-&9:3����G��/ļ��r{�	��Ov���vʦ�m0G�D�"מ�(s�1�s�
��C��!�wR�$F�+��a׻�|�"ˋ!�JƲ.�SC���V���['�0M����hu3%���h�A^Kgz�A2����S�7�*6L��8�@4������:�օ�j��1rAe5��Rھ�HD�52��Ƚ:��Pź\�\�N�e��T�r�D��e�.S%-�*:bC���5�D�~��4�A!`_������S�XWv)d�n��	r��&��R=�'��?��ΡG����u���H���{:pe�����搣C.Y*�`��FT����,\���áS&5p�/�(2h_֍�Bq��S��g��2')c,!��R*6���e���"wb��I4��bM}�t�_~5#Q,�V�ܬ�=�{�I~��; ~a��P���I�5V��'I9�X���o�&q��oU��W�>^�X�8����D�H ݈?C��v9��J0��t�jQ}��/�>2e)�v�3_��n�A���<����t�*ݚ�ҵ���ن�9y�Q@g��܎ՙ[�=��E���R��Ƈq�g�PO�j]�T�X1�Fv�vN�����e|�A
���գ�nRM�NV2r�N���230�o�D���-���Ӊ�n#�ʲ&��Gm�ֲ[�:o�Q��+AZ��D���׹�I1^I'�_
�������"� ��t��B��9V��E��Q�{	���\X�KY��ﺃ<U�oV�"ډ��I.��$�1�(0��g=p��}G���@r��FI��qԒ͊��i�k�\��b��P�M�mf�zdj�� ����9���jiW��S��K�b���^�e�,�����YڠW�����������K4���S���t)�x��Lٖ�Q�S��a,�W���F�Y��%���e%�ԜA��+n�
î��������x��ё��O+X�PN�f��I�������D�
�s�a�%��4R��`�Pd��-㏥q�;����PV�c���W� ]����Jr*���+.�B��JbH($��/!I��B�e�J:��ŚE�f���`�A�7��w� Vˊ�{G_�T�p@�/DN���$|�<��BB�J�b.8�cڿ.��]�l?�u��yY�o���8԰t��->���S�Q��@�<�~�E�=ޓ�T��B40GaӪ���(y3���IK���*������=�t�ǉ���2���g9B×�R�T�{҉�	����l�C���2g��>a�;��2���Y�4�6�){�[/��"M+)jTQ���m�W�{�A%��y9�CHd8'�"��h�8b*�ی+d���1��ɂ�K��T�W�hk��W����J'�t�sh��Q�[���@��r.��\he8�G.\���5����՞ry2��/�|#���ԛ	��ȥ\������i��g��&�`��0��ʗ�>��Alʒ��� �JA���)�� r�E�*����I1�RW�%-���>nX�RY���\�GF�بã�:u���V�w{�A]3{���}�R�q5�Ѻ3љ�>X}�3L)��PJI�*(�7�>rA'y���9Y!�mQ$�xk-���)g�A��ۍ��*z��7�
�~e!g�]}����j+R�8�;G3V���'���bd4o�o2o��	W�ǌ�he����q�R�.v^`��u�unw�>:�����3]��G�x�C�֦�O>e�Fx�u`����㝱�d�Du�/ ��H�� ;����1�O�25�-���7?rJY\%b2�_����ضuC�A�.���(��a=�L��5��_��8�,oP1��׿��b��8,��O8��wt58-�
E�t�������t�F��M� P90�4�@���������<����vNC[AD��٩q��ip4��Մ.>�?�!��K]0M�9�!��<�]���a�	� ��`���'��ZP;z�y�21����%5�Z$�-��,��q�8����K�/��L��O65��3��V����<�XA9����⬛��k����~�����Ac�̵߇qi�Ү��,)�-�Q�d�^B���d�m��ժ�܂����3i�DM�n}���D���+Vr��se)�n-�ũ��S!�O|K�^�^�����	,AN�4�9W� ��5��q{p�Ͱk�Jm�&��	��#��7h�9u��4'=C!|o�K禾3d���'�?�7���.�u�`#T��Ɵ8S5�o�3-��R!����7Yb�M��������vq1�J�P����X�En���UJ�Q���4d=H��L}�<XZ���gI��)Yuftd'B�@O�؋S��ե��9ځږfwx�)��j�O)a{��ֶ�U6^�\k��D�ȁ�Y���<F���׼~�y|��c-���Y�m7r[��W��Fi���i�v"��h${��ELV6U��~������A��g��i�Y��LX��1�1[}��cs۩i
Ç)n�뱕U����yu��H������~<����X�u�"�R�%)9���_��c�#�j�j��{�e$���\���a̳͌�V��U��������W=N;��ȥ���K�=ס�������8�@����[�ak)� ԮV��Z�nC�����zP�>L!����^�@� ��7�����10�g���
�%l �j�K�&vu�7�O����*�Ә}��+�� ,��yc�����f�t{J�����T����|/UxD�zn�h�[�����O'f*�i-������FظWAE��4Tm,���zXH-V�ux���V��Y������kg��^o���$���trRt�agE$N�G��� �����?���[�϶a��ȚZhBr�4 Ip�f���k��w�A����]�֑�
��ѤMx�J';��b��u�4�$�\�*O>�N��L�<4 ���f��,襶���US�����E)~��'��	�� �l�3.rG��<�\�|�^��~�ۏ]F�N(�'u���XJf���v�Jta��¿/_�
ܰ�.t��6����(� "a�I�n�-��
��'P�����G�3���),��gA��4@�St���_���e�?��2����E�p�o6���KC���{+O#�DP?�<g,����O[8�-����4�[_�>�IK&n`�p"ح�q���wM
60ęE��e�Xn�s�����7�ppI;���,�m�0Ț�bS�d#�%w�\09��������?���5+�9M ����Ƞkଗ)b����8�]q|B�N����$Mkc�vI$�o�bɸ�֤�wo�B����2�r �ŗ�<�9ނ;��%��v�~�� ����u��K��3|u?�Z?��A�jH~�Kue'�n�1�R��lM�9�9%��C���Q����,up��T����#I��[/���C�X��)q�h�R0�0�s��G��shq�T����>�<��H�'@���Hi�ݠ{W7�����-aSn�����T�>�?B�7��%8�n.dm$��!.쇂�u�����a^I�Ĳ�*��e),�C�G�� 7	�����NA�Fq5e���"ñ�\���?�?�c4�n�6jJ4����� � ��9�V@^���t}���Y�7�r݅7	O��)���Ae�M��ff��
�����U��})x����7�HRG���O��c�Cb`V\,9S��Xd���S�X��\ڹ����&�8�d���O2��`�VI_ˍ�Po)5����Ʋ�J�}�}�2����Bg��%g���Dө�+���,�;ء�T�9�IaP��O��j[+�)%� }\/6�4�Y�q��Լ�#KY�~�Cw�L"�PM���^���g�.�fFFQ�{̶;��>��4���OU�O��"��f7/�}R�t�/[�@�K���(���b����Q7����:ߡ:�$`��{Gk��Ĩº]�݆�z"�%�`��$b�6>�b�[�&�KV��`�	��H,���dsu>�$�XN��)���l��U���>YӨw³�4����yo����C�
*�B��=�y�3�[8���q����Q�P�o���=��d�T��fU�R�vO�6��];��lM�R�NΊb�%�]?
��¬���w����z'c�y������K�w�����!�x:Rn�-�%F�e'����|n7�Q8�]@�F<�HZ��~���BQ��zBA���'5�鹤���݁O6]'&ʁ̺�w:rv�r����c�&�]���w��iQ޹��>I6� 6�ٰK�B��6I��h�u�~/�D�'�]��&+ߕZd�\��,<��7^n�'�ӃL�P�7�����_|�Nv�s@S�ҹI�Ƀ�LrɃ�ֵ�_͒��ݒ�~��=�w���;3�ʸ�M����V��r�x�_|�:�.�;y��K'�VN�Cm�W,�<M$|��Lh&��x~��W6�Q��w�[�20�FV��sN�����PP$Yj0�H)+�U�W�Km� ���X�5б�f�{R<u�}��L�t���l��f>� J�RZP�a7��9.K�]Q�=Md�|��HW������=�1�M�L��v��	�m�I�`̓o���J��n�zy=jK�lkS��^��,��K��'ҥ��e��׾��H�5v
a1NX@ԡ8�.r>,H^�E
ib	7���� NKWo�ί��g��ޞ8�G\ؒ}��$!�.�f�������',,���u�����T���H����&�N�l?��>���`�Ċ&]�Ի�6hD�Y��"	xe���.�-�ٴ�۽bj��{��c�@���C��$��]�5+��N0Joi�2�QbN��9���i�?LG��\���F`�f���T8{		�H�g�����S�'�T믇��{V���u�f�
}/lE�$-S�bo����6�(8ug�&�0M産�ݨ��[����;�k���?w��!�������Eլh��Gy(+)@C��l|,��-����u�V7ت G��3@Ex�rf�r>��%��\�t���9?�v�@����Ǿ��K����U�v'�O��!�'��{�~۞��Y-x��BT�B�
S(t2�G���-o��䄮B�/\��=p��C�$�� A�iםَ�טY��Ƈ�֠�29��dW�i^�R::[� ���Y�*U��D6�zsx���l�:��/Nerjx?mL�e�	�����N��)$SfMKFW&�$�`����I�F$<�u�1y-d�.���0�m��
{v_>R������j��A檲��J3��!��8���]b�2�ą���X����������ݟ����4��\'�m��~�ʟ̑�a�0y��9�A��_���~QAieѰx1c���$J|%�Q����g|�ʘ�0 ���y�{}P5X�w̾�P��8ݨB���G�����a-Dǳk��A�{M�.���~�_��G?9H[AP�G6�>���z��;�&8��^��� ��F�:^ZJ����ƕ]�Nr�Laɩ)7�U��/�#0\��«H�Ʒ?���ڀ
q�/y�VV��m������E&��C��ţ��f��v�� #��'W$�ɳ�U�*'��G%��Ґf(��O�vX8�.�b;b��a����b"��~��d�Jٶ4Y�v-�x��,�NU��a��1�l����L��+�km��aɖ�A��V\ܴ��W��":��b�˪�|ۈ_&�����s�,]/��>�𽍤���f�$�ߘ�>|�?��e? Yp/�ax>�߮�}'��U5�x�4���nN�\j��L�5�y�u�W�ş(�k
�|3e��i��M�!���{��`��a��{>4��Qo(��38ݬ[0�א�́,h�	�*����� y*Dc	^l�S4�К��8A��FO`�Ѳ�x����ˁ�t��q{�fPJJH�><|  �Fp�z0����T)�|��P�.�0�q�0�z�\�@�v��M�y�����q!@@�`CaG�b��@;���C��ӕ����\�-��E�br;�ܘN�N�sn���-k�2t�/�G1�iy�͐��$4nz�;q�]�-E3��p�=~�筍-�'�%��L���R�S������7��)d`�K]X��k)�'�n#�%�L ��O�"��L����B��~���z�W�۲����B���ib~�~��*/i�z�Ώu:xZL��~l�s<qxP�F/�S?p��0=$�X���A�`@�#U�C�FD�r�ή��3e�0��·%�� qo�^��� |��M���Ԅ�-���&�m�U��v_�����_�ˎ!��Ք'����4P����޺�Bƶ"`�
~�J�����#�,�ݮY��b��f��t(񈂐�CS6�ھ]��8�Iu�k[�	��e�b�d�3ѡσ��Ҵ������ȫ��nz;���̶&�}L
5"�0�)��f��8�K,77�ll��w��9
�d�p�b�ЮI�r�B�Uե�u_/2 ��J��q���>�l��63 kFwf��%����Y���	�]�/��W��+3{D��7����3�澉������*n�Z`�&PE2�1m���O)6ҙ�\ȱ�)p{�A=o����֟E�r��~
N.H��傤����Ϙgg�A^B��H}g���Z1;�IӤ'�A��)���F�Nơ��A��`�G	��)�Αړd}������,��g����Y'G����C�:��M�jQ�����Ɂv��T���)�}��H��L[ʆ˥e�n�ʣ��)��C��%x(�WH��Ot1��9&�@�hQ~��^x������y��@��B`֭\��-�iT�O�A���r���0�~����1$�)�������T�190�f,=�UO�yȑi:����d:+zɑU�E�٣�4�I}�	l=���R
{h�:E��7�]��)�`�&�����lr>�R���֑�5����S=��3���N��h��g�b^E�K�� r3�⎯��^�7}JB�v��+�YWa��U�ގ����&_Qj���u�PD�ӫ�EtG�R�<Gv��D�ԽT�e|eh]�3�u���
����m#��������3&�/�Z�q� s�V��k(��
������$�7���\��k�ɏI��Ng	w`�?)1|s��E	�\�R�����l��`x=�rN�e�ο���TV ��\�#�t2�s�5w�u�� ےD��_�ٓ9-���Ė����w�b]?[eB�Htg�2Ϊȶ]���V��c|{�)��C;q߽�ފ���1���������_%&>h�#6KwY{y����!��G̷�l�gj�R�:�ÿ+z�Yx8��rݘm���d������77D.�E�ҿS��Joϳe�V���rׯ�Z��F�K~TNuDcM�B�-�w�dA�R�˧_2����#:b�1!ڠ�_D��r��� i�z�Ud�=���K۪\���v�&4+��	� RxL|,E�j�TҨ����Y��9-��x��É�1ňe�A�pf9m<F�L�[3^J�ˆ�����b���|���8�I�֕B����P�C*"1������]Q,�ֱH�W�D��L�ʔ�բ�D�Z���?),���-d�d��ڠ�t��Ts��Y���6��<we�&�;��3{l����pW�?kYt�3/�f��[��'��L7��n�RY�����A�N�:�{�!S�ahB�`�)���*��P�VD���R8�K���V�Oj�|����~��(x�m7]���S�����s�""�;�Y����{��O�
c�.-�<Ρ��.�A^>���4֙�4����l�cU�[�GQ$nB�[r��p��?2�@0��He��1A�\S(f�R���tX�U�>�:�)cG��@M���9�=���@Ŀ����WkJ�4µ)��7�'lT��<�b:A>�
��b���HX�z5B�qc�}z'�S����:�j_�Z��52�-��\��`b�v������o�К)@X���|Q�� ���w�i���S�s�����d]��A#Y�0�4�2��8
��a��X���b@3�	��;��i��y��zǉZ��l�D��$��:v�v�7l2��ݎG���a��yk��ʎߤ���ɬ�����l,4B��i�
YS}���k�� �-�Z++��M��Wu�;�1{ش�L�PZ�T�]@����9�~��j��=�Ti�n�P�ј�a�s��$���v+i.E�0�<��$
X����l�{\:�D!qPAc�ic�diP���/V2Í�j!�;�.(�S��7m�˚�R$:���̽Pz��W� �q$�,_Je[�'(c)rh�EP�n@��ʳ~Ĭ�k�l|�{�Y;�8��!׃,aD�[���fz�A9�7Wͫ�[pr~
���B,�F��'��
�aIR�Ѕ