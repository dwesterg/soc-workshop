��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�ʖ^��
ccֶ����$����{�����m(m�P���yĻJ��!Oz@����Lʠ�1X�i����i��� O���6F��Ǡ*��<s��T�t�b� � ��ƭ��݈u�w�ч��w��(��Vf�nT�WSu^3 }G�1�� Y�mƻ�.�F�[�6_�LJ���j�p�8p�U��Z��:����(��q3~8a X=©�������
1�R���!�t'Jb�Z�NI�D�}��G�|=�A�a�2=��M{�<�� �����e�?r�d��4Zү/���<p��1ԃ�����yA)(,���Q]DbT1f;{�^�8�U�4�<�T���
����O�9���:�$��\�}=WN+���F1��J�V@�	�⥡�ryѶ�U�1*ʂ����<8�m�o����A�t� Hh��q(�#��&����b���i���X�mS;Ԑs"� {��V�y�O㡕Z���Zid&+$Ӹ���$.9$�Y����G���0����+�Yأ\PFU:N>4�U!�v�˝��ށZ����?�X#ubla��x�R�~�a���mr,5��}bHҕG����?T1.u�*zh,B�I���&>7�=X�9·[g�����'`PdgV>�?�#�m���u������X#\%�X�l���GxH
'�O���� <�J� ��U��Bym�ݸ�������ð�����IB���ҘD��grV��|6���Ύ�͂�˿��U�r>X!gzP�<��>RlΓ��j������N�-$�D+^�m��4����5m.��:A&r	f����OY�.�g}\0_�i�-���g�T�v`�N8l��=ܚ<����b�+�HZ9|о[V�8�H<>���.wD�D��t-^�9Ǣ�r�jS<D� (�M�p���J����z���&$�SS)iy^�H���ٳ,�3X��;�#���1��m�n)H^��3B(}����RO�\�I�x5��q�b/�[�!�;�3�s���=S�xpkoF���_7ҿ,�˿�.&�L�5��7=�	���vܓ�ͷX���X�}�2h����.�A��?���UL���:�X&��9��)X(�ߣp����2�h�=��n�Lkr2z)&�L��?Rv8|@Z���=��V�0�G��"���&s�z_r��1��
 ��e|`��SXq!p��ݞ��
B�.�����Bo}A���M�f�>��(齻+��5�hA�ۼ����D
�j���:�u?]����-Z�%C���v�0��@�d���:z�*��]��</��icGq��[��F����˃�!Ʋ��2��������e�T.��[٠�пR�k��űR���j�0R����.,qk��iu
"�9�s	x� 6E8$�l2~��fC�9n�B��\�g��~8ן��@��d�ybU�n�Ԏ�,UF��:�#̐�VL=�/w���nk�e궿7[Q�r9���>����o4p�'ٓ�����ݟ	i��6���\��⊝Ԉ@"��vzOC�<���ȏvE�����o~V����!�f����joLs~�	$�Z��,g�P�烔�DSleEpi6�"�x��f2��SO�T�Bc�d*�`� 1�L]�)�� )��5��	�j�����)S
A��d�`��㰐�bw&���*.l��)�i�4�;_� K�Wڢ�W��qA�o�A��ƕYs"7�F���i�3d��d0[I
FU���.�aa4�o5+G�[���l	��E0/錼0ZH��U�Vv@�{��j��k@<�l���I-乆���<��XPS8�"{�^�Q�J/���V�ܦ�V�E��� �H�9�ɨ�V�m$��jL.q��#��B�O,]�=�S�[�YW����2�~��n�1C�?�&;6���/���4�2í�]�]h�N6p�x�ް�}R�o���>�ME����n��,�R3�5E�p����z�a]�kv�l��'-�:���McG��h��<C���T��m��v�T�5*��_w�n�w�B9U��5n��(�|u�WC~$��=�Z8Wwi�4�S�T2
�%���1��>G��~g�zL�B������-i��Ff�S�G�5
`$��G�O}�\Ua�9\�<��޾�FC�8����̝�_��w�X�3C%1-w�t4��+��G��`'��##�&��������&b{�r������LR!;N\�8����AKbt����r�K�T��s=#��{9"u���G(�4��
ӣ{����Ƹ�|R73k����J���\�@���\��o�n�ֵ�j�,<QN�_>�
��e�򞁖��z�Z��O���R�K� ���+	��^��b�E�m=|�����nI&�$���C{6��D��������覯Sq�{����6O�
��I�H�,�R�@(�t�r��eS��h�4����˒�˫�K���P"���҇�3���~H��7�[^�Go	���17�����9s5ڿ���	2z�no#�!�z��ƃ7XHr��c_R��:��d�h�T-!�!f>�pG@�6����n	2]�²zlN�>+��-�p���%q�^b-r�/���������+� � �6�$����%��In��UE��Z��f���������c�)�r�lc,s��ȫPɢ�+�eў��w��a����H%�ի���FUq)j�΍���`�p�v��`4�9`�y[�^L���瘋/��8<'߾�����)2��A�W�W�s��m/���s[�D�?�Am�f��-6����n�~D&u�ӵƂޝ ��S�r`t�ߐ�㘪*!15��k��u�p�i�[�?=�c�_<�[VwFl�]z?;�հB��n/��z� j5�/�t�x��rO��(��S�N�@vM�ԭ��'�egTꕳ@�=W�PdKE�W��.���|�h,�V�N%�������O�������#�U��eyM�P���wGgax�ϳ�a��pR.'#��e�\�s2d��/t��s�<��O�]��=r��} ��[B�Rh��A�%�
�rǏ�O�>Ycs����B�ds��fnJms�֠�c|uH��^�A��V
� ���ÇC�IRbx"������oJ��tG$>:�U����~����h�]����9�=��;JR�������_�Q�)kw�	���ݐ�4P\JȊ�8����PIn��tp9L!Q���3���~���D��q���N?��Ψ��M`�M��~����i���}>�%Q^��i��L\2��{[j$y��'�/>�?�(,�ʜ:��E���S���SZ��~,\���;3*7�z��,I�U͝�7,�	������uĦ�#��cIM��]�Y�Nx3Z�x&��{-�	��|���K�Nh#ϨH���%_wxF�Ӿ�����[�7��/�t&%�����_�+�F�y�W���C�i��8�-ل=������0��{�݈US�S�J�=߸��6���&Z�:��j"5fMU���g	hȩ���B𹱨�؍#'a�3EPb�#�ts�_|�UE
]ࣷ�I2u-o$��xɆ(l��� j%O�N�
�~glc�0J���t��g��\7��gn���v]"��3\��z5�%�R�����y��m^*A>D/���@<��s	J3��56�-���9%����>���<̻�l]o�Y�g��Ǜ���+��s���z�F���	Zc������P�}U��w�Q���ʛ�T�v؀��$���ڕ�*Q��" x+��G�J��c Gh^Ntx�l��iϼ�`����H�����*����d7lp���	�Eo�q�����`MN�����������z�A�s�;��;��>����u�yh8�����q���]�a"��vm�}wȤ��;��j�����:�|a�by&VNE�i~��!]
؅�].~dl&M�R�FFɨd��kd�עJ�^�Е
�X����a\��
!Ds~6kv� �x�n��Mل���U�&��}������E��c&�d�:&cS����5ꆈj�R�uYi��3�Tq�� F�͔�_��v,�0�<)�"HG_c���Y>㎛Nw��'��o j�=�5���{�W�(UL{H���.���m��������blsۑ]����o�X�=�z�ݤ����ޖ�9{�Ԏ*�Lm���q����jn�������_~�4K�7��M2�i��e���S��P�#�co6~[��g���%���<X�Ħ��+\����B�v��ޒv1%�5�I���&�൙����e�Ҍ�k�r�#P�/��|��pm�c@����t��oU�XQ��Odj+ ���y�=����\��7��q�*hvu�Cr���:�t'�AB�1��]�u�'�i�7E��`ӟ�޽�	O8K�*.�Zq�B4-aC��ƒzF�B0 ���������*1{E�;�2����ѝ9��<��.�Jxg�MR� _���%7��Q	��X/�#9�m0k��Ǿ �0]��S8�jw�V��>�q�7d�^�Z���}�#U�m�fc�\Q+e� �|F@��].k�-�褉��c}|�;r�%��k�ߜ�h��cK�~���o�<��ZB7��;㊗�ʋ��rI�kfq���i�8��.����������6"8�.Kr,*�����j��#�xh�R��?�H)u�ˁ��y��x6�'�v�?L��긩=��ɺMg�I�68�	�^?U��"��R�ؒ�}0������9�gm/tܽ��8W�y)�6Ϭ�ph�w"�ٝ�p�d(*�� �n�ld3�����Qm�:X�7�s/��0�gQ�z��9����GQ�5�?r�ƕ���q���*CM�h��沺���JQYu��	t��"��ҊѠL���e�A�)�H���=56G-10���P-�ʑDh��6�np��A�	b��'��3SN'�`�R5��m��ٜwu2E�ei�ʎxJ$�`9��z�@H�x��a�8��FEn�Y?�ZH��b�
�4�m\��Ov�t&�$���[E0�ȂMC6����_�v	��G�1#c��)��6�Dd�^,�������z�~�I$a:�6�{�ϙ�6�����>��=q88�`_���������'3%'�U��	^���*bsUJġ�EQsgc��8?r��wa�J��m�Kd�� #�{g���Z��k4��u���+SRl�{�PV��5
YK:ѡ���Mō������2pȓ��#���o"ܴ�=n^�w9an/�ʹ�C%��,!��x��c����;YW��^$<��=|y�5�o��#���5�-��������?J�.
b,r�Tߦ�H_�6|2Y�_�̿�Z� �B�X�t���OF3��,xq��X�X�q��mPV�82�=�*��`ְH�F���=�A�f���d�'+v��h�7�H�5"�$�ϒ��H�<��z�]��`�OjѤ1	���Z��)Ej�y����| ��_(���a�ص��}�eU��(ӕ�#)��ձ��0��d���?�������ܢM_�+
("c���������f����?7�w��.�������\y����Ӧ �A6�q��ႹL�\ L��e��R�J��á8|��F�F]��K�u���>�y
�����kr���r�)Nc��W��W���B�b<���+�9�5Uqߑ�ۘ���h8�0�d��	�'o��k��<U�]S���PIy�X0y��\���h�oS�7˲7�#_�p��4l`�ᘖ����NHJQ����,9J�;iӄ�Þ�'T��3O;h�ud�7��{ה�G�0_�!>/����?�����_�ĩ4@^���JH^���X���Ν{l��x�uR��/�������W����;�{��I���_��Ļʕ*��рg�� S}�dp�c�]�[[�-��K�x?Q��p۴^�+�Ǿ���l�