��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�,(ۍY�Y^5��=",E����VF�?l/�YH��X%�A�E�	�p�,�?�$�d����e�Tv��!P���� �a<s�����uq!�l�o��Y�Zw��P=�ī��ᙩ0�8�(���n2�*��k�oaa:;�pw�/k���<�2,�H�k6$�~��r.b�\-�r�t�%<m^�]��'a
^�#����}hr�M�X�6�w�^Ֆ�m�s��Բ��~~�J��1��U㡼�=�zF�O傡�}x��Y0)��gS����9�	��1Z���cb�
��lo���c�g��)��+����3T^�Op �Ï	��Fd|OE�󷙜��P�e�L<���Q2�*��'����4��v,Cs.E,��q�Q6��k���� �`ؖYnz1��vl�$�945�L�r�Q��*I˃E������z2��.�8G��
<��L�vΘ�@u_�%�c��a�K@��w�tUA�i0�+ʝʍQ���_s�1�!_1E��U���o��T�F�#�ft�!W�k1x�H�_�~�&/���3���/C��f����Dq+qt=�5�!���߆u�)�W�ܼٟ`K�54�q,��y���M�H@2
<�ӽQV*J�H��}CL��'�lW�+��2W�"w[!�1��X�S��prU��O%������hI�T���<�Ȇ��{�K��~��=�
h��x�\�~LY�l�M�����q�x�3�b�u��b�rNP�c�cSS�-d�D&-����Cz7=����@�����:�n=Րs肹���S�	���91�c��s2[z:�P�قȆ[T��v�Y�'��98��N���9����{N������qF0��m2��f�6�ȡfސ��8�f���X�Dj�m����D)��Bu$Q�I�� A&ayk�P$���`�)R�dm�I: �;Z��S&A�V�OGz~��^���U�Ǳ���#�ɯ-5��������4ֿ�ȯ)d��Es�!ŨlM�)/f�<���4u�ɜ��Pg��_������J1w"�$��<MfZB����yz���CǤ��eݴ�E��E�)�Wk��B!�)��r��7�K ��-���k4�^H[��$]��1�)�2]������-q�<���؞��D�.�gkKP�����K�a�u��}�6�q2�)�u2{��n���0�����On�n;vt%�l��L�������]7��b�}���v@t����<%&�7,s%R��]s>��]�����a�ԍ~�CȲɘ����E�؛c/{�jZ���M?5��ef����(��5W�.��D1@/S��7+��t�� dl�����7a�h g�E�v"�y�1����0o����X&�냓�������`i�E���5 ����@�$),�Í�� 8�u&��BP�b�xϭU+��E���g&����3���F���{��k!u1���l ��j	<�J�����x�È��� ��f���0Շ�?!_��l�pSe���k�2���|� �o�I�eA�aAg�L�_�U��	�joi<�oi-�#�4Y,~z���s]�jq��Ӄyۡ2�%g�"r1���)2���AM`����@��cr*�I�I|��L��N��ĕ\�Z�3�gD�����0H��Ґ���^z����&��?��Bݭ�汍ώ���yLH��s� ��=\xb6�n�t*gQ�Bey��UDN?�;yѓ�Y�����@7�'pQwڑ�yg���й��oWv$��!�.+�=��{x&������"��M:x��a��}zn}�떚��k�]����0wW�V�T��Ҡ-�S�3:�j�����]C�]�V �0 g&a��_���X�Ńk����Y)��W��ؚ�|܎!t��,Ed����P�3dߊ��yK�FhV 
�>a��c�U����Z�O-���n�:����JO�lo�1ы���.�ɶ"jU }S��q�"���1�yA�5����\̎j���|w��������v�����={.���m���U�x���Cpnv
#�q��*��s\C�W����&�A��A�����u��ၭ����ˁ�m�z JFY�`���X���}6�l4��-C��%m[�5E�Es��N].��^�t���P�b~�<��a�����%��O��d���.V�}��a ��>����Vt��U7���O�l��� ��F����x�诲�cM��B��%`���faN��M�:OYZž���YR�R�*�{�ΖT��o��(��;�=���7�,�2<���~D�����xȄ�~�f�
x<4L�$l�T�*C+��IF��ɩ��.&���9f���?YIj7����,[�/�}��V~�6[CC*y.����:-D�Kr��K�i�5D��'�&��\_�矟~!�y%kM=F�:����|���F�
ƾ���WJ8<P	��k�4�Td�x.@�Tͳ�/lԣo����WO�W�,޼���nhP�~%���>�F��WP���(b��P����0H-Ͳ��� �sD�-����7��c,���"\*2���*�e�B�5\���B��	�e����n_���i}��7ٜ�񺏚Z�Cp���
c�%�<v�?VoOo�����+�+�ʶ�g�(R�-՞���Xw�L2���G�/����K��������Ǖ���c	JI�M`"�^j�ol�y������IX�Ld^�A�!1�	��N�u��8���aB�"sy/�-��>���K��r�$�RPo#��8'ZAJ�&��˺!��f�%��@��h3�>q_��T�4�v\�=�单$��T�� �_�i˅C,���t�g�$�B
�g��?�Ʒ�K�����tj꺸*#P�]�,�H$,˝1Z i�0��̆�����V��� ��J������D�F_�<`
5����rNS#��C�)�� �.�&�m2^fkf�f�j�J������*�o`�1eyK�!�P']�O�uJ�l��D ��X1���Io���� JX�$P�F�zfpԦG���A�n p�RL��țvy.����y'���׹Fc:ިJ��HA^��q)�ԄكM8uǠ�RCGd��O����ݿ��ԃu��I�ͽ������$�+���W)ˌ6�oPB��F��R8�VM-�Jε�$�1��0�PC�Dp�u�nK�h;)|� �uky]��b�	q�gb��P�yH�i�5�}�TN׾��	�-�V%$ zdZύ
�I�B
�nXf���m��$���u� u��C���6c�� x�0s��L#vu01� �NP��1��H����X2��4%U�%0%a ���l^q��ˏ���Pi�d��E�iS�\�I��fE�v
7���yn�:��ȿ�gs�Y�~˸�4��R�w���)"���$H�����:���%7���O� �s��E�t�-���@7�fQEѫ@;��@G��Hb�z咵�zkbd2N3v�-��c���[�?5���(�D��JTa?[5{���'7�[.ҹ��V�RӖ?U���D��������R���&���.�("���R1�9���(�'Ó�QAb����Ed�6ύ�����R��Z=�4���@N�+!3������#�IvT��Q�Rom���������؁q�I���6�oNԧ5�����,��?���v�[�q1��M���bAP��H�I�Jȕ�jS`7RM$�/�hp�t�N�+���&�h���ŦzZ0G�.�YM�S�Z�4���̰��)�5D�^p]Q�^�C�c�����q���l�/g�h����*����3��W�D�=�Is����#cx���A�.줬홱��1	�}:l:��#�X�]g�B�q4�ܧ���g��ro>�烗��d:����rpЇ������P4x,�v�ɍ�|h]a{,`��<=O�c�K�u#��#n��"�/��KH�B
.K�8�D:�֨V%�� �	�\��S����w~���@��(�i)Q�؈o�=b�*���A:���8W|V� i�}�hye��Sk0�5��k<���n�F��tkf��*���C�``U� ȕ)�����n`;�|~��[��E���8$���ЩX�<1��Q'vܐBf�!��B�ܹ5�_���w��찑�jn�6��둶��fV�������+2���`V�X���i<Âי��J��@n���z�S�_#���G�h2��)~_ʖ��,��5/�U:��X��9"�-n�^P�Q���I�Etx}���f�Pd<3�.��i��I���5W��״/0^6fj��2/5;_���#"�{ʥ��OX]���* s\+�7�3�ܹ��6��؛3�Z��զ.�4E�,H�vQ΋���0 ~d[=Ʈ8�'����8������䎨0:a��8
�Δջ
�/I����lÃ����ظŽ�|���߿��,-Wճ{�o�ȍ65����:v c�=w&G�6���Ԭ�i5k�t�z>�4?;�-��㏩90��UޥWջ|<���=����{� �]��EljS٦IaH+[��Da�bW.i*l9ܧ[�Q��)�S9�(�R���z4M��_TR�ws�\Qn�ܜ�O�J`e�
i�:��;.��:ԶsH�ޘ:PU����`�F�eJ��[�xYh�ؽn��$�qXD�d5�8sn^�j�����]|d�{%ZGc�;�Q��\T�7h���P��J�����]��\<��ސ�]�[8��,-�r�v�9<-��~_�`V����;U�nvr��gm�ֿ�m��E,e���mT��R���k2"�遫��{&e)�_�������J�7v�Gڼ� P).���Z�qZZ'�:̊>Z(�O��)4�'&�.����	���̘1�Wc"�M��Df��<���DA��M�����>��������~#F9�m��c�琡���ݑ�۱/���	%�!ӳ�?��nr'�
eq�k*TVCˡ��gP�bWH�Յn�Ňf@TP`K`�9�]��N��DC���K3%<ts=�1�R~QɆfx53XF�}o�'{K�и,�����$��"����_s� x���;�����k\���BN����y�[{WL�Y���j����+�,J<";����bJ	�-�n A��9v�E�w�Q2�7�6�[�ˠ�!�٪�?�3G7�?J!pb4-e��1�s������/�y�.��#�(����JN���3qz�i1̈���9U��R�v]+��)�\�mM�J:����5�S�����)��7�����l���$Jy �t3�V�Y2�bf]��om�˞���A�r��V�SBK�-sk�s5�(�&�\�N�^��pqǞQ}G�*�iob�S�>���
4D�!�����/���b��c+��z��[{=�<��b���;2;�\�������fqYՑ�?�N�օ��"%���hkb���bQ�������4�<wEET����\)Dvd=S�,Y��>QMK�"5�c���� ��B��� k�����"Qj���^����-<�Y�!-�J�?�]Cu���۞��ѝ3qu:�$�i9*0��Kx1D�F;��~��8�9B8����ه���-:k�Y���ku�b��=�n��b��sN{�i)F�Y��K(��>��:�9v���n�x�Z׋�h���&�wsK��0�Z�p��̄a m����t��B|��C��!/���i`�i$��u]����Y!(|���#��ypJ�8��,T����L9�̉�N�-�ђ���Mlm�}΅3� \ ީY�)~5�٦�n��s#0��ݚ6)��rTiC�ɻ�~�����t�:��ӗc���&��u�;�ݓ 9�N���8N�1�Da���!Ǻ��PK�$�I'�����&��R1-�z��+��rUrݚ��P�eCV��G��|-�aڈW0yC��539Ą~�b;�)��]:j~�\�!��p!��G���v,�8��iF��|���2��(�n��*я�n���9Z���\��㥞��� a ��s�0�8Z@�2"1������H�P��W����a��X�v.�ΦEW���)�P#���
FT�'�fdo8.���^1��)B4�;�.���H;mɈ���Ny݁q���A5�?�eh���dC�qC�B�NӣS�Qm���M�Z�l������n%���B�!��M!%���x&|��=���`?lfi΋�����L��/�R��2`$k!�2�a��2�Ht��O�S�B�/~�Ak�����s_:���M��b��6�c�D�x���햲�Qڽ�$.^ߤ!��Ip��p�JBrR}�(�HL���D���""�pX]��h���G��ϔ�[q�����h�&��
���8�؍� :�(u�5����bZ�������CV�l�q����f_���Ȁi����Ce6y�l�;�!M�խ����a���[s�cW�;�w�	��6������㴘}�����q��)�ʯ����Ƿ6�]hP�� �4�_5 �W����H(EC���p-L�J���*�"��x��a]��d+��}x�8��X��yKΟe�$���P��n�!� ���ͲwN �d�s@������?��oo"�FU�U�M]�T�ߕ�U��0�^8K���al�-~*��Q�!�������X/����R���@NH��m�?��˼04��^�#	74��B��?��x�X>d��V�L��.VgO�]Aܞ��\uCk�0���:�4�:��S�,(w�b�_���\qv��$\��P=O��u���.�T�`��e��u��vA pY�,��#ǀ��'�O�x��-���:^�>�����/P�����L����W�����vdB�Ϛ�"�\��0���rA�B"���'x�J�p ����H������������(T)ʿ��m�ta@�i>������	�zN����%����rܽk�u��L�&��J0h�#{y	��\�e��M��WF�δzRA����t%K*�Pv�#�.LB�%�3]��6�|�L�hZ�_��D�a�I'�d4�r�;��te��b��� ZF��2��7���D�/�Tn:��H�dQKz��t�0���钄g����ldR����WG2����"��;o-��-�7TpU>��MT�ao�{�ɭ�o��yg�����k*ݰT]F�J4(6��&l�phzm���i��W��yA&LN��$���#�fY���,���a6�z�c�f��V���W�ý<7���Ϯ�L[��p�|����Q�H�~�t͟���цA�-�|<~��]��B��B��齞 *t?j[�4��S�3������&� }ģ@�A�5��î���T��{�j�!ThN�Q�1�Cg6�I������al���m��ˑ��x�\=/f�4�(:���۪(l
o��
�;S]�E-�A��×��al��ٞ�>��bVD*��t��S�HI:vg_\��ux+b�c��>�P�J�d�����=x�y�����X��Y�����7�(�t��!�q�H}6��>S|g.}[���h(�~��TBI����cT�a"t,��6T���ߝ�Y�+>c��G"�v�0��6��h�*Xފ�9���_��%�%5\(�wB��ח�]�uY��^�#��G�ĺ�w(��hϭga&7�gOk־\U��(�!P�q֚ �L�BMa�~rQ�͌� 	4N���~*�dhP�U��׹FO��;z�t�^�mYPG�Y��nh���iQ[GA�%I�N��u.3))67���,�U?D�-u��6�)��M�d�E�t����'�:$�Hi�yk���PBB/ݐ������?���L �KSz-�$L�0,F�t;��k�����T�թ�\���VmD��<�>��^�_����g�)����	��DR11�,�p��E��9�7h3M�A��=��wlZXX���k�}3����7��٩�:M�|�Wrz�7�<��� �2�/<4��E��S�0�T�~�&80�>'i����TL^���������.�f��=7�?�����bs[C�}T�}�J\���)����M����R�Qi�O2y_Л�j�!�U
��)�jk�C�*К#yw<A���\g����5Y��\\�1��:@���q�ג�h�g��C��b�\��0��{�b/�;�z]�iX��2׌7G-������@�o�;_Rx�-y=��mB����>ϒ�������b㉑����q+b z~�Ca�/�:a�*7`�S�D��gjfq�D� Nr������QJiR����D��%�p��V��0��ەu��7C>�L�3_p	#ar!�%�F�1���C[�0�3}`7Մ������{FMD�����9�u���G|T�â�࿦��J)d��m�r�IkvUN�[�n9��&'!8.f^�+�`�&���V*�!�˓E��Fk�6���~Đ(�Ln]��!}���ǔmC(4��inLJ�h��n6|�o��,��H��"f���:�vC��^_{@��č�n(�t���[H4 lƒcU7�+�r��7z���WW����P�x��@�p"p��^� �A@��:	���6A�y���zm>�lP_�V��w;�u�d�c�>>�Zf���x("���JG���|��d��LJ[��\�'�
Qw�(٤��4 ���D�J"�
��>�+���2��m-�]���$6	�e21c����敀�%/��"��:�@I���u���6O�,�+O=
�QZK�UaD��e��%��rv,J���_��/,�|B�c��zb4�>I(�~$��Mi��G�}{�O��1�?(�C�ρ9!��@��"�]3I,�� �W��(�JQ�k/|F�z҄ 6 ��l I<���ߥ�zp��߇H��RD�	o�fY�E����/�пQI���Δ-d��_��k"Ms��+80@�h�SX�k�B!�.pP�ecs��
l?�:�W���yǙϯz[+�?�˳j2�\G��,�h�5FU�rO��a5�>���ؿ��4��=%Ԁ�n)oT��M��ф*W������<0�=���;�[?��O�+2�
.��}�t�)1 �b+d�h1�����cB��V�g��#T/��"�[��{��՞�.i���}��i���w]VԌ/��&a�������¹����Ɇ̇����ŝ/�=B¾��l��c[M�'D!��{�ʹ��t�F��T��Ga�Rc�{�q�bv��kbA�$t"tM�uFC�)]�]ufD�h�蛏��
d�a�̉�( WGJ c"h�7�$�gL�w�W�J�3I�O�B�š>�	ղg�Z'�(��.�6�HA:��4��\��MfDl�K�@a��C&���	���L��[��*�u���к�an���T�;�u�|�[G]lH�@��ia���^	�6�T�h��@�����r��Ӫ����W	BfF;Y� �����+��QrIR�3T��>�ړ�q��X�����RS���jP���,j)>��"N]�C�ecR.]���l!o۱�
�1f�C�LZ��f�DQ�4Q��,�H�L���
��93?,�V]�N�ׅۈ�媸�Gh�gb�����=�����~�� ��Ȳ+�ܯp�
X��b���EA�к��,S"�a�^}`~�����i��۴H�i�[�1�n���T�Hs<-��	оt-ka��V�O�V��Cl��'r���A�d��<�����G�jd���bo�x78=}����P�Pj�gݩFB1�5=�E�,�όK�8R�#�FoTv�4c��J�\hJ���,�㡶�)Aht�\k*������]ac�c�Ca�x����.�z���Q�pr�1S�l��@���?�O��Hk#.\�,��<7	m�@iw�vú�.Y7q>7�R �|89�mBV8���w`	������iTXx�\	�ˈU|#��@��9@�xΟO��\���7M�HaU|��o���o)�%Z/z�a�q��Ț�����dZ���O���NP�s�vNF=/�k���VԔ�rrl�8]0h�a����b��h���̟R�)s�^slL���W�_�*y�ac�C�+F�m�]��=��[�R0�/″�*��]K�;��|2�,�[�D(Dƈ�_�+��.�]�>tB�q8ہ�a����Į:Im�B�A��#����(�?����(�i3nj�{�Mj}�U��t�
�Q1�m��(G�^<����D�ꆖn��p�5αL����&ĮL���T��֛"�QI���$��/̙R'0���VP�oc�,��Rm���ď��hH2!���vM��諆�%���I����U7���KV��d�.5%�!J��2��J��^ڝ4��iXW(�� �AՕ;N����$'�r�����~�"/-9�u�m�|��-����4M���b�۬�MPG�H����QV�����W�X�D8�Y��"����enT2��|)f���y�t�V��_�9�v�:
�찡�v��\Y�L�F
��/04s&��K;�����>%bc�$��?�l�Xݞ�%� �Qg��d%�k��S�igp��)�YC�5�g�M���2�_��x���^�P�b���A�)5+�f UEF�}�aSޙ.u5�tB��P��p�A�3w-�#� k[�5	�u�ZD0]����cz��Y�4���͐�����̹C�1�����{Ox��"�@��B�Ie𦘻w�.�> �D?�ʥ��;CU�F�Y�逐g B<�
�H�w��|S@�!��c����
I�RA�\,_خU�̂6v��Q/�0ZdU�/�S��)tU�^d�6�>�>v�S��f7fhz��C�L<B�{�bѣ���s]:�1�z�!�z�� L]=58�zkq �Gu�����R�d���'��槩l�1j�o���
q�H��+^"���h��9/ft�;�p�n�}���dl��7(��4C��Ȕg��/|��Aq����3�o�3ǡ���Sn�j��t�&4�_��)$�5��O���1����9��$
����1�<��ku϶ͣ�SyVΦ�
K�c�5�'���a�_P���4d]�n������}�>]A437guM&��əD|-�뫭pѻQq�.��n^�	�&�P��}�Gme)Y����X9�_1[���F�H����>q�C�&�1�\�]8.Vt�o���$ �n�����O�w�\�	'�X�����,��}�g������oh0�B���H�k�Q�&�Y���c�	24-u@2�HU�`�3LY=����_e���(f�
>�z�]PT��'�����R%���_����6�r=8h�N#̦5;#ev���CI���d���Ƚ=<��������v�Xub ��zU�����x�������^ś@ݫ69k�>��Tlm=�~j6�/���&����3b�;�bM/ā+�p;��9`R�Lwh�(l��C��|�R�B���&0�͊�FFn]#a��+InZ���+�	�U����7$Z�lf��T&����[5�P�|�ͩ�g?�(�W��X��GŚ
�}w�J���\˜An����l��앒�Q�^�;��O�e`P����7�q	�rw�$]2�C�Jٍ��,yYd�?���R+�JuC����.8�U!���p �%_���+�ƛ�(�sp����4��C̵u{��l	�IG��J$�Ab 9��	�s����?���W��ue����n��.�D��H�!���x�V�?�u��2Gq>K��\)�Y�<�7�k�(�<��k��[Ew����U_�a���͕�@��{�]�3Ex��-�r�c�o�y��#*u�B`i���v��K�X'9+K" {�}_��X���*� ����&�����v_A�U�zc\��6�p��5��;g���.{�
Q�g����מZLRO�/H�kܸt$���m�#T�3������P�=C�4G��k_��_�)����j�T����p4�����Vo�S�'�%D&�� ��f��sT�S�/o?N�ǇD��&� �n�x�ȝ{��nm�@E�d�x���<j��iQ�������S��+�)}�ڽ��<���܎�Z��ts�����Mn�*���鵌��gʊ��t67�̏�ʀԇ.���Ie%T*P�QJ�
���!���Tݣї	Q�3T��zO�
F3���zZ)���]_t������HbQ�{N^l��r2z�s��=�&� ���ڱ�b���`�i��Z"��7]Lޔ3_f�-�xM�s��nG���/���417�}Cj`"��S��]��
�t���owkR}��Ƃ���y/���'���$׻���#JQ�/��Su�\r��K�����+Qa��������nL�����Fh��MF`�m�<�>�3�����k6�z�����ʣt��z��4�I�y������ڗq�5��y�v��W�w�f9����[����ay�|�gj���%���&X�@y����L^�RshJ-]@{Ǵ����/n.��?{��t2�'9��Z��a����V�;I�e���WZw������53A1'���F�:|�i��38��~�n�w�R!�x�vz���(*�#�����<��e�c���T�;�x`��K�τ�F5�O'�+pS�P�R��%ݹ����Q��bp�d�}˜^�nj�36�43�F�u�`YҐ�&�3q�w�[���?X��fk)ii�Q�(�D}<�(�9�,�E�rj�����gKf. �o+������
z�{�4Y�0�����nR�P0�C�M4vtv?+�W�:�v�*a����AK�.C1�dŲ'��T׼����i����^/R���:�\꣮������a���-J�	1zY׹S^��ȁ��o���V����O���H]�KX�1�fRc���l�:l���>1$��VO��'��#�T��E�1aRwr����D��MQT��7�16�3�S����ֲ�������4�7׾��m=�\���rh��y��L�
��&�x�"͡��E`���!����r���g��t�(�[��Be4��_�̞؎����,a^՛�a��y)�s�(� w��4�a��$������<�D �n�s��W��/7��6^V��������C	��(��5�|��n�J� �đN`�0S�e+#~��/׻L�G�%C?��iw�T�y��Qo_ԁܘ��m�ڗJ�̟��U�����1kD2@a��@�9-�2K�`�K6�@���}\[��n�e!g�J�a��v�� 7��=��q�NmQ��_]6��\[!(���5ߗ��.�Q�k#�����5�O܅�"���
\,(�(vx�<;k�����Ũ�x1P�w~�'l�AF�n�-Hnse8�y8��B�!͙/����OŵJ3y�6EЗW	�.m���2Ӑ�I�%��8�꬐�g�w����ퟦ��l;�;����5혓U�cM_��މP�������)�A��(�r��qCj���n�Lԭ�^��d����C�/!��
�خN�m�R�GHv��d����pt4w��o�T�z1�������Y���@$V��)�
�sS���M�6B�ҏWZU"K��/`���BC���߈�n5A�*��a��aď�ONڣ���!{�β3��
D�TG]R-�|�
`k�,�s���k9/���͸��_e�+~`�zy�j�c
�>u��S�̑|7Pn����;�Z�6h�j��=�Q.�M���c���/�5���aw��Z�]��k�}g�0�����M�ϱr��u��\u���M�S�kқ��5t�OS��0}�|�!R3B�n��)��;��L��HS8�C���H�Y�a��8譽9��^����W�4ޯ�R���|PqVn�\��M,��~��%2�����R!��.*d� �P�K�	ZJ��6-~�$����cl���������9�!�3�t�.8
TI�� +_R-Tf��E�jq'�~�P�.s���{�>�'g�]����Vpk�}:��2�$Cp�Td�%�%�ùfb[5{	�?��<H��h2�d��4���C���+�W�(��Q� L�`�m�����g��d��7"��@�p
[�����$�}}Z�o؆��('��\�	������0f�]8���R�ن���D��Ǐ#BP"/N@�=+jPe���{�ȓ �3����?ZP���m�J�a�n��|�gO��������o��n#H�52�S�~>�l��Zȋ���6�~;^��-t�w���ߎ��=�R6dqU�])���"f���F���	�������H��t��z�155u�V
9D��}���y-γ�H��U��#�x�q�i���o�V�ƥ$q]4��N��2R+�t"�~�4Ah3�V_x�~z?&(���3��Iu�VV�>���'�2/ ���!��A?�b֜5�E�̦95�ϐ�o���Q�b\~Q�>����>cyoH��݀��-�A��ꖁ*���z_tu�_��'��>��9��"�ֺ`��)oa���sl 	�sA�0|\��!�\`Nd��:�,}Q$��h�a�V�/�$��/S	w^~��+SK�<Z�]9)T�#s��]�3�K�fS��1�d�m�&	Z�L�iÂv�x�\�=�X���O������c	�:r��ݬtSwuN��0N1�Av@qWP|��j���	v,&�O�.ɵzԐ6A��b�b����6�CI��%�=��f���)��<��?!�����a�Zr�,���t쇋\J��6O��ޗ�x���s!���D"2L�Rl�)�����U��d��.���/nM��Ť-o��������Y�T��v0�>�$8�`w[��	����5ϋ�n�F��T}�x�}�P3x��:��f:P��|2�>_a2)^Y�q��utc?���'�{aOr)l�c�䆴f���: �,?�֤9�[����� �L�y�r����w5������ �Zg�N�k�b��/��뮼�A&��QT�;��U���]��o����HP�$;pu'��F� �a��ժ�"릅�}��'`�/>��LN��;��[��2D�5�]�e�[�`j����gtG��\�u �OkYϬ�Tey���؀��*�x����S��a9\��S��m�L1�^,����O�2��Ī 6����5�a!C�y��Gb����]���vb`j��	KMH�}�*��{򸞹i#ʖ8�a �df�a� 1��Φ�t�5u!������*c �JVa�ސS�پ8��Y���{�a�1})f�&����O=�b� �[�����5Fmf��.<���O�&dv���c��nv��8�׏'ZKF��2�Ֆ��6!��݃����g/4��JF��1�4Y��_p�������o�$ǩn?�s�x�y
��H�ݣ����p9�a�?���2��4����j��F�
����j7AF����������-<W9>��|���� Κ.�'�6��0�s:�g�}:=�}!��kH�|�v�B�a��~�5O��3ܔh6�l��Mw/�C�(���p�s�9��j��G�YJ�כ+��JE�$�[-�T\.��_v�UUC�$���I�B�*lK��Y�k�������_�x��:�}L����P���6g9�"�=b�R{�H�/Z{�
hA�p�F(Ni����'6�z�\���	B�2{E|�b�]t@�h���
Ri��T:KǗ� M��r2�uN�b��Hv�����%��+":٧����(W�aݱ�������y��{��|�{�x/��KWYa�q���E������Ӣ!�˘OG&���V�z�̥�`�)V$�y�D�E�y�"E��*Z��5��jv��S�FmG��Z�پ�DO�5FNl��v�)��~=�����! R��W�IG�p%�y_'7""-@+�OmD�2	C@�J�"�萁��aF��1a;��h>2V��˙>�Ipk&�x�ۉ��4 �A��.,`2�;u��X�������X�av�ݱDNW��܂��	Oɾ�/��՘���Hr`�%}��ȯTn��:�l���h)e_���{��fĊ�*�Hb�p��aY���S5��T�Ҩ,Ӓ�^�����ƚB)CVt"��/>n�>v��O�cE᪚4��A	���N�5�s��%P��D�Q_�\�E�M#d���4Ce9��v��*V�$;�I�sFY�D8��<N���"�Ti�o[��}���/�S�}˃sЙ��7y-.lo��:��������R� UX����1|�Cq�;��V�1F��"o�rk)1Z�&�=�j]���p
i,��"�\�.os/�ކiK�
�T6'��53WX�}!Lmm�xP��}��X{�`���6�0˓W�9,�,�����׊�q���?��֢� 5���]�=��K��,~gͨ����'ɱ��G��s��kP�c�A� P��	)'\�����@Fl��]�hj}�)D(d�*X��a8��M;o����n���d3!K1�?���|rӘeJ����ZK��,�i�J058�M�N���{:𛙒In�Y�,������|V�8'h��)�n�A��-�r�}�}ؖjNҳ��yw4m��5r�հbD2��p��u���`Et�y���:��SWb(�Qz�T(�����(���ğ'U8gJT��7��)ͼ����d�ӈN~���2�azA�w�`�
����D�=|[n�\������^�{w���<��rڙ�TXk>�e�L��yeL-��O��T�&8y�h���J��n�Y��*����x���.��1�Yޤ�hO�z�5s��w(�F�Ⰶ��M%�=��P9�
��lrw�K����_4˛�4�5|=�\���*..]��K�Ϯ����X>���<��US�2'�fɌ�Xq?o�(��
΅����H��8��&��԰G_��]�yoчa EDc�
^���5���E�e����#�O��ǒ���2�D�*ڥ��q.K���R�ANC��=��$��2���1�:>rh��&�U��}F���'s�ʦ�ڶ����öc�]�ϟ�Nk�����<f���ֽ	[�p��SIQ9����O3�����~qg?����߉r��:�:�f0�P��1 �-��~������ńֵ'��P5`b�1����j�x~����^�u�_�-j·Q��x�0�|��[lp�t���C�f܍���eɚ����B�ed�"��(ߗ=Z )u��+Z��.�44�J/�h��F�h�� 36���欰�?����̟����(O4VU���I�'D��� ^d`�<��|�����.<�Ǻ菎�F֪m�"�H�tn�מa���\��oڞ^"����	Y@0x�Qn�Kboԧ1$���'[�D�to��,�)s�%>]��͏��oL���l�W �`��}+��#1E�j�"�rMJ��e� ��A��<��uYUào�Sd�)9�#�C���"YD�P�xC���Q a��Mr�}u�j�� 0D��[Z���v�ii`�� }�������cpsQRlc�Ȓ�DR,�7�e���P[��j�P��u&P��q�޳1���]��X����]�*G��n��������Ox�-=��K�em�Y֌<��)}s������Le�0�[W�;����Էĥ����Z�u�"^2����� ;���!p�	�l��q�Úϵ'�)L'�TE��g���J�A�Mӱ���Gw���RĠ��9�o����	��tZ������E�D+x�x��bx��\GfC��>Ӝk�s�9�JW���c�^pq(���zN,��/v��|j��WU�D�?Y:W"Ӥ�s�i�O*�Tv��{�0�B�h48Wm�{<B<�g8>#�V}�W#8�LZ��*"B��d���9���m���?�Ma��?Q?�g��M�V��~�0���k��]#�w�-d�^
��^��4C{*�\�˭��T�=�<���O���)73۵�8���p>�Hz��Ȅ���w� �'���r���
F��w���V�!Qwt)%-���*D<�V�e��1!����/��X[b�A���c�
�q��#�5qw���tZ�^$@<��T{`�fw�m<������0�x�֧��(��H�}�a��W6H讖�y7��ISn��<��'�)��J]�jTa���K�0�̼tZ�;��:4EC]�5~���ͅ%��Da6i��p�mE�' �j��*�j�[n�2�a��mC��r�#{��6��ָ+pGe~w�/z�"�׬x� �
fsD��i���t�z.\���e5"��V�X�.fz��5�J�1BFl�ZT,���K,�X�VWȌ%ֹ�(�}l��g�R�Ĵg�FM�]�{�}WQ��:��jM�U�Lg�dj1Soh�^R�"����TD�D����{���3�侹����^��UL�:�R�j�A�-0.Ƈ�s �W��P��;D�`�P�3���%��e�'m�e���tf��P��>8�V�M:1��5à0d����e�I�:��WГ.�1��9˱�{${�~��Y�(�6�}ڥ�ڥ�ݠ�]�Q���ߤF��U����9�zu�t�b����/�t6Q��O,L_s/�gx���%�c�'0S��Q�u<��e�DS8�Ȫ��.�m��^���"��Wj��$�e������o�.,�J��/$�}*0�"�6�&ܶ1�l7��\y8F��\a�8�z�9};���J��{�iV���f�GY� lbuۜ7���j� \�XD�Dx�Z �P;�v�=���zZ��#(�6X,J^wS=�Rz-(�����~��� \9-/k�jO�)�F;�K����Z��4s* ��6=�N����W҈<U\&��s_��G-�j)����n�15�������s蘞#  ��)��Z��`� @�M��r	��j�?��G?S�,v��sK�L�\4�3wL_�D���4��C�b��T*N-�B�9q�6�B5^*�]R4�����j_�HeY��@/�h?��p���N�T>(,E`(�p6�e�����OU���"�LFV\�YoE7��t��b`�@=L/X��d�!�mQ�2�����%�I�ߨ�w�F�Հ!pW�����v�n�4�;��݅f����Ϲ���rb�j��P�@P��Y����<��P���=7Kd���z�+>4�� ��J��4��Q��W��/��w�2,��k��pZq�\c<� nͺ�ۺ��[��P�K[[��ܯ $��4b�p��ۃ�n,�fq��B`z�>l�f$�Ds�<	]�a���� �Lz�t-G��'=��l��R��i9�0U��A�.Q�Q�g�U�p ��mQI_�#�#RJ;��iPc^�
|Y۬;��^�)�8hY֬&�xf�P<� �T>CV(4�B}����[��9��B�� �� D�C����i��@��MD��#�4���f�nZ����QGi�%z�.?���j8��I�m����x|�
�Sʠ��9�\C{8 705$�ji�>T��r���݁�Q�i����4�΃@�����È�^qL8u�w���Y�M�����GOU�\���_��,���;?���6O�և���ë�λF�H�f��\@_�@��߰�<&�>v���I`�n��_ݴN����ڱ��>?s�G������V���j���<��y�~�!P�߉��Ls�� /���\hX��$'���4.�q�*�L[+4}g:���4^0G�'�.�)��~��G� [�*~`x�;�vf��_:;{��S���H�i���1mp�j,�(B�d����[Cϴ�+��
:����t�)B��"�?G�	bFle2`��T�na�1@�3���U�J��52(�" ��mA�!�� �xJɨ��+ϴ��Z�6��E/˜Y,.�(�7d���:�YI�Ъ�\�&�R�F�����w71
N(�#s@����c8l1��[���a�T��# �u�Yi���I+�B���>�7ah�e��6��0V�5�>�?ɓ䍘���Q*�ۉ��&OJ�����C֊9-�����Q�>� w�ָ�Ū'|/�N�.�D$��9���"��b��g^
��o�������x(bYdkc��{�%�Ռ"ٽ!��H�Kl�!�T��b�ಱ�0��I��}����j3�e-4<�f�p�_[+"��H�����'��Q%d����� 1�
W�{���,e�\7��r�(�Ȳ�9g���ٯ�ݱt��������R@P�(Yl�e��^�Zޭ������VH����1��&���m���N؞�v������ �Ђ��U%�g]���_}g�Qo�Gs��s��L_�Ȅ�qnZ��3X9x0�դ����nݔr�jӁ-w㬋�1g�7C���[�a�X�������ޑ/<���l��L�^�)����u�!�s%��_��7���$��l���j戢�lUf�����\.v��O�}���6kur�_��5�BTM�����B Ɵ�Q�gj�A���r�
*���j=Xh����D de�Kx����a���n$a �K�+���M^�{����j��c3Qܛi���ʾI�����Bz��f�F�o�����z�����^�:'y��:7T&�x�c�H�M�a�a�w����_P�V�곭�(���?>��-)4u�4��� �s�T0	<�A��}:���U�|��C��,��?Q�I�j�������֦"�3�q?Ʉ��1`j<�����)���ߞ��4��O�d~���"��؊�(�Hh>�E ߅t~�p	-��m�s�/q;j�X�($|U��t�>��[APs�����(�$���?���z
5M��{#)�8�</L�G���W�Ľ�0���ga1�Y���H�-��>󶭬�����~�?qjK�5M7ğ!�����9M7~-켈�F�14���a����ɔ|Ad��TӅu���ӓ�}��m�g!@
���v��
�'8\ՈZ��)y�z�Z�иG�*��u�,Ak���������@ٺC��8���?W�Kd2ʝ�͢Vپ�ʲ7�Qi�0�ĬU(�{@l�-;{c�*��~��D��>��_����@2^ѬCQ���*�и��%�� 	�������hO%��2��t�.߭�Q��Hv���b@��fNޏ�r�<=AA,B�ʖ�������9��Ū�
��?�т�Zێ��cc�T������a���a�������i��֓��fy������w^���Z�P���8�����e���f�6��
w��}]��T��Bs{�W�]��f��I*�7��aQ�UK8׋ym�Y�X���?"����6��n��;��j�g�����etX�<Vu�b�A=_AΔ[k�n�W���}�s���>�|��E֧�8��(O!-�z�h���cb����Ozy|B�tm�ɵ�s#�>�8y�n�&=�M(��������x�[�
��
w�>��AlG�H�@��G	&�#O�Bf��xRZC� ���ؠٙ=8@��Џ�'�n�v4���	�a^�y��z��rN�6h�"'X��bݰ$nGCҐ���P�Ԍ0<l�̳�����Bo��W�KIj�ɫ��/�Bիd��I�y�JY$)���6�@$��(Y(?�s�ۅh�1M��h+�QuC4�y<y	������JB#2�IZVb���3�%�՜�`V���e�R5ϵ�հ$�Z## -�2��{��;u5���8¶�.��~7&�0̷2�=�eu9���v��f�V�d�Ȭ�\��g�flF>��d�w,<�SX�HV4�qe4�=��4 žM���=�5�I%�;�nj�{���@� �8��/�{*����Z�D�}ψ��Y���c�< ����4T�.�rTu�_�&%���ͥ�l�ԁ<_?�|�H|����98w܌��)�e�<����0Z[�D�Q��a�l=,�I->�#�K�c�ƃ�0��k�8�#��u�@hۮ��������1'���/�b�\�7��T���Fna!9:4��Һc��r�7�W�֐n�"o⠷ya�H��5�)+m�L*T6)?��$���G�]ka��b��ӆd�u)�hazrW��#v�^��o��U�ل�΢3@^Ӽ��$��6s���j*��%Qid����E�����P��bP-UN�p�<�xV�;��zb9��|�z��!�k�[�M�ox~��X3.�7�$������o3�;���AhQ��/���/�q��E�`Fn��S���_*��������n��CA�ez_���ؒⓇ_�BU����X��[����7�5��'g���XwӼX0���Qe;�p�s�S�<[���d���7��Qsr�������_�� �L4����sݹ���x,��#^�����������ZWG"�~���Q	�u�w.��!��=,x���SI�F����N��A�8����Z4�$9�y9.濱D�ȋj�Ue���7�[AS�O�)��w�� �����] x����^"��i� 9�����D��cF�t]�)"�T5�/� e���n�Z�	��@�����+8I�ѹ>�R���[�$�V�J����)�x>3����6 ��A������Ŝ��l��&�L�*�\����ø��Q�=�$=�{��.��L]^#�r�����P���H��\upmHD[�iKz�9����|��T�q ܾwa��(�6z�$	�qZ�VW��,'��l$��̺P�z���HŪ�^���ޢU/َ�p������)^w����A�3�W�/�������q)bV�ԩ���r�h[�(rD �AZ�*7�o����¿��Y�k�YJa`�M��@��������S�>�f"��?y`1@L��%*��_JT b��mi;O�k��ӻ�^�=��#hw�� (L�6du��W�oo���E�
�����C��~��L'$��6zU��ךuq QϢ�d�hF!�N�IӶn��zCu�����v�R��-�a+�M A�J���䛫�_
��Tk{�T%�_1��vOdL]m��P��o�,�c�2&�2�7�� �C~z��N�FI����.�������L��a�RW�fp�����	O������IN)�CxuV�V��/��E�y�G��GbX�{�VԺ#��| ?�T���w>�Fq2�mt?�%X��x��aѰ=[}���n�i�A�7��e �T�cb������SdD�s�b�+��r���ʀr}iNχ���~���#�s����,u �0J:ǽ�z�}��,*���I�K%Φli\�i]�t�{�������m+u��d�{ ��v��&�V'w�ɉ�2 ��CX�5�>25�0A�O��/*��u��	�_Oj���w�ك��ބ�/�eK���o�s���8�gc[ɤZ�<U�Ç���"�\���S�;ׂ�L�E��a3�R�$�� ��Q	 @�Bp�ȩ(����@ݓn������A���;x�`ڔQ���.���Fw_D�Ǿe�H�����00�oe��OS��[�N��I	�E���m
0(դ-4��<d�_�0i)n[�u��/~I9&�x�����1Ķ#j�̰����z�s�8a���=�g�]j�dl:s�RkUݼ���.�\/.=����4]�O~[�PrG��~ب��z������-e鳬S���G^�=x�731JJ����ڃb0e��{�j[c�UQ�#�����G�m�{�}���Ɨx �"D�7���n����l�A{��
�[�I�D �4�f�XI(ؗ_J�iR�vNs��i�n�=Ƌ`����5�L"�!o��~�w��Z������ݓMrs8f�k�YNz#^��П�|ľ�V(g�%�L�(J*䭳5v>!bЋj��b_�b�}��ؒ��G�,�L�?�EqP��.��	ތ ���� 4`�)L��z�21�_�;?�wU����M�Z��,a����eT�X��p��5��&k9.�I0��&]�^�.s	�s	@7/�+�)P}#��C���0�|�l��.�R�@ʕ����v�VC䯅zl7�;^n�Q���4�J��M�����l^2�C�B�H�����2w�4����X.}���¡�1Aw��2�ec�
i�U� ��p�쌊�?�F{iyzR���2ʡp�0r���	V]�{.���^��Zľ˭F����]�Y7��/�g:�WQ>��^���4KBb�����:�%���i�tp��A�B0�↛��E�ze�KT(�.�^�[���nZH7����,	�ڱ��R#�Z�e�����C
"F�6��pho#�@(/0�Tj���+⪢�x�Տ����RR^�t@+͑AV�%�v_cҧآ�#v5�Jٽ�	+��U4����tj� �e�0vF�~)򂖛�1�7��4��J�c�<��	�[g�3nC`i9��3�\�!�I�$��w<.m�re��y*� ]�6�4��W�	!BCy������4�*g1K0-��H)��P�6��G7W�i��y�xAH���P��Ea,�D�5���:���U�
�c�^���]i%�_�0�0E�J�f�c��u�������2�	;Z���y˪�45wg!�U�F{���u�i���0��R^ZZ$E�)��,��@}tnF*�4z�/z�oﰎ�.j_i{kfȘ�,���N��^�]G�)"KJ�'�}s}������T	�Uјiˀ"����ᢵ�^�]��C{�t'��?x��x���� �X�T�&\�n�#g2�I�:g]G�HE}|w���F�z�t(�l���T�y�6%�moc?����U���W]t�Z�o��39b�{�>b�z2<�l�B���.j�o�q���~�&��"�� �e�I I&�T�Y�{���P�x�ꪭ#�k�2�������������Nh-�.`����ъY=�Rz�����ǋ��z��s�r���:�����ʏ�$h_`~T��4Ĳ����MPh*r fN�O����Mq�
��C���^5#����W�@��"8%-�y�]�V�]�t�I��Y�\�E`L�Sw��k�G���I�_Rַg��	��	&N�S�=��i���?vR��&9t�3��-�m9�0���7R����C& �e?`\���}�K�5�=�C[��G�%!��J)�I�Yѥ�9蛩�j�׈�k7	8<id��va��� �0l�u��֢��򔤘��p�>��)�̶�U�<0̩�l�>1��v���3������؝	�D��@]]ّ��[�Y�La��,qči����#=�;�J�Lڋ�������*� ��������o$���˫��{45B�j�M�6Y���w�j [eY^\�6�B�bK�K��hL���nF�`b����*�@ʇk�����S��B��u�,�jd*��M|�8��:'Cx�4�y��R���g�����!�8j�3])�;��/!}y�G�۷�`Ȑ&E�\x:dE��ƥ�{��o����azPç������zH&���[Y2���,x��ig> �
�s�U��AH�W�fJB(����@E&:�J����̻	k*>����Y4���8?t��<�&���$����C�
�4�����(:��b�� Wp��Oa���z��&`�% �M9iX�s0ӫ�H���L&]�U;�2Ti�u�� �����x`x)���UG���Ɓ�� m`S`���H	�Q3�C���Mm��T�1l (Ќ�9�@�
j�	P-�/
����ݧ�V����Ӡh`��LU�1�l�:����qә['oXnʢI�����-�y��9aF]t T�I1Ҝg�AV쯒�b�8lZ�<`=��d ��	�x�9LS}m�w�\1 ��)	������6p���1�N4�>���:㞑n)T�[Ҿ��@vŹu�+���@�Cah	�Jh�_)T*�@9gs����O���*�RK�-�U�s��]���YkNOG!����tdָÏD��΢��yy%����|����~e�Na��;��&MK���(�}�Y7B$%����qnGK�Ƭ���<�a��eF�Hd��fM�+�IK?��j��� .9gU��*;V��I~��$A"agU�B�\�1C6]/$FZ+^����U
�glNIR��&�.r��<�0��aq�,3����3�j��+�?+��Q��+u�{"����1��L�c��gمC��W�����*+{/���!���xrt�Υ�φ�#-t�B>��<I�:�V�U �$�V%-UvC�u�hs��'�~U׃� ,h6R�׶iPZ��1���@��� ��(�7�����X��zI�A=��xC�7�{_3�u_�`��ag�H�/T�7ǿH�� x+�OZ�n�f����*6�{�,wG؀��,-H���kc�yu�P}VRJr�(���Y W7�0:v���o�P�-��NTdh�/�f�i��.��*v7kg��dјU�tA�+�@��Y�_��ˠ$��âLc->6�a(C:��AA��}^5�:.>��E_��8:��p����u�K��w������9��L��1ԛ$F�p.�T��F&����/�x�}Aw��@Ӈŏ��;��/u������#6����<�Dfw��ʹ�-B��9��fۧ�*���o߸�2�2�8�b:j�5 �3D�)�cK;p��#[�VÜ4�jC}o���s޿�,�}_�DL�ɽՎb����gj�E~�Dδ�=�O�Y��Y�S;�k��N��U�E�vr��{!�_)����ԟ�0���H�8KfB�+�@M�WiŜ����[�^��o2~���3dj�c�p���FUvwT3Am�%<X�ɜ%����fN�:;^�>�G�D6S�P�o�Ɵ�+ )@oj�&~&���W�+XV D� {vl��G+���}��:<��\����62�����d
��
Ò���~��3x��u)����ǂv���cuG�CڮՔy����l4��(��գ�l������Z���h�ȫ;��bG�6�,4�0��-�.�O�o�d�'a�ip{D���������n�]�Q�.��]@��_�&�_tC���`,�a���b��'���1�K�r+����wN��Е��Y�>�@bmBo��%������'qbKA]Z}�ظf�B0y8��Z��F����2��A�!�c�VՇZ�b��ƷX�>`F�GI�gU�^M���Ş}��!�����[�V���MK�pj�m\��}�P�Z��u�#NQ�:g�q���/���V����x�N��&l������+�Z��{0�%�V��)���bМi���!�sj�s��_��Z�^�aD^`!: �G;���<�,`��݃�\5/Q%Vmėb�_m�P&�Zc-g�נ�"����Ip��|���O���}��Zg��_��.T��I�j���d�ⶤshedQX����K�O�d,a-M���AP�M�U�3ﶪ}��	$�"*�Җ�����g�3Ь�=�r�N�,�,L���V5pGM| �M���|�ٶN5�v�S\e�i�<J�n�Wy-OQ���56�$��W��ҝ�2�ő1q�������W	��@�%�d�5��h!ڿ-I��s�� �1^�.�5��X���Zos.�BJ�ˇ�j�6��AF��!d���4[@g�������c�|��"�P,u٨LʯI���f�������������׶8�?)F&��@XlUpt���@#�����߭���0��T;�%QYO;���rǣs��2d��(�?(i���U2S������׭�Hx����z���r�=E�������=�T��1��(X;o�5Cߑ!A��F�b��֡��Z�L���)Q�o�D�z7���R��I4G��UGV�U���s���:��D���k,�]��h�Z�K��(��Y���kI������F�_���CU���,K_����7ez�!��+cSpCh	��J�.����ihWRK������5��8M!n]�h�3+��C��Iҩ[�nZ����� 
��"�[���%XzS��8:[�?X�OYRi�g����a,���U�S*�����ni��/�����O׍m��ѝ7|1 `jM��� ��t(.�:����$��Z���IF1 �����̮�g����LәQ���
R5�e��/��(���=��aݖt��2����S�X�]m����[�A�M�`3�g��Ҝy�C�iQ(��cAM<�Xn|�3�%�� ͫ��wp�+E�/ÏA�L��~��2��[O���i��Yn�be]ۿ)������b�����QE�d�a񌻁r�Q~��]�c��x��f����=�>='KN���I*W���!<�'N�s^�F�fT��^��o~�<��rY�t��E�9�n7����ߛo�BG��ҘBL(�N��H�!!�{dmrN��6ׇ7^q��|:c��G²:��N������Z��e��Q��/Y��z֤E���rRm%.�:Y~a%�Q��W��g
����g9%ʰ�b�)����������Ҍ������o'����:K7�X�r�������;��R>���v�TS�Q|��D��5�	��7�"+�����du��'���ɬT&�+P�՝*���%�2��3l���V�Y����q_�d�'Ќ̀3�bՑx�b@C�!R��-��BB����KU�IR����3���+9ɥBd[��X�[�p����ĕIlx�TL�R��PgJX�4���n׹�˅a��Җq����+]�E��b�1+�$��`��~M����a�q�Ҽ	.�`9r1��rL ;���Lܫ�UZ�wz_в.4A)�����.	�q&�nۣ�[9fl�����jU���P<�Xp!����Z?,����/0+_%���._ӨƱ�te
a=�]�X������ʙ"��6Vz�7�M�Y��2H\+���h�j 
����A��zt�����6��{�o��Ȃg��%V�Z4'p�8�C�Lx�/	Z���0��ϱ.`����Y��l�ӮA3�[�4�:Huy8+�.y߬j	M�f$���&�dZ�;yT�Y�`Z��v؋@�M�b��p���P���?�Xp�~��S�Vr�Nv��<QmP�s�59�0f��)�=	$e����������G;s����Q�;�y(pN'~7��ˑ추#ޣ���V�R�w��lM���D0 Ͷ������� 5�N��C1�3�\��s�x�/I�ƌ�o�`�P>\�Ce�*7[p	<�FK��L�0����kν�#�֦���_f����a��`���:V�͖�i4F[�2kr=#ve���ܧr�ojv%���ȩ�'ݔv��ܚ��"�
��hu�'kߨB �W�zS���j������L�!?5݆^�E F2�L+���@E/�V�5̎��3ܓ�!�!�
U�����5��w`���P�p`����y��I�4����j�61ՖB�Y��0^V6��D��}�m-_�vs]1��x��.��V�Rz&���`x��(4���)~�@��f�Mz�1"��0�H�kw�r��H��Y1=j���kя�1m��Ǚjs4����,��ge9��	��Q��l�w67�^�u5'&9�|E�(2���RA>(�]�������w�����u���T)�+��~�Gp�3E]~�X(����V#K"Ҿ0(���e*8����m�K1c$t.����W�7iE���l�ϟH���<�A��+���%:/
Nā+�{H�a���\�-�(��Z[�]q_&� $�
��6S_��M�nU�d��%�������|�P�3���؛k,�����a��_�L�H�����pI t�����|J�`�4^;1���l.�z���6v�}��8�M�W�y�/��s:u��4Sv^ภD��x���Zc˔�6�&o���?�#����s�S�����d��Ͻ��n|�H�C��9��
H�Ni�f�7���b|XBƢ�}}�=���G{�5�1e��¢��{��!K�F�٪�J��eT�uDʢd��]{T. Nz%���	-�`+�-	����Qx���;�Ү�	�t%����`8�>�G�4<YՃN�;�deK�(P��o	�����1��؀�]���<�ܯ�p�9�]�%���s%��L�"��=�pl�ۤ��U�Zi��I��N��(��<�NX)$����������[Z���Gg2��Y����3 a�Pw#�8	��lߍY��v}N���k�5~`3Ll��b���)>1&��[m���O�Pz�A.M0f�XBo�c�o��S������2td�$Sb�G��r�]�Fy�J����^��:�nܓ��a�#D 7�&i����5�Qbªkv�&򮿤�Ar�Y�� o��t�A�Ch������+�-�n�b�ss��r)	K$���ʠH�P>�?P���
Q�,#�鶖�]�w��J!
sI�A��+"�%�G�0St~�����2G�W�>�A;F]g_���+.�DՒ=g��ys `mT�zaau`�F�dE����N���8��P�Փ�k\d���M�1����7|$��E6�:j?O��w�,����\��W4��P�EW�xk�]V�V�/�����x�V(ڐ��m�RZ����X�2�1Me��ĥk�\�*���O��9�_�/�Em>*u&�%^9�Toh�����C�QF>W�)�&�Tc�)����w��J ����׳���t��ȩS-*���/t����h�%��&ǿ�.]�ߊ�{��8���	��LGS3���]��� �m@�`7�>��i����&��u��Vl�Ll`�%�%ߞy�صR3���̎w�_�_!�yb��1	a{�2xkB<�y:���ֆ�Iyv��LU/ߐH�!�({�l��e�����'�H\`���u?�k��ȽV�����.9j�Qy`�z_�թwP,J�c�����V���u�1	�����΂!B�Ny�"���E���KW��5�OEH��yy)���u0���U����wPH��J�v/�J��v��n�e�}��z8��W�Nr/x�$���qC�{���|03������*Gd���7�a�,wV���W<N�|	R��?������7���ʂ����l��0x�"��2	Pp`#�9 FkVcRc�1��f; ��.�23Fn ���i��J�^�d��6o�c�����D�^�3����M�Gݮ7v����za�]l�c��U��	�FT�����=(
۸
qo�H.�.���>�"2;]�� ��� F]���Ƽv �����U��#:SV��
�9��O~^�6�6�K�IN��I��	=fX�G^uZ}�7�C���TU}j6~�uqU&����v��p��R��.�8J /��T��SO����{0�a����Qֵ�Ch^��V7�!G`��;�'���1�oK٬(��0�|<�S��M�	e�{|�etIjp>�/�8��N�k�ddc���i��~���b©'�8�w���z$��I���V�����'o�D8 ��v*�ٯ��A.�W��� :���9��j��B�\x��Ac�����ǐB�ݮwẘ;������=3.$���Ԇ��
�6���ol�?���}]в��Yqn��T��s?�	���q@%u�x謰���� ����+���>�?xF��+�!�\3׫{#k@wNP��v?���@��"1��+@G��a�'�=�#}�h'���/�6(bJ"�R�V(�3Ɵ�aQ���M���
�90H���Z�\�l���BiB
���_���0�$$��'�{��WR/��*;c��9I>#�b0{^���WYȌg����^|�Cτ��.������ዄ�#��|�_�R��Ҡo��F,�qL���AC\`7�%��k��o��e��]��Q{E&(]�߶����4��@�uS�)�$c��b�0h��r����3���E�Q�G4��w�l�$�>���� �л5�a��$?�Zj�P#��kVj���
���N�k=$�:g���U&r����9y{G[vM@L�y�����4���PC)�%&+ܼ�Ҙ����YF��?!Z��!:h[_�kLF�#�C����6�/���ßp.�`�T.����K�a�`gӁR�+&��-�@l��)���#��OF��	��=IDy�]����^"3Z$q�Z�q�a���W�)	�$���u�02H �Eǿ�����k�������Uw��;C�D����|k��_~H�CG�G�"[q�ьr��-3]��=�4�#�eM9���'C/cE��\h�~f�ONu�3Ϟ�/_4��
ѷ���Vԁ'2Z=BQe1�<���db���n4[ ����*��3ϧ����_�7>]���F��gO���=�:���`[�;)�r�&�S�:���o8�u]���o�M���M�.�B��R�[}H��-ԔE� �&��9�w�
Ē�z�m%�����ګ`kN�o�*��������PN����ża�v9qOj>