��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��˲�|U�eu2���P�1����J�2�@y=܆��X�n��t���+-1#Հ�B�H�b�~"�{����;GH��Y9�QR��c��ׯ�b�i�j��Ñ"(Y y�AG��) lW;#��2��rn n�c��n����dӻ��4q���狙e};�e�h����ήr���[�̉���Y~
�-�ʙ�d`�d�Y��8���N����j�B��M��tI na��#B�`��f�v����+�~X�<�V���~�����p��ӕ�i�:[�<!n$
�� �_���zE�0
�O�9/,rFw��)'9� �Ԟ|[�w�C��6�Ui��g���
��]6Y��uV
��u0�cπ���7��"�[/�`�ڃ��xQ�HPEIڸv������F*�Y��u�L���/�+m������R�y��E�0�k��^V��0>>G�2ʸ�S��K��h˽�<7�D�}B�r���sDf�O{���~oQ����� �}�X=�(c�!@T6�ҰH�rQI��r��`���9��e�j$T	]4��<�� y�-p~�l ��ʳ������`�����-��|`��D��h)f9�K��τɺ��[h�������kκ?gU����UV8\�i��a,�':��sJSG���*�����2a��ƶ�{�wǖ�K1���E��x=� �c��U�,�/l�4@mL�q�x�tʤ��kv��vo n�m"��fX1��5�|������ˎhkG�t���.��wg�%��Q��(�������s:���S,h��Β�p��rt�����E�e�[��,�0����֏�|�þd�P-�^��3&RƯ���:�]���GA ����s��Q�'���g8א:�4�u��Py�˃�e���Q�Y�.�.S�b�k�]�C�-�5����T��|ɐУ5e��5c8���г2�o!��cn�H��XM����"�%��d1�daѬ(�"̊f������7��	�>Z��������VE�Q�!��3�Vs&�SR�lXk;�Z"@ti��2�������b�|���!_�z�M2�QY	v*����y��J��/:���Lw�rl�cI]�-������4���6�]�n9����Dfd��<�1�j�)@�u�4�+G3�ڦ_� ��A���:\Ԧ�vϳ��Q�2��)j�U�1ŔG#��Ri��$�������1v�Dʿ��뢞�-W�
k��#��9��g2U��'�V}ߨ��݄�{�q��;�1�Ax5׊4��j���aE�zF�xd�-�&\��~4����T�����;�ًt���jrY�f���Pz���~�Bw0	>E_B?y8�E@�:�80H�h�Ң��:��p���%�������0�OO4)/r0y��3w��0q#����p�\�͒�ˀ�ѿ�w�И���C;6Vx��h��b�L�O��B�Y-�t?�c��̼�z���������w��=�fF�ٌI�Ã��@D-2������LE �h�^pmN�K��A�X~"�&7����GF����Z�����i.f�j<�\� %��k[��t/:��9��"�1���<3PԸL1jf(5���0AIN[P{Rct��A.E>يK�h�w�T�Xzd��
o�AZ��O�[+s�@�٫����܋��p;( ̊f~�|K��O�㉾jb��Z���^[��f��S�p� ,�� �4��;�@0Wmп�(=ঔK��(��3��J�E��A��%��-��~Rˍ�� 7�V�'��^�n��Ӥ5r1G�tw[Y�5t2J���:���T���o���2���Dy���T�K����*�*����@�oҐ� �6msz�0H�/kSɈV���䒮�O[�a�-�����؁ϋ*퇛�	����9&|��Kf�ȡ��j�H��iQ�U���`�}i
��Y�i>�S�0�	�Ga,�P�pT�$	!�/מ�����-����R8�&��{�&~
KvZ�E�1N��"7rl@Fe!XC�}����Q���A�z�;E!`=�E�|������z��g3��*��2��=���g*�q�huAóT�r��Ju˘���Op��ǰ��(��Q.i�z���4�*Εa��1YI)ʃB|���Q�x�Ƙ6�R�b��=�.�}D�5��J�gi�B�7�u�ܛT����5}��7\�\�\d�M��y��Xm b��F�2+���Cښ�I�Hˏе���m�������:���i��N^��9���@��¦�F��|�L.�I������?R�e i{��B��#v���w�y��O��B�jwQ�x=��x�y�cz�k��g�H&D�~���RoZ��X�g-���0�rN�6ЁC_�рt:�Z�7�\��^�Ƭʀi |_��#N�$;���z���[����HN�췪���-gj��9xLjK�����B��$���Ɂ��%P�xղ�0�^F@�� >m��v�:�ר#_�����g�@��O�kZs@:�RW[E���U���q|�:Lz�J�(�V����?�o$/�[��`��DS֪ny�%�@��[�o!|
<0�+PB�(,��d��u,h���{k�m�|��0�B��B�-_@�Y�}�A:�Y�E0�x���� �')�t3�	��͡�8�Ӛ��_6�0��X#�O��qi�G�(,P�<&r���A@��TX�s2���pl�D��7��<!QT2���a��ם�k5�-�+3�����_K褼F ,�@��
 5³���m{2$3H�k�B�ŷ�t�L�k&�`���8y��珒�0�ˈ�5�%͗Չ��y0��߁��<L�bw
�Op��s!m���h�
�MF�����9��<���y�5M��t��KC�ZdԜ6ݚ�
Ҫ���=#�J�0��wN f��6q�ה흉/�o�q��p� _M��ݤ.cQ�A7���� x\��OFk��D�5G=���Ldc\;�����ŋ�R�~�)&�el��)`����+	@^���)<|���,���$K��C#$[�Lѳ��\973K3x�30}t����<G����o�26��tR�T��6�X܉n�6\X�8e{3Gژ��%�
n}�9bAf5�h��>��>C!-��B�����3M�]�:q�f��`��4��;2݀p4���q Xu���N�u������5�,Q���(���Q��[pe�}BRz~v�]쓀Fs�9O{��C�1�00|K��s�͋�d~��Z�|�{H�,]�S��c��ߟ�JU�P�XDSߜ�d,����K(O����)�O����._�i�u��;Q�k5[��3�����n˹�'��]Ւl�*���A=��܆�o�!t�z�j�P�K�*�u1����<n�t\ᝁ_��zʗ婯�����{d�w����7����Ӈ}"�(��j!�N�'���ӴTF���H{J�g8�v�?��IΏ���e�0̇Zph9|����=Q+��Y6)��!ot��ڔ͑~5I�P!u���5����-���*>�;QY�����x��1c��T#N^��\��Bz<�|ē2�.뗖��ë,�R��Mӎ�^+2iSb"x�M*	��c����d���.��'k��,!��x�%b�2�|P�eZ)�/������E*N�!��>�W3;!l@;�֬��=�n��T��t�®�@�[�h�uE��x(@�-
��H'Ӌ�}�����t�XӒ��a�O��@s.��!��wbi��BM��s4d�^�CgfVj�4W�;� '&��u���U��P��*��ZjI*%Zs��E,a+[���-H�%3`�B4����Na�F�5Az���-v�%�1Q���ӥ�}��Ae���˦��%�$���Ya��ƿOm7�y�/Z�e���;��(r�4��,���,)Ѵ���9�n�KU���?���_�ԗI5Q����7f������~%'bފ�E
;F��Zo<:+�����^L�G���"��,Y�֑SӉ ���>�pG�.���6��cR�NB���-�ˤ}ܕ8���+�S����ꈌ�:u[���0'��٤����Ü��CiM��T�$1C�[�*������pr��뻄�"���v�𒦾C��w�����P4ʣ�2H�m�洭�&���f\O����{[��OF�`�i�����1�Ͼ�+̖{A�#���0�1�?�!ͣG��מc���z;���NÕ":�g{��Z$��R0|v� �S�MR;��uX13����sϦ������;jN&���f��=��iI	T%yg�P�d�	%��e�Vh��=�p������=0��z��mSN�Ǫ��Y��s��M-]� ���lk�g"ڣ8b�}-;j�:YU����-dp?	"�����ʊ3�F����roU�3��H��t��H�\=�O���sX�<O��C�OlJ������q%{H7��rM�+�P.nɛ��� ��{�y��tĎ����Z~�6qu��Ø 1$��`��� D��A'S��zɗ�`զ�P�ڙy�(�yaEIm�x�3p��։��f�3�c����H��
�f�Gx�mAD�7}�I��?JjҲRWW�Ɣ�Թmh�u�g��G�x��%��
�c����Rq�V'nW2�K}���h�G��+$��3��M��~�b�Nf��Դ��@pt�m3X<o�=|��� �U�N�jda�ٹ�u�DW熴��XԮt���#��|\e�R�����w�G)��PY[�8���v�3��!J�`�X���"N�j����4�mv��^u*��^*��8�t&��r��V��[]���Kk����&�pR�~$$�������e�y�׹u�o� ���/+2%D:�f�O4~�:_���k����
 �w:c`7��7�>�6���!������t�S��JlH`��	�����*��b�M��Q�ۿq����?�0�Am��:�B�����F}]hY_(�P��SLY��5�=���D/�FrS|�4�15������olhS]K�zv=�ZU�78�y���1p$�"v�����^0�9��R<i���Z~`��K���U�A9�� �'�F_:���d(��P�~�����%h�_�X�+�gh8���ƍ�|R��_{��F 9�A���7���2n<꠬��u�?��=�X/'<� -��V'�h�����w��l�0�Y��FD"�����M�*K{�y�Џ,�9J�{�ʍ"G�&Cl�r�l����BC��9����6�s�b6�d'Ի@�p|��|���)LcZ��n;�����$���`��!�>Yu�Ӗ��
B����1�J�K�zIG�|�ﷴ�*xQ�gr[r�'��~B��=�K�!��ED�f{��#yv���t
�}50А��"���͸킮y��K_/����y���-�F�����+ļC���/&=q_8h���ڗ���Z�T���b��}���j������=��2$a:���[�W��+K��-��|oV�����F;06O���f��n�x.��A�8�vJ�Օ
�M��DA"���#B�*g�<�6����/���<�)��-��<R{v�ȱ<�:�iP�v�fʄ0��P bE"@�0GJ�Ee�h�F������-�wwQ~�m��f�^9��wsR/���oo=��4xwd��2�!��'��1���`���]<@#g %����p˰+���aA�J��+��!�pi �FA�(���B����tL��'�҉JIM�q�%�N���"Ȩ����}?��R��Ř�>���ɌR(�����&a��48�]X�5c-�m�A�
e���%}jQY�p�8�fH�
��D��GZ�X#>U�j��}�m�P�..���nCy�P��<��@~e�DN�,2� � ��;߃���S�p]�.��<�,̝@��L�Y����=D��m֛�T�����x�Z���~mQ޳����Ͻc���%�rAHQD�OQJ���3�6���G`��ɡ�9@���ߔ�>s"�"M���.D��mRC���c����+&^����[�E�(��W�d���_�S����HH7g�k�i%'��_�V�P� ��WLΣ���1O����J�"us�F�b����X�ڙ�>���D�~����������UvNۂ;5Qx�Np�9w��'Wh�
�q�͗�����T�{r���~�đ�����M�HH��M�Vz��+Ơ	�˚��h'��fs�5��F���K!L ��i~�� 0	5�(9q���3�x������I+� >��'4�7r�^O}A�ǫs]�(��U��{f�g��a�mBI��eG��R0 �	���.����gѰ�i�˄O����뢾- �|x���2EC��!m�jl�+RA8H�8����Ifw�qP%�t�ە>BI{~QB��K��Ud�#��P�� ��uIM~P���
��4�����Y~����k�8#��)PQ��՘��˝��3u�������#����H�X����T�IP�Ot23u6�r�i��>?��i������� ���9��"S��������Ŗဃ��B�ڝD�B�"h�5M��c�^!>jwYQ����Y�f����<|�y9�f�+0s�b��E��.�P�b|!hn_
WoV�.r�w�#�z��&�p��d���$�Źԙ���z���ac�#�uv����zU`Ƀ���h�OF��>���s/87��NF/J�:��(���|�����s�o��z���w��roա#%:�G�_)��H�������~�ٯ��6�'U���@���b_�P�߃M�v����@��t�}/�vGd��7#�����;����*�',
����C~Ҧ���5����+��]]�	��ʠB�	��߱>�PP�j'����X��L��	W�%�9�\C�{�]��\C�E��_8�nJ��^�>�O�O����QF�.@D����dA�%ny&ZbX��Z�K�&.�lpc"�Z
k�;I���li^�G,J�%�\鞄��Khy҆uxE���a	�q(q	کTYY���g<|���f�`E��̧�Qf�b��=��)|�CP&z�Wi)��b��q-U��_^掂�"L�DX�ԍ}�y�� u��Q���v��������R��f�*(�A=��g��(%}V����?sX'���o�i�}�{���4m*����г�V�-��K�3kt��
�s[��H}i���5U�U��Մ����ϭ�N�S�,vP��ԕ���ޚs�h"�����>�����am]=1,EZC����Gzi��Ze{ӊ
@>ƾ�[8]fq�;�9�I<M�4Ŗ`b��ȮP���e�`%}"��gWbe�UI���hS�e����h
w_i�H�����SJ@/�S��D�@j��� �6%������.���{�hA��lf1�?q�7d[�	��Q���&jYY2Z-��\��;�fER9�F�dN��1��>v�w�-�Σ�x�v`��o���n���b!=V>j~�*yt��w4u��Z0�{	++
ma��õ�fq����*���
�r 0�������0���֧�cx�����E�����7���q�+�l������f�}���4��ǽ<f`S_��v�EHc�$:Z�j�随����Ae��|�#�CC,c���9�+�\<���CxjG��_�%�[��}/AXcu�p�e�ȶx��v}xEȮ�HݠО�2}y{:�%�Hޫ�~�Kʄ��=z,`�+��l������-�ՎQ=9:Z�5J��T"`��<o��ѧ5u1*��q4�r�	���3��������vf6� �AU%h\��;��G���ti�_�����O�
j�X-�K�g�@�ox9�N�t�s�l����jj'W-�6�{�c���� �\�D�w��Q�`�%�ի�M����o��{��N
���jd������Nq�%8ɳʊ��J�bO|�0����b>��ӹ&�[�5�M)"[Z�,�1~.L5~���Y�_�"�[R���y�4,8
x�*�(W�
eD˔cl�(��E �@�;WqELV���/� ��^?��=��)MhL��l��) C�-{�p��eY{��NQV�SV�#Q4Ifh����g��|�����p�#��̙�-��/��и���X�B�5��q���>�SF��~�FTX��~����Ê��O�+?\i��7�D˥9�h:X���~�dtj���o9��.C�7�Ih�D����>Sߴ@7�1����~�Sl���sz�P�1V$"�f"�q�͉���$����O��_5m,h�ٴ�%w�Wۙk����=�Fx�ꦨ�1��i��TKh�ç:� �֌�;+��;G�����R���ԍ�x"�0�\J�ְ��)%����V�\茋���D�E�ó�O(�U�q>X3=^����"L��f�S<P��P%��)�Vq�jt�4�2���<��`w�ý��%�k�(q�ů3gc��K20sá�sԜ=��6bS𑹟�ilH�:٫r��}q� ��3�ǪK*X��p_,�sJ�Q��Pm@T��;���&z5��_G�pup�B��=���,pk���E4�J�p�����E�=m�G�v���(r�<��I�^�5�٤?/~`_Vqw%j�{�	�U�f1������ ��S�"z�T�V�!��
�^���y�.O[舼�m�ZC@�;�z����B��FY��z��x!J�� 0�y�
��qUx�P`(��f��t:h�(R�^G�D?��{M�چ��h�J4b^x&��'�p�[&s��h��>���炰��~a�G��E� �qH�ѝ�@�W
)Ue��:
ԩ�84����mb����X�%{��*?ˁ��f3�G)A(t&E��1�S
��O̔� 3l�^���z�nqn��g�{��n�0i,`sn��V��J�6��Z_\�:�0����,��m-�����6@�7��2�gQ)�Z>c#�3�� �'���â(&@��L%�ג���X��yp\c�=��!��i
�>�l>]��ݑ�&O-w��Nr�~j��Bf��s"5�L-�:pCN=����f�4�)	3>O�3��-g����N�$�)���8=HkU%�S�j��I�����B�Ӑ/`���xw�����*?Z�{O[�ô�7�_.C�-�;r�]Y�b�kR��%�
���N,�t��tR.M�u'�����v��wn�����j�
)�q�RH�����Ѥ�;�� ��ٳ�Fbcr���ST�Wޓ	ޞ ���}�{][7�N�
n�����eS_yb.�$:`��&�ݐa� ~���m�XQ��ZP����#o�vH1����ƻ��Y��JT����ԪI����VZh�b�E��x]E l �w�I`�s�?��� O�H��������4'����<��Ǯm�C�B��ϩ�t[>��e�N�Q�=	[b�Ҵ�j$#)Q��]�iLJz"����hY[ݱ�����Ø7�ȕ�ܼ��q9y�Og
g�)Txy���p�o����W�Cϐ���{�#c�`���33'��nET��E�OP��;�v�ύIb��E���(�Y�S�z����UYD�=E��m�p��@f�5��"���N��&�`x��<{��`�*� m��u��:P�䍾���r���p��^i6
v><��1wnA�l��ꮚw���[mn�:�#`�a�y �Ry���
�����q�'b��YM$^�$p-[h�M��!���t�hN�%���'r8V�s��-���V���Leg�,��s�J��֭G�����	��вdHp�7 ��g>��r`,�Ŗ� ����ڮ��fH���s��N�8f3b��t"���pI�pb�*��r�u�f�b�� �lW�5��>�|�ą�+���(���"&R�y-�d���H���@KoB԰Ocɲ}5H�|9�~=��w�:�M�L3�*�aw4��ɐ-��+�hLE���<���(�1��DC%)䲻H�^���'V�	@�a)��zG2n5��H�<�J�@�C�'h�[V�
{��w���y�dY{���e����^R�=v8����@�ޭ0�d�̅�4�~
!��z'�rטUQ|
^���!՛r�+'��4�/Xd�ڗ_���3�4q�{��<C�H�����[���@�`��vGM�Ԍ�N����L��]�1��l��� �2J�89������N])�@C��jZ��FŻ:ŮX�c�`8"��ҹ)�����i�`��i�Bx�ܻ�w�G�=�#�Nj����Y�S�S&�;����/�ۈ��v�b��t1�=U���z$LGnE�`��4E��@��!~� φ�ǬW�b��(U���ޔ�fI}��%�Q���
���� �|�!K��O�S?�٢�ӌ��)��.�$y�ǧ����ڒ?��+▴��ձz�;��#q9�Iq���f��:O��1�ԋ9,�D�����L�#j�gM+��r'`o C|6��Np�fm+�x�kr[f�#���u����ɟ�x�dE��Et�O� �ZJ�E雐Yl3�e)���@��Z9A]
�׍F�O�h������=F�$1���@��|�g��_�Q0mF�팮�E�؎,K0ފjZ����sW�Q�2h�o�|R^UU�?�۫X��Ť %�
�t�%�6��I�Zb��k���\�X�N>�CT-C8U��qVyD��˻!=#^ �)ֹxS2�hO�����v\j���ayl`���spK`\ƾ!�+3�[�k~�7�Y!eT�ρ|�?�G�K���������޴_1��u��F5�=@��>5p�S:}u8��1P��h��Ѳ���o=;E�'�6kỼ|Lj��0sD�be:�[��m�3߳��=�i������'F[bLI(�A�%�I%H�@�<����&���-��ݤ^�!h��`�ib����{��=Z�Dn�
p��G�s�Uo�(��K�zKل�j��-5��� �����Wo## �L�������k�h$`1�.\\7�fE����U�\����X�&TmߤF���dO�c��R�J�RU�V��Ū�3֖���~���O,G�ȁ�}�u-��C/x���M��(�X�9�g���#쉴�	�2 \��"�c�aSZ�gm4 �a�^�,�2a��]��\�Jf��Hpʸ�j��01w��q''���4��<��<����p]_�,f3u��:�ت(�޴��C&{�":�U���R�� C��[���!�<�3&�����N���,��NF��MZ,P���7�Ͽb3+�CHQ&[s:��%�TZX�͘��I�
?[���$�0y� �ua���Y-e�w�5���'$ ��8W+?��ܲ9��XҌ�џ�D[�r�2�"Աݧ��CV*R;�q{y�`�Ǐ����I��Q�!��r�e����}�����n06d������17���0C	��[!-�=C�EG�cL	��-����+-5[S�L��,�>�4����lu�y�zWӡ�!�R��G�|��lt��։��@��x�"��m��1���$��	r+��
��I'O��҂u'�����%�a1����i���vۣ>�ܑ1d�ݠf��s���K8p4{ʊ��~��>�ӆD�蜢"Z&6a�X�c�5K4@�R�����(��!Z���1���m���/�*�W�ӷN���|:p�'��<g5A���c���d�lq\D�W�[���d���.�x���PΛ�����M�7�\VBR���	�ت��J��!�(D�D�	�	���ڲӋ����$(۽������L˪f�"�--�'Ӊ\Lː@���ݕ��$5��0�� ��d�|�X�::�����wC:�>���W�P�s�M �������ㇹ^n3�3u�h��������su��s=���E"f���eFb��"���Q�����}�=��;��~�*�J�7���Q�e�jd|#���) /�l�GS-d�fݣ,��91���o�M.��Xـh�H���V�E�`��#�2�*ֵ�jvǒ$}���J�$'�b�M���N��:�,��E�c����Q��5B
{�RsoF��IC_sK
�G���L�w��%�g�)��K��� ��^��@	L�#!��� �Y�>>S�(������4���XD�0��9+%���'��i�N���.Tu鄯�q*�-�>��t5[�ܮ���
�M�vK/�x�oi�9��IN��:������[כt +�l��s<�~;�V��#�e�⏡QtUR jR�t.b�0��,-X�TXm��fj���d>Ԕ7��ض����d�1~�0�;�c�]�Ά�&"��c�:�j�V���
*�1Q�]/m6���F���`���2� x0K�QL�Q���iݾ7On����O��<c3�ǘ��W"��{�����ƃ*�x�׻V?9UC6�n@c�ݡTV�~���V I2��ѧ򥟚]��[
�N�^��n��8��)?D�;��AI�]x���v�w�W�Ϗi�~��Uu�#�ď�U\�E�%�f�RZ��ý������#��n�����%���ZKq����v�UW���\E�3���3��� �q+��O�V��+�`����T��;S� ��?���	�H��I>*�����K��p����2�)����,�U�եI��=��T5���R�>����"J����c�����Z��..~�6W�r�3'L�̏�E�y&ib-�㺰��D�7X������O�To:�1f��sw�Ѿ��ش�D�c�@�U���8@ �l��l�Og��W�E�|�q�����y���,$S��U
���xˮ�K��X�J(�PR�R
t��^��/ڂ��-nU��c-b�CL-������E��]�E��@�j�Ph� �tY,���3~�����U�IjB&l(�;��O�Mҧ�g�E��"�М���>������ʦ
�/._C��z��[s���������YK��M�!����_�*4�fgOv!�e�?���#y�CJʁ��ţ��n����:���Cr,�Z�Ѓd��?g[��G!�v)�BL"^�����8N��NFOL���AܰA=�WNO}���h!�_Um�'dwg�Vr����q��q �af��(�r���
@#y��/E��P��<��j|�'��|%��&6���(��_y�m�c��E��A����:����#��J	B }����W�/KS��uV`T�Б��Z?��ܣe�O���v3OA�o� �5�;E���v�m�Q���s�Ř���:�#L�E1���/��s�<y���~���2�0�d�����+���8�h��B��f�T��H���K���К?	o{��rI[0��rS��m'3�3�o��s��1 �UҎ{��7�Y�����|�-��^��E�/�
}�g�3�b��֫r���<��Ɵ}��Q�۔II��I�h�U~�kI�l�/��a�u�B�<Y������%����f�%極i^���ڹ �����lv(�<So�aV�"��bA��#ϡ�Z��h�
��AW��B��_W����?ς݁Z"�G��XTᙁ��xöI�	Rw%�B�S�6N�U݋_�����
�1��q�,r���	����ڔ�� �l��GjF�j�&$ҳ.����ڶ�C#{½�[/w�ȍ橌��W$ ;���۶�b���C"2�2qtpj3�v�}��}��w�V�IR�2�Ye{ e@��Z�PQ��<�`�Z��� �g 2�; ����V\_��ןy�56��[Em�.P�%1��c�"�*�i��u�9�*�Yi:�i<��l+�I�D]:�=Q���h|P3GN����H��z�f����A�b��u_u�<�4�'����_�%[)�|%A>"��DA'�{-�	j�ױV���l֠�yË�E�r�A6��}˺K �-��c&C�Ʌ�lV]y�:�b����T}�m8N�iό�/���/�%�~�O���{'�����s���o~jf��dG�cO����m��L�d<n
6!&����K����D����b<��pW�&�0O�����w�����?�
&���h	�e�x�A����ς\S�a�SKy�sO�b��]2�� 7L�9;�[���9sS>���?O��	M*���a4g'�k��y/a/�e��8ԏ����1u��g-�G�ۘflj�w����26�� I,42��*J���
Z$�?%W�����p���U#M=�K�������-�}Ul��r�_#=�蒞� ���Ň�b�Sm��Q8G5�.�:��Yv�&���wj����tk�<������2|2��1=��,�洰z�+��8���FXU���3�%"�g��]3Ο�f�<�t��I+���r�3g�,��������	Vy���ƁP�.�>���,-�=��{��tj+�00lW\ASu	��b9ޕ��}�H8�7/w�C�\�����{�� �!m�;��AgG�A���<�Ȇn"���O7i_�?�դ��G��?�-�E�������u���E��$�0�Y���[z���_׼:�9
�%[����Ok�5BSūɫI������u��D�3���{A7�f�L�#��4���%|��Do�?oE�ǌ�A1�^�����/�DHf��<ao��	<m����[�_�[:LM��؁XL.2C�B�u��%o�=��p�(���yh��$���#.���0�����S� N��M[�"[@���{�>���º0O8F�Yַ�9X��T�l�xb��O���F�Y1�p�O[��?J�����Ԑ�1 �V0#2��+гS�`�T(�Ψ�b���H��N\�ů�La�Ҁm,|LX��A�`��w�+Z���C��^���=۱+=��:�����y�rV�o#Ml�ݻ��n\��۶����{%���j�h�6���w�c�ւv�������1a=��E�]���
>AKN��s�m�T˕�)�M͙�n��Fi����p3������إ'�����e[u@��W�0W4���t�X��FGC^�!�<e܉QO��=)r>弦�$�r�O�o6EÚ�|��c�*��C��ƍ��k������7���$J!'��!�c���|
f��Irx|���j�c2ބv_˦�|����x�r$!p��w-�[�yS��y>�?�����>R��r�w�VK�-�ΐj��8uX��
�m{2��g)�÷${
�#@<�es6w�n+�VO2�\���G$���բ%��)e�`�l7����"4^��'\z��I-8�o�:��9�9�zƞMC��#En��*�)ɤ���Q�}�X�.��2��k��ҽ�do�[ �o��C�� ��<�Q�l�DA�z��/Zى� �P��`���h~\$D�\�P'4�;��W5�3ܢj���6��( 
K�Wn�'VGB
\�޸��Q�F�?��'����	�1��:Q&�+�}�2a���s���^D���?��ab.�AfQ���I*��n��g�d:������)���ȡq���gOF1(��l��Ǫ�z��%�Q�h7MfA�K��$hq�3���h=���C�i�e� ?����Ǩ���4 "����(Lq�U��C�&4l�"vso
�RO[T�[�N� 4Ŭ{����xMk�����ei#�%{;l8�~�1��g�\5��S/C�`���>�N �6Z=�!"�SgÚ��A>Hd���؉��N���ɇV~Jn���nf�ɸ�̸ z�%���W�>��xɩ	�,5�T�	��ԺQ�Za��ݹ�@�A� �E��g���^��t��^5�_�W��-��Q�.%R��VN�H�mF���������@��я2_R�T�*-T����T����M�smT�lС�`m�ݿ8S�����k�a�5���賛��/����yu�J0���&
�DRۼ�&���<"���q��}.gt�a�7�+���X�R�"�݀�&��j[Z⌻��!��-��y�8�� �+е��O��a;
�:,E����� C�BHW��1�������nc �5�ǭp1����S�S���~3 �u�7["3ii�|���6�h)����ʇI�|�r2�H��Cf E���L����`�IXr	����';�p`���� �V�k��)�Z>���2����w'wXؠ�ml>a�L����9��~���!>zS�o��y:t,������S�����X�fw��0���3�[&�������L��>)��-�؛���M���S���
8�h�{WOv���b����I��>"J,	�]����B�6#[J=3����Q�[K���8'�)��<�4�ߝ���+�fI����!��� �����̩gx��v�U�gX`��EB�̵�6����ǆ쭆�U)����ҟ�!�H�Ŀ�)w|�F�*:L�i&�aƮd�Nu1������'�9q g4�Z���d���O��˟�4kYF�t��>�Ї�2�Y�u��Iq7�������	�����o�S�u� ^��9�wq����&;��n�����t{ T�x�e���A?�>!ک��ܝ�cD����ś�)d�j3�S�X���LV2����;a�bQC�kP	-�ɾ#�?� 8��Y�y�iQR#B���
NNm/�C(4��x&�/��<��[�e�x?d+������lūR�;�f�*�;;b}\P�iCK$,��}���oDow����Êc�}�����R��&SW��1\��v�'U̎�X��g�3�$+�
�"���q$	����a��Ff�&"Erc��r�k
J�D�P+R��`^I|���q�[��e�mY�����{�էю��jX~~Q���.K:��6tN�m�9:��Fci���V����xr|�NtWEl8f���Hǒ�1��j����j������92���X��Ӛ�����V~���N�R>0�R���WuL�[Q��M��%���K��y�r.$�)^��"O҃�h?4#<�a�>>fi@k"Zm��Q�Cc��/@�9��;���O@��Ba�<&��^*����	AN0�l��V�I���֘�`���Hp����d��D3���F(�\ny�b���Mi��S�U4��`��䨦$z��]À��|y���ӳ���;�M��Cv�H^���<�e�?R)|���h��/�ԹH-+8`c��S$��F6@�V(,=�rڣ�pn�#��uw"[�]H�o0��պ{�'��^�W����(Y�M��|���.�;�ei����Z�K�@��_#�8A�$���rK�u{�i�����&��� ���ؔ[����'�]<M�8z)޳X |[��{_�N)i	�Ħ$w��4� ���A'@Σ�[�zϽ|�%���OK �l�OˡZm<����Q~:������{�{Ko'@��<��RT��C�ƴ�]jD����s�A��*�B�Q$��T�@�r�CtID��p���Z.��O��ev2�
����e5�X���2:�S�����Ի�����-��|A����E�P�J ��Pʼ3:�C�I#���7\}�@ȸ��@�,��ȌV�\���{ 	u�Zљ�1�����B��9�Z��E$B,�.y݆�b�VK�Ji����Gm�C�#k�C�>]��b�7��+g���І�$�n�Rc�y�:��=��gc���g�r�&�����8 LD/��^�PKre����r#����K��<��X�^/
�j%�ɡ�K纸���,��r!Q�Lk�[�ǵ)�w��?�?q����}���9e{��>\e��O�MI4��=���	.�ҋ�^��$6��Rx��I�,�L��m��<��Z�G�?�}��S�MN����D~#�R�n:
�L1�>"XI��4̶_�Rj���8?g7��wA���\��K����K�Y�"��u"�U���8HЗ<Dֱ��#�M�JƗm�*� ;IA5�DS��n=���*al�0�T9�X&c��CەXEx�y�d���4"�8���iC�
��.��¥4�;�*��ڛ�~4m��ؒ�[N����|�)�]&��R� ���Է�Q��C��?����">��<:[a��.�;96!�r�c�X2�ԏ �L�e
�9�׊���/uZ�����v�:|bh�H��>���[�8<T�|��~$+7��`�'ޱ���ܑ��- �Z�1	��M唗��^��⸨B;�t��ڼ^��M��>�>�
�2[�w6]���k�<�%$ $.��k�҉�nX�^9?6S����w�������x=r;�ȓj41��i���i���g����Wj@�諎�ܟOR�BL�{���u��i���|��	L�V0T�����"�F�c���rBUE����|Ɓ�� �(������sϼ|���ȨK5^N F�cP�6cN�'o�B��,���n��GPw6o�d��!<��V��<ICU8� ѭd
��!���s����*��J�O��J|_�L��l�b�8g�@b0�5"5�6m�0�><\&�wȋ����)B Z	����o��L�XO�re��|0^kjh��?���4𒏥��a}�6��`�~�����a��8�C�ɮ���8,�o�mI��it�����Ìh�������.��+?��2��A����UF�;���,�ԍ���Sn�mePz�Śƫ��[�Q����ط8��@d�����'��9ЏXA�!.��[���MB�6��j�����	Wb��<�GZ��V��fm���������]a�ذ�7��Z�ݓj	�Ҭ���0�9b�C���>EZ�����SY���HE��R7���>-�*(H?[��4u�ƽ�?�� ��T.)�7=_����_׷�
RF��\��-ٸ�{�ג|UD΋Zfo��P��'O��Qw�z���vRi���,�|y���b]ˊ(pg"$C�&�Rԟ�t��S ��Û�p��G������vV��a����P��+�;�:I�0E��h m�U�fJ�rY"�jug�a�]���w������:~�V�Ƃ>���$�z��A��Ё(��9Lϴ~�S'��5w�ͱE��ﾉ�2�З�ۼ(}r�
���Nұ��@*�/3؎Q�n9�w�%<��r�e@T>�G�ETI���lg#z�Z�������]�uFi���,��Owh[�ѐ>�>����o�}�����B~zD����
��W2+p���>��kL���Fdr����rc(co)�lC8%!\ K��W�x�i)�U�~]�~~���#����A]x����C�U�C���Tq{#�m���I	�0��,�v��!��T��|7�Qd��"��Q�w��qZQcml��X
T �����k2�OH�1}���KZ�O_¨�#3�D?�H����9)VJ]�?�FL7B'��#[/�uH�9Z����T�j~;���d��=� l�]�s�6�c����˯��t�`_
-��?!��j��u����E���^�j��&[��;|��IQN�T�H�k~-5�={�~�\��yc���!H�6���<�MQ��ԓ�3yi���ڴ���i�ػ"X5s��؟��&����C�?���g�� ��̑8��>��@����u��]KӴ��ƾ��K��'��?�߄��"�65����3�"�3�U�l���M�Ch�?A����	�0�zY'wk�b\�{j[Y���<gw��ag7`���[c����9W��ۙ.�!;۴T�4씕e^��a5$�t���kc���a����&;��I�Sr7��k����s}Ֆ�*�����%&r��i��A��Ƥ�p������=���}��)��_�7�v�2�vJ��У��Vξ}�f/2W	�%��``�=p��hm;?��B�\-Tq�|ΏYl��sT~�� �Zo�%0��P@o\ۉ��:�wĂc�M9'kn��^b,�q�s� �4���(�m� G��H9�JяE��*���s?�����6���J
�d��|
���uA�0�I��B"�s[�-�v/����լ&֑�3�x��[� kf �a�*�΍>d��b�����Q�8E��0��,N�el`a��].Z�-q�{J+~��~�~A�T�0�x�g�k�o$�$M������'`qmŵ����Y���T�<���l�h�;1|��Xb��T/''_Ǐ��}b5@�x^SA;�2	�"��&�%��~*a�?v��:E�95�K`=4Fe&@�'��auź���x!lIa�P��?4h��Z�`?O_�9��.[GK�< �s-	�#������A���)�y9�	4;|�N�O� d����uN��Pĝ[�!�����3aN�����>g��8(�T��v�m�1�ÓD�.�=u��{ ����K���+�
:�'aGdN�L���cז-[Db�y�G抂�ʂ�f�'1��!P�y �/aK�DD���⏹���������.�q��O�ɛ��!W3��p��1�^�#�f8�Ѷ9���O��άL�'��Q���c����\��]�٦��A������V[+zQG��B�T�Ė���s7������#Wz�䒬�, 9ɞ����~����z#����ʫ��.ө[�3�n�\|�����˹�P8��+5T|uw;0`��G����urs+��c�6Ж��a��&wYə��#$o��z��Y˵�5��/5�q$�\��
|X�������m�Q�	Q}�L��2lA���h��B�m��I~�\�PT�_1���
ߜn�!t��\!�ʚwA��2�Ңځ�,�!��*x��˴�\����BJg5���(U겴3�#��C(�Ѕ�G����s�^�3����"(���*�$�4<��i�W��x���ή��&p�Mfb��������A2J�4"⻭�� P͋���,^,��Ҍ<��� P$����h]+���|"����-�T���X/��[)�P>sY��-��ͼm?����+���\?�d��el�-C�%�j���fѺ޵�YA�9����/�����he�B~�:����H��j6��8��2��t���s6�ZE�y�P2J�5F*眚)ِ����wt�;Хy�-����k��@��͊����\w-��f�Y�p�ɲ�uJgiQ�`)l����QJ��k�<���,�c=lk����wπ��"9{��٢�o+�Sf�7/�Ԭ�K�;ߜ�kz&����� 3T_zt\��4>��t�x�ϕ[�ʒ�~��٩���Z���C��3�(�\�Z9��A)�+��f�����=_��L�~�լ��󋚽��cq�Û���TK"3ł���vV�<#�4��Ty!ѡ��|�g��nM���������0�_i�mk���ñs���'���=~O���~�44����:���I�_�bW�z�
l���R	��m�� �̛�N	��,%�����-�x�t1Hg��4�al�3��p��m��C66�2%ծ�m��J6��I&���*�Ì%���u�J3RP�������t���A�w���.�*QcCf��P*
���3=���6�#��I>�px���u���佲�
6 YE�ғT����s#��:6�;��?o�x����)�<��Խ���7 �l��P�l�	�<�"�����&_��g�h���߽zoj�+��n���<��,v��.RJ�թy��l��	:��{�v�Y��<�J�е�Q#��U�>Nm��`�x�׈�e��Ec��ƄQ1v�d8����q�`�I��|3X��fEۢu��u��Q���sD�n&�xu��i�x���{.q8n�n�]��|C�:d��9��u������Շ%]#�؝2�V��P��m�j�Hj�~?mu�����`��D�#�3<zM\�� ��$2�� 0�3M��u���\�V��+6��&(Y�n��u�x����,z�jN>@X���n�X3-����9��-5�+VΨCqbg!&��ŀDC�:���(��{�?�3G鯴���@���>�0�n o Y��@�k,���7.�*9���E*~eP�����Yf�;]��Ysy�6���� �^���0C!O~4r�$�9M���^[J�JH�&�K3���`V�/1}�o͛B/܊�� ��-�vrwE���AY	Bhv\)$�<R��e����y\���r��j��at=_0Ak��h��(N>h�btp$��N��mn$�5�L���2�h� �����YjOv|A�z(���0FZ�����ʔ撁J�]�,1�W�����4.�C��)TX���-��ŝ
+���,�R�K�s�	b>�t1���=�,��q����!u�,4��E�x�0��!�����٥�=�Η��t��z@୍-H��ʓ`�\R:�=Pn/^`o�OwP�a:{u���<�2�����z�sn1��ӈ&ڬ~cN-���XD.B9�tI�Ǝ,��N��ob0kR�ܽ���u��5֥稽3���F�J3�?X��LQsx��(�n�i��7�(�~�WҴ�B�Tp��Œ x�X�m1q�����[[��`�Z`s2)w�i��m_y��8�=C%�@�H�\\���M�A>7��~Z+��\(������Ctb�}CR���� D
�B �eWq���.�c6������tT16E��j����{m^��i���a��a�!�b����d��!ёq�t＾id۟z�q�5��5�I���,D���+?Q"��k���9��׻�`�����eg��k]Ks���S�D���iC`EJ���>1q�vPm`̻�5bQ�~Ѫ˛t~,C2�����>���D
�����0xL�y���.g�:>�7 pn�����kz�%~�p��0�l���P'"�.}�Xi�U}@!˴Z�ϒ��P�uKF�����x���B�7�2�t^�#bQ ���������0��x���
B V/�U�~��_�ͪp�ݐ9l�_��0����ZBwW.g/�
��|���6u$�ULyeDS��q���������Νvd�7���enL�jDMOGwɄt���^��(Aѽ�����N��p
L~>�JH0�#��`dW��c@��S,b4��E�v�L�J\��Y�Ν��W"��̩��BN�bs���~&v��c�R����F=��&�:�`�u�Hrf|����'�%�{�8:�p+ĺI�ڑD�S�:��_긜6�!;Jj�.}yjF��L/�Qqt����$B�tq��G_�Vt���
e�oH
BHh���D#\�
#4�`�3�b�qa� ؊ɡsc����g/�ul�s���-�ɏ/�@|?bJ2kWsG�,���*v��N	u�%�)Y->7[mS f��`Z�>���!6um�V�`������5���S :4�9/�-'��,����π|�X��>��}?Ջ.��O��qk���g�B�Y��O�&hə��.u��`�~��*�b
��t&�mw���!��m=�$�>�I�$����-sc�ާ;��r������TCu�<�_s)0�nh�<��f 5oӏuc�)�G dv/�]V&j_2��^�r�6��%���'7[A�wɷ �s�^KƧ(DQw��'l�M��4��5��S���ς��c�M8}�@[��6��^:�)No����7?nwg��@k���nl��1⎓"?�Vkoğ�����#���X����=l8��|�w�i�ԕ+y�D���Tjw�<���+&��3H㌟nw�I57�b��9��;C�a5�"�5��� ���Ǩgݚ �����	�� c�P��͓��3��m��^�����B���«���L�c���'3��#Q�oTK�z~�QT��:���Q�!V?��L5OY˰58�Ǭ>JP7��S|�񎠳�
z����]k�Sa��[���G���q�{=N�>C&�G)S�2���+O��5O��0�������T�m�� �j�!��k��az��V�`K(m ̶H��m��zj4�Zkw|~�d���d�vߟ���,,��FZP�ƚ��6	�M9���EAp���j�gE�~����Y���5��z+.�G<P�#G(3�"��3x�礑Ѹ#5<�v�d#Z��ޘV���a�.Ó��F���<��g�2\9�g���![�^��.���*(k��V)�(R%��|�iZ�z���ۏ �P��}ӓ�I~�o�f��J���w��t ߆���b��9�����Qo0�c��ᣉ!��}0Q!���j_O�	L����%*�MA�>�X�VuS\T�_ǿg[��WoP�&pC���0���^��Z��<����joB0cο�"+�ג�1�[q4�@Ƭ�k)N�W��j¼d¡�t�n	,}oP��?��	���4�>AK_[f����$6��jq��q��Y�������a�\34啀�o	��K	i�s��
UY�'��:� F:��Z�Vd`n��!m���3>\���|�!�"�T����i��c����5L��J��vg�{��`�������&7�q�E�����U��2]I ��T"������y��9P�a�t?��xa��$v��l�'Ӫ��C`���<�B��;[�͠==����K�F-p;]W}��^P�	XC?��e��
���Ə��m}�+�A �Z��F���B������=�<��,e��LHmFq_�=�G�'n齻�?��|혍��Y��ny�I泯� /����L�m +)��Ӑ�[������ySJ9Q�闼���;���������oH�$��9��R{�y���B�l�vj���H�/��\!h�>��Ak����P�������us�e�q���/���A��K �L�Ҭ�.aӵ³�b�R�I�f��2��MDFm�{�q�[3���"�Pul,��^�^� �@y�Y�iy��i���lk��DjX�gU��F�t�_!�\)#�͐]�R�~�_t���&)I1�g�Z���V�e��~#כ�,�yY�Λ +��i���R{?�?�o�O��-DcN���k�*��9��������GX��4�*�m���1s�@N:V8�Ӥ��A%]dR2M�w��ޣ@Ҧa�D������4��ꢔ�u�t�c���N���R�-���,5��g;�[U�7׽��1����0��P7���)(������}��@��:�D�����ĺ�k�o��*���5?��^�v0W���W�8���f��j,�Z_?�� �x��2^BC�.��?�5zb�Ω�e^�A���D����[M'���q�m�+�:m{�K�g�����ՅݙV��y��3U�!B�rcgM��Z2�&�R
:]���ڵ����]jK���KR�oĽ٪�(�����N�Ǥ7#����_�ݢ�@9cz���KG���;]���|��L��BE�ҳt�L����:o�n�J����{	_����+�׿�&A�Ub8�0�yo��W������x[O�|3˃�2�߳�#`�V��4p\��3s[�	-���/o`1\�/G�hBoV^�X��_,|գ���ks�_C�l�q�Ei0�����՚R+�):�u�Y�eY��1���"�m&�(h�T�� ��O\?���J�K%�k���Ws��CZ�«k��Z��@�2��B�j�|�N�6e�a]�pu�/��[��L
w��/�#�4����8w��D�[?ilk��I�}��3c�'�mtb�2\�兽I�I�΁?k�w�Ӡ	��<���!�Ն�19��ꮷ[,�X���)a<|*Q8���RH�ȀG1P ����.:'�b�#��n���W:���4 ��|m��Z'��뽵)yt���s/͊s�,D��fe�p[�����~f�t��,.�>��Pᐛ��\c-7c���[�6���as���y�l�;
��� �£�K��`Tc��l�`n�����Y<|.�Kq�D�����0d8��T�D�;�h
~�l�1�ȹ_5+�l��S�j��� �B;��r����=�W1�}R'!���mQrg3K�+ �\�#qeRa��.?��۵9������
'G�9+g.&g��˰�T%	
f����ƒ���,s�������QHu�)��Q���8�Q�kT@��y=�+Yٚ>T2D�WhV�'!����arғ�>��f<�Cpn{V��r�P-(VYՇ���^�y�=��mQ8��:CG��br�|?H3(�Xn9�2�J׭�	Ow��1�U	�{��rvC�T����[ye�#��:��G5k�f�q�\�;�[ɥm��ϗ�bcd�_� �f[ �e�~H�0#>�xܲ� �*����[�7�����m-L;Sx����PNo���zN�py��JY��f�RXκ�:��T:=�u�=�}���>��
b��!=����|�|��:��C��
>��G��~T.����Z���3K�>�??�b�*�R��*��@w-�,�)�:��4+�ߏ�����(��_���wB���yI�Zk�0�5���$�����/��ko�l������x_�������^9tq���={=��od�Tj�](P`���Ί��@Yī�>P�"��C��
ު��O���={O�r��+�p��@�k�ş�;{<�N�t���={0վ��p��(��Pʕ`ܳAQZ(&�Bٴ���␩<�۶w<R4�~:�o��~G�K邩3�>��a�	ɓE�ŏM�( ����.{��-��������ֽ>]�6!��x��}y�~J�F\l�pO�^`])p���w�gG,��E�)�'�ci1�M��������R���?����mC�vÃ�D?Ŕ���k9����x�=�H������;�̏�_�^0x� �����e��Ɛ*OB�w�u��&~M�.a����o����(+ڡ/Erl	�I�B��uAB�r��_�\�������P��~��< ��v�ɵ-�Z8�g3,ɷ4?�7��ߨ�];�|R`kW���W�����m�q�`�r��i���8wM�{�M���n�%y�^|�Pj��嵲A�#��:���O�c��L�,��-����U��W+�ec>5�b�`�i�OrQ�v��fH���p^�^\�R�=��nB�� )�a!A���No\?�֕��TK �b0�q��Z��B��ew����aD�_��\��ޝ�{�t�K9���BLx89��S�(8�?z,�Rє$�t�1W����Ĭl�e[><���9�1��.񳗾��Ee�b�g&������wz�r���7E&���]�($6��yZ�K��QA?�O(pY�А��|�d�����5~h^z	�*B
9�����Z�s�i�P����	a���jf)>�� w�o���@�+���b9Q���ጧ\dVl.D�f���H�Pe����-�{���r����QX��H��^킽r��@QN7��}r,�P�fݽ�B�&�"��>0�����'�?�B\2O��綬1������])f��j�4�.��k��`B�����	��q9ܬ~f�5�a�G%�<�帀���e%����JM
P�������!�����{y���ezf'w�hI�'�5ע�c�l=���6~��h�H\�e��z�'E�/��v��+�<�?��}\`�]����h Na�zN��L�G�-��sY;a�FӺn�qh�#���#	Ɏ��Zű��0ِ�˔�2�������_y��0�}a�"����vpB5� Q Bm
�h��M �+5�l��c�����������SK�1�h���,��i���'���?��iJn ��"��5�T�gl��3Z�(K~��(�������\����s����M.���7<,��(LxH���uP�ٽh<�>ڠ
�\ƻ�,��g�(�v��Xs��
��@�S���U������͡E��v�7)R{b_
m9� �:�F�4�#G
o�}�n�F���%�'�����YAY��T`K�0�?U��c��ڑt$!�Y�h��� <wK]v�?SC���PF�;�7G�j7�唋ߎlu[�'�De����j�Q�+1LN,�3�7�|^Q�$���1*�p��k*��8�>BO�Q��t�_��J���R"�Ef!��6��?P�X|��#�v��;�r�������K��
U&B*��y=j����tĭ�_"�;��§0�WׇeS&g`Cަ�T�bM*�w<N���d��$�9��q��͛1j�v�	����(�\��I�$�|/�4s�EäȞՆ�>$&@��p�Q1��6ᕧ��p� ��`bSFUᤂR,Rj�X3"I��U�b�!©�5[���������0O�(1��'$b�O:g(d����Nb�z�`�L�C��{Q ��r��ߢ6>�[+Ñ��ú9��ujE�F�acE��>!��of�m�-Y'�������3�����t吐ll�p��������mnl���~ֱW�G"@|,R�[��4�z^��tiy��q|Yګٶ�����}G�2_K1�K�>Cǹ��/��o�$�ǻ:���V)pF8�0F�TV����8�6�u���+^�Z��H%�s�$6+ok�Z�(o�q,�����{��&�����zHr:��i�E���U෇��[�Z��;��(ř1����H��]���ͼ#��O����8��d�!��X��Ȁ=��m��j� �)ށbI^G!�h��rXj���W�H�w@�I?�}���] �Z���3>n��uK�ە��=ʵ���Sĳ��~*܍��[��N�9@[62ڥ�6aK�%�]e��71��g<Z��D���v�3�G�w��l"�(�pS0��b��ni�*y�7� �JN� B״�Z�p���{j�/�Yk��Ps�D�:ѕ}u�m6�	[�K�F�<K�B���۫������)Y��<��]f�V�_U����ˈ)���cC���Z7�*K�%�h�{�6�H�m���+����+�>t@��-ݏ��Ҭ��4���ǭ���o�u�P��vinЫ��b#cuS۷�Q���e��� 8������`�f�\�1��U3C?�$����"���:���0���K�{s݌8�??{SK����nr�+�1D74�d�R.\͐��k�����p|^�C��[��d�E8�05��1��Gq!?�3PAh�6ι�P����B����%*����$h��{~��ѩsq�?@H�{G�W��%�0�;E�in��:º���Mܯ�5M�� m������x��M��S�����f�n̥"��3�<6���A7:	�*s�9;z�H1J̓{.����J�'h���2,'���b�/��~��7���ϖnR�̰/��`#�iI���Jp%�m�Ld�J����}�h���zN�Sb�eXӘ�g��-�a9�֪��h`�E�hT;�K�>~E�=hF]�+�`5��R*p�k�`�ޠw1��چ�I��Y'�%��xvK�z,>޴�H�c�4c��+@����[R�1�R7i�]�h���B�<�����y5�m���)��2wy�WvTw��$����UՅK�caY:>4�RUt+�7��������z�ұU�a��J4`�� 
�q5�M�VP�dT"���X,0؄|���@��ƹy�����g����3��45%ݠ
=��5@�ʹ�U���	�Ħ)��o�y�Ѭ%����1R͜���r�e�����Bt��s�4.�\d=ř��ݿ7I��Z�5$-��[�s4?���T*�aN�C�1�O�Q(�ݵ�f"SZ^d3$k��N���5�T��`�ݷ���6�8W�P���!x�渻撏l�.A��Of��19�ѝ�(��oí�L��i���E_��q��
��##{�p[�9/�}��5H�3��dA<��Ah���&�f:�ނ����(�Uc˾�kLȩzt4. ��0�dt���v9�3.k���{�'(��f�]<�BqWR��i�n�{*E5���Z���j�-�tƐ ���:;lL��B��c����㱄�gh9��X[pJ*�Q��A1�����e�`�f��b@�NT�h�n���?�}�H���C����Ar�����"��7�B�޷�MQ˜b��L�ൂa����O#ZWwA�A��Ѽ�!=F�)8O�1r�	7`��m#����u aЎR�xb��*�4)�o[�hv%�Ee5�l*��D�l�iJM�"`����<ޗ�aB\�/�&��?*"�z��K��W�{K�zs?��O �ƙ�N�vXE�d�!���vn�\C8�)���܆����zgepH��h�IBLhqӴ���&�+�g7�g/Ku�!�h�lh��[�voΙ�֊Wm����� �lJ���� 0\�����}��F��i�?C��k�X��]�Iu�p�J?���ƣ�MB\w�lS8��`��NʚO�p��a��{ce��g�:�-)���uq���'�/DT��fg��BE���p�|i1�����S,f%^d���;}��=l�Kzm�o���I<ޒ^m?�
�(a�MM���ł�
GK���k��ShY�my�	._Ƭ�i��n�`qӜ��]<7��z��M�ܯSN���l�#�Ƃ��eڅ��Z��eϹt]"����.|�i|y�o*�����*��"��I�4�7��b=C���]L�s� �a�tLZ��8M�6/��BT��C'li�j>$���Ũ���-c͗HfL;��w������Ӊ���C����A}�6 Ek��ľP�{���.���[�� ��!_�A2��㏨�*.gnI>V7��p�����F����YX�p�Ơ6
��Y� z>^$�{�n7J�!�����N->�:?��&(g�Jŕ��~0P8P`�D3D��>�Ѧ}}���oڍ�3���+��1~�?���u�����b���!�v�6� �-���8%{침��R�g)6l;D�=����{���f�����Y%���L��/ޭ��zJ;lkW䀁K��a��N�v�;QY��n��&�8B�ۤxǅ��=J`���F5�E�6�Q�q�-����>�şى�9g"������u����eP�>S�����I��Dy��1%dZ����HwE�5?m�?���6�d����J ���Z�%>�P?��X|��eA<?8a�Q�`���/�r�!.ҩ�IK/~�,J%������E6/ۄ�o=��Ez��Z��d�;J~7!9��?c� )��li����e�����1Tc����u�?\gT�0�s�(���#�l���)₼@Y�{Rw1�����[���h���- �9�k�4��1"8锟�E�Wn;Ձ��FA����1Uc��q����]a�isG�Z�ԓ+�}�O�(a!���Y��6k��œ�߻#�;JJŗ~�����@�~dHҺ�$s�����+���ܫ��S�c)M��?�5��L�{�j�œ���[F/޵h�ˇ7��
�D�U ����K�f�"�Z����La��,�ZĐV���g {���>%?�N�]����=�8��0x�vO��K�[y�dW�1����a#�!�F�A�Ҹ^�po��Ӟ{���&7�H�^'��,|;]4F��_ �1���D�y�f���l�+G����Z�{����W����S���{bW�ծ��aj��G`"�)�mx����_PC��hf�gQ�c�]���þ���Aq�A��ӡK�/�	<vK��ٚ�����AX��КN�$����:��
�sS�ʎ�BXJr����~�\�R]y�5�V����Ӳ$7�:�X<�z6�۟���o�KȃU�Á_KF�%�r�H|$e��IRL1+8��MZ�ݕ����D����?hPE�5�}��mZ����>}���T��b�=��������z���.п)�����2�M�h��m�-w�`I Ě�ӄ@{��]���D̃���$���ࢯc��0n��6\�읨:�8��?c�g�S�J��q�q�>'i�X0i�$�e���8��owٗe�j2.�!�U��X�I���
���U���.Sh^�PA��J�W9�>�w�<�$�i�I[�b6(��	�sB�: p�B_Z Ԇ�H'1(�0���$�������)�I	�@'A^��º0p���>/��{�I@[��i�"�P�9N�+������>|��W��J{ J���h׮���f����9��=�����am�.�0p`�*�OK&���2��5Eh�mO<��]R��E*EKv�y�E�u����k�4p�����,4��R����i]�5T�T&^X����L�/���vv��1+80��<�m�����<�3B��S�t�}�]��5y�e{5栾HR1~)��/�&0�\��?D�{S�AW[������ﱂ	��ߴ�]Uh����y�W�~Dx�P�2�W��+t��U�Ȫ�g�r���;�L�ќWB�E�uL�$��L�Yp�H�� 
�E��N���Ҋ,"k��&GM����
�c�|�K���ɋQ�^�a����B�I`( c�S2��-�h੆��`t��[��w��3����V\6�7��M�w�G�{͡�$%dg7MU��B�-�E���^,1����@-�:��@{�/<�m��UX^��rN�������{8'�kd��H�9��jy��Oచ��kTO:�=��.+�������>�i���&zL��Kv�u_8�5�v��'+fD��a\��ۍ��%c'Jm���:��*5.�][K ��������.���XYo2�8�鄩�M�i�Ap�[���δ�t��.�)S���Kl
 w���\�Б�� �5*c��){P�:/8Q��j�[�V����Rti0?%�M�$H�R[	��2�1�,�nZ��em"2NA�N:�	cN��c#,$FLk)��[ ��^�^:���8&�e������D孍Q��E�CbR�>�"��C�����ϸ��v�_�q�y�x��ZmFJ��9K���©�������,��DS�/ _Of�IԜ�V��p��)5_��OkrY�i����Ưmpѕx��0�����eބ�.9��X4�s2�{6��ċfZ=lrԥ� �%}�F-�sJ�Q���V�=�Sk¹�g���J����_U��=�p�WK��W��F�������.�"�.$#��'��,�o�_Eq"P�9�8+�����i�k��7n��좸C;�)I�LQ�p(��Z��oq{^,&LSFo ����g��Q;gU��$�G�)[�OQ�@����.��.�Q0���W*"�Ϳj��:��� ��;����T��Xf��ƍ��8�����r	�A����'gm��
���U�W�A�{7�C��?$�Bp0b�������mR�T긂��Q$׭��_��F�wpg�.b=��S��W�������1
Ȧ���\F�k�K�F�b!���+��%���B���*7O�5��Zt��䗲������^���l��:��Z�B�nݪ_�)	���?�X�\q�ʒg߶5�$���Ke���X�:�@�*[��`�&h���u���Wje�r�Bp�q+Z -@�C��w�Ȱ P����(�u{Up�[yB�<�����ᣧb�N25���p:����\��:B���J�����z$ |��/ ��_�c0��w�D�&"�+ՠF���z�t�u_��N��T�X�2�c�n�e;&d$�@Wu,v�x�j�b��l��9o9�jZD�u4|��X��JJ{��'�Q�]���kۮBK@Å ��K�@��쨶ǜ~u����,�k+��~c|�ρ(bRK���Q,��V��M	]�+�k�SB�T��z/�~w�Cm�pc��]`�'MI��;��=q������>��t�R��"o �����5��{�bg[�����͚=u��j;���*j��0�A!?��U��f��*�"*Ad4����fh�^�D�G�o���d�o��֌��{�9Fc��U�B� {�¦���TF�WΛ�;D�I���!Y5֖���֔�F��w��n$t=<�TS$0{�k%1Y��B4)5��M�JD�5Nn�Jhd'�S;����1T�~�����q�MK �Q��f$��g�7�-5��p�%y29��Z}�nD�K�$�8��
�.p���ry��'*�'�
�6QOP�"hQE�3!=��_7��ޙ
��u�gC}�r)����w��X+''��p�R�e��R^��Gp��rk.Wl�"�V%����x�д���c�;��xr�����#�L�� ����8$g�]�:d<"Z;&���zj�����7���`��jH�.���|4L1���pMB0*0gr���7	�c��J�Yns�Il��xd�yIo��a���j�S���R2���9��[���#Q�'�-1.AJ;�.,f�3�k�I������p�	/p���5P��#=�u�T#&<����~OwUB���{I^��Rc�u14;�+�j�5���߾yB�������O���"򋧙\��xE�pԟlLD�nW|5��+n���սވ��Ep��Z#y[��X�D��Z��+U.̩�aXX�hO��� \Qu1}G+��s���4ք�n���I���*j �����!�O�2��ˢ`����#�L��v%�ϛ��R;cc�l3 ���8L!s�J���uU���R���awD4�v���ۣ�Rϼ)�C� �25A���pz�M�,?l7�h��ӛ��A��O]��g�Je����\S=Q�t=�P��L�Y�V
�S�DY����8�T�R[4+�H�&|����G��W�,�ط���C�:���GB֏ƕK�p`I�����*� �����t+�8�$<o��7E}f5"L�u�cs:��SZ���/����[��@_J���'��V���aV�|�z���C�3�b{P����/UP�RNK�=�#��`h;
{�0.�w帛c���9R3UI�Ѓ��8�\�A�kPb�IF��yo�N��h�%��V�[SU�[��qtdO"�ǲL��XM�) k�����?���B�i6�.K���B�17zC�n�n�'ָ�(���J;�o)W�Ɵ�����zE��\٦�S�A�kG���������C�u�^���$:�Dʴϥ�س�p����% ����_�O���o��C6�o�䖂0�a���$����֚4ն{-�@o����_
NY����C�4G���D�㚰Q`�O�)�	��2J�B�����5�?{�V��w��ҝ���`�O.��KɄ��(��f��KIp��ܾA�.�Cd���R���O���ӛԅw����#�����2i1����"]?,m�k���E7x�dj���Cyv���F�jS�E����R\>�(�(�0;`�><���G��w��B�x�e�� �.��/6Po����i�E�x��ʩ+0�,ć$������!XS<����/��d�Q.�)�mw��.Wm��8�P<�X�2H����>f�h<A^4�@��lC/�d.kە�J��V�L�4j��4�br�z�eT�M7^��p.Rwo�9�}q�����fz�7�j����%̜HYI�.��7f��2��n��Gz��Hs	�ym���ۮ����jpgC��m��� xz� B��s {�v|ԋ���PZ��o����#\�}r~��,P�K�>�wڧ �d�W�N�~f�O�#�GQ��5>".O���6lZVz����-vA�������3q�Dw?�$�9�b�<N�S��'7�c�S�!�H���]o���(y�����U5*{w�83I��������d���in�"�n#�~��9��ԇ��N�!rU{�΄=����y|d���1���f18�P$�j'w���W�~���j��;{|�O�r���{{�i�eE'q1@|�V�!V;&�����y4ٯ�uo�V�����A61�TקUG��'��d�]������{���&]��٬_�=��6���Q�k~���'�n��	�h?b�3ί�{��9+"�I(���/��V��� f�Mn�*Ro�%�3➬:rH��w������o%�#�+���+�-�� "/�Ȇ��'�/�!2i��u����k��"�3#��)�#����⎲' ����.\�n,,�vK����հ�91�	$[ÿ�Vw�~��K�Ġ ��Fk;x:�lK]�����uNFje�n4h=�V�G��X%�W����3Oc?�!á��DJ�Cq�����I)�0A"b�L�ٌNqD���8� $��N�%_a�sØ�@&c)���Z�I	�'"�㤛�ۏO�WƁ�I���D-���_z�2�Ɉ�۞{,k�߄i�׿���E��#������>��wҹ�˿^���-&�X�Z/�켿�;m� e� ڃju�5�$7��E�N��;�̽_�m������#}rU,��鋀�#�k�F����b�%��
��>J �2���F����[1�I R��
V 2�(���y�`�<^�m1�-���w�	8�������sI����.��i����V�-G�p�4bzt��M:�����I:��;c�
@#�&]@���s�5(���;�n��N���̂���z��N�C�I���D+��˧y�P�����2`d��FwB��B3����Z�ӻoz�,>�'��+3٤# ��Hu19F���?~_l�(�i;Z��@�:��� �$���N�E��5�X>J�!Q"(f�̈=�Baʀ��Qk�����~���=-����k�fr�ע�d��0mņ�V[�w�)ֲ�i ��*2�M�U�	�������K������@5�y�(���MKɼuת�4` )���b9�1Ke��0�V9sۃ�~�UGm4�s�	~�4D0\� 5��+>��X��P��Oy����HjܽBlr*~[��847 
?1H��Y��\馷�t���I�b�z��q��+A<`wu���#�7��:9��7K��Oۘ�P5�"�ߺK<�q)�e�Юd�.I��q8@�6���: �=|�JaR9��ɺ��ψ�T���GG�1��@ 5Vx1Ha�n���vFȀ�d5����gV�5?��Mv!o�D�9�b����7���HwM�N�aB�p�m��+m)�65	�i%8���3�|�$��	w� Ĝ1΅���hؗ�
q�T9L[��G���	���N(Y�����C��t
���
�������-�el���,�Eka�fa#J�݀w�ʁbv�y��+���[6�}:��"Bv'<�8��j�1Z�*O�[V��:����ߌ7G3��B���KFa=�L-v��+X�=跟��L��i��$ �T��YA���1t<�Co�-}���z\�&�9_��ެ"��(�$2R��R��˫�	��\s+�����Ø,�A�q�e:��~}C���Y����N�S��{��'���r�ɾ�go�?'�(#d�t3��7�&׮=�ˀ�-_��g�e�tU�)�}�EЈ��H',� k�lHdඝ�9���x�)�v8P��W��bJ����x�������_��p5��*��W�@'�J���
PQ�����f_�Us�\A�m�B_b*�T�%N�Cq�m�ޛ�z-x!��al�02�a ����g�f�;^��f(���I0A�tJ�cJ��mO7DMM<Oe6�Kh�㍼NR-�}`����'a�yک۲N[��P�c��c(�30z��k+:�2O��[߉6��HH�6�p�ܙ)l�o��k���J����ض	Kn7	�Mq��<�xEO��_4�4���g�	�m{G)����}@�z$+��s�Ym����+�lL-���Hǉ�b���I��6Iu*��
�R�R����Y�A�wk��U#;4l��d��∔z�-A�Y˺}��\P(��J	@�q#Uͪ�ě�N!6vj<�J&+[�N^aT��ua3��x�54C`2/�NLO�਍
��6�,���v[$����'�&��vN����樄؈)��"��O��*U�5
x�����Nr�&�< �5�ݭ2��jy[��A{����>N^��+ڶg|��Ȱ������~M:>�j���me�wWW#���ήY��'Zh[�'K=h{Hi:vp�K�/;|�.�ڀD����?Ti�y."�(�-Dhiќ��X��"{8��*%��0۪����ɩ�א��K��.�Sº�.n�"��P��6 \	]�8,�����Zu�,��@[e!?�5]�N��+�&���u��؞�^gb�c�,X��#P�_Enb���xX
�H>�i����P�����w���7�2�$�Q&��\~��_!<@K���s���KbZ�n}��l?�H���#l���J�c�PÖ%��A��H��w0>g/m�v���h���!������1�G��!x7g��,��e����ӫ�,�A�%|�� ������~����Ԭ9�`�ڗ��y�N��F���eP�g/r�������[���dScq���eewn�f�4:�T������0�ch��tC�yR�sdl���m�n���ٛh ��������j��,B�Ю5С��^)�N��ء��B:N��
ec�-�Z}�qz�kk�;!��~�poA��rt��zEf�1VD�^n�th�'�/Vx��{.�w�TE�+f�E���㊪��_�i�f��݄Ʉ�<��//
�����oZ�Q�,7�)L#l^�c
��_>��!�k���MM��F��MΟ�6C8$�r �q#v"���" �F�&�]�OE��������<5�y���#Q.�;�Qӏh�T�[Poy��ݵ����Ưl��Uޟ�v�a㕶��g)�Xo{V4J��X?��VLD�G�Ŀ)�`z���ZF��� ��Y����4d1CO��d�WuI���a(�#�;A�g6�8��L�3�y!���I+os)�����
�S�6B�x�t����,�<��ē��V�� ~ޡV����F�F�"��L��&�j���w��	ۅ�.�'u�H�3瞩��'k�݃�+�6f��wݭ�y��9=�q�"�B��dRa��������S��C����R���p��'�<���26����?��/�Ҳ5�T���dƮ�ňF{�s�w���DWH�y���ך(`�{��u�L#/��/�qC�`���{����RF13���6��ձpn��L^���I"�3�7@Kk4�_umڷc��_�+Q�=�[o��]�A�����z��3 MR�y��|y�ï�|Գ�˫5����©p w�&E[XV�l�j�(����I��At��Xz}_'5���34H??[�~	��H����d�ٕª�T��[:�,3w�oysg�f/*Q�'�*ǾK�����xV�%�l�Qlĳky1Ȁ�'_͓<ݸ]�s����J�?�-��mq�r���r��Eb<�7*!��¨�ѯ2��w���C�EYM�Ú��Q�Y�JTrCB&��?Uɪ��1���e�|Α�z�ji�Ϳ�a$k� �u�jV�46�N���S �s-�qˑ<Ci�[�,�,:�E�b��1�RA�M��9
Tvo;��E���[�ck}Q�m���f�*�S�At�ev�jIP� ͟����!�ڍ:�S<�>?�C@���SWoFT��zl�9oA$�L��|�ۥ��LA�(`��pގx	����vt���&�1�l�P��qb�G�K�6�������<�Y>2�pZ�R��Dy��u�6��ԁ�l�!5��Q^��U?�7Ul��bz@Y1Q�^��?�$�'���3������\*^?.�p���Z���r��u��\��%�Vg�jYg1ML\�w �� I���r\���a�>@����Ƈ�e���������P�?�sH�Kx�����͕�����!���d|��F%��k�-�y�<��/`�D�-Ϝ�BNHQ��S �u����DN,`b5�h"�_�|j�*F>-�C�Q#}Pl������R�]Ot/G=w�E��vL���k@k f�_s��Z��?Tw�h]Ћi��-�f��\4���@�1�����1�@�m�LY�쐑���ŷ��G�)U>��5�Ƨ�����Q!s�CQ¸�>���WOҬ�m��)IIZ��"P<M�s]�:j?z�I&	�I��45��'�<K���,E"qU�,�G�d!R+V@�q�f.:Ĵ�G�'ضaʚ|��u�o�`ҥ����[�rq����`>,u�`Q����1M�Q���ΰ��y��8fP�js���i1V�St_�7����Rtf#{p���:H3g������Ynmw+�'�к�vBx=n�e