��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��@���_���2�pۻ���i7�b�D���V�𹈙�v��#nv;���v�N�ͦH>�E�/G��KI��
�n��Io�i�;BlS�`ar�^x�ͼ�ZB��˶��9���q�mE{��1�!�$a÷N���Q>���;�
�����P�6qG��A���W���(��C��ˇ���Ú�@����ޫ�T*����*S�p��G&��"p*6�'�����d8�5�^�;z���d�[^��Wd1�!̖��y�&�
ThC)�o�&��]��v�B�(��^=��0���y��V��{'�c��J�b�%M���Mb�Q�"��j�#3U�$��+Nc+GW�ʰ���S��o&[:�����#	ڍ�.��cu`�">�1��7�����2���K�3ǃ�~&'4QHW�����-���a� BWw*~��C��)�a��Ăʈ�;|Q���ݴȲ����}����c"�vwa�.G���ջ�6�-;p��<tu2�����p��@�x�E���~��D���_em�N�O�x9�(hS�N��tKr�}٬����;ͣ��WC��wp��-:s��2�
;y�)�Z2����AjX���Z��kѣ񪃖�t�_���{\�V�xv�:��Q&�ŋS w���Z ��6/?<�l�sI�Ee2��f����ǟ3�5X��q�����Ӧ#k�*5�kɇ�o=�ݺ���|6�qf�
0�@����ޚ��na�-�aU��������]�m7��]~kQ����Osh��(�9��R�ln�v�{V�g�{���H:!�d�����p¥���*��
't�@��Ф՝����;}��{�u�fN�'�LZ"�i���4���9�׋��5BU�}։�Y'z`9`�J�I����F�}v[|Q�O\`����ƚB��Tc��� N�1w>��[L
aó�M���Roj5�U��2�}���O@6�?� �G���eh�������c��6��@�r?�1{<�V�u�����Q�CCY(�g�����mi7��
�N�[��R�
���@��Ż�(�:��� fP�!$�B�.Y3�����,������r�ٲ�!���N官�-NfK���Q49��ۘT���%��l�v��q��A'}6͖;문�6̵P;cN�����oHC��,Mh�Z&]��_��?&.�r�YAE� U�SQ�S��K����`�F�E����VM��f�r!�84&j�,N?@�Ι�c�p�1ST����P_b!WS�o+D����hlp����ȃU�X�7���	(��b�ņ4�~e8YӮ���� qCݜF��V�Y��$���gi����O&�I���B��^�p�;t��^�6+FV���?`ۣ���CA�W�ǟ��/m���ǠWc=_W�9zE�Z�M�e���