��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���KN����[��Z��*�T�Dr��[F<D�z`��D]Ñ4���ۘ Z�����h9Ľ�%��(�[�%���8�m��Nh&��sO��8���8x�߲�X�6_݂41�CƩ��r8��N2�k �	�� �������S\�{����2��e%Ji�U�6C⥟s��Iɣ/j�Nޟ1ou�J,.�����!�8fw��bF��������&�9@~8mAߌ��Q6(Ϙ�!E���l���]2����=TK���	[6�����06g�cx��
���Ľ[b�c��t�"���`�A��t��2+p�/Py�+@@*i�A<qi�}%I��$5�Տ�
�D,X��+޲��?�h��Ւt�ډ��L<��X"o�܂��Qa��G�I��t3 ����$Ic��Q�r�?l��W��n�4:���Jo���u �۫ ���� �f��ǚ�ne��!�m~�5���rW���h)��=2m6�+fY�%��ܛ_c��{�ۅ�yU�߸�Ңf��0K�4@L���S*{� 'G���=�Ou�G�kzR�X�/6�H]�9��_�8�_�iU�����&v.H�*Z�v�z��b����?��ë)��%�Q�C�I�/�Qv�0JV6j �{��::e�.�7���#��J[[2k�����[E��%T�7��pk4N;Ufí��m?�I�E�:�"����|0K��3�hC���S��m��ݢ. Z81����$���ܸ��	��TJ�� Zt�(Hu��V���h)����� �5;%�G�t�u�OZ��}�����Z�G*y���ό3 ���I�.l^��g����[7�3���_޹�#���Ė�v8a��h��N�k<Q�N{{`��P��|rY��k��:*&�N�6��~�
�r�]��ck��r��i���1�0��1>�KQ�.�1�N����zҙ�P�φ�}K�������`6����|�b�;"��cӒ�\a��ZѾv��>Ԇס�+j!��kc�΁��pȯط{��Fr��@y#:8ϙ�� ��.�Y�bXX'��)�ܔ�za�f�k�J�����}��Գg�x�v�Q�Y�P:h |��w���|ExM~��I�A��d���@.%X�[��^~ٜu��7���d>�9�h�B{��]��vt���\�i@�+˩�4�����"W�dcv�����G��B�_�)�RU�6��۝d�ŋ�_#7���;ʬ2�s�����IAF�"����6 ��p4�W��w�wz�q{T���&�>��0�6��m`g�Eudh��Xr9`���i2�Ă�X�c�d\�:�tc�T��0gU�m =a�����|�!xO�by�W-7EXd���XY��<�e��~���iF	���"�8M�ܼ�hb������?�KH���U�J}ɇ�a_�ح�X���F��4z.��Zn��~�o<�#�p��:��в��M����{�S���2�g�c7��;9����
��C�T���vY�iWy5^l��5�g�U�����7^���gIV�+e���g���o8�2�RI0�)��y�Q
�=0f�!�Plt�F��ާ�
~#�s�Ahw�H�Ё-�� ��2`�93�9�jV���x����f��T�I
�$��O!������@@3������<1�y<���x1�}�9�x���������%����p��0���R��P�e' @��Mm�G�kL�;)�Y��D������Yʁ��/kќ���)+�k�W�l3ꕮ�h��א��b�i�#�D|}NZճ��fA��}]Z��T�t1
Q�E��E���%�t�Bʸ2a�qB���;&^иO$����`��C[�;Bt�| ^�9��=��B�f>8���68*��~�Ɍ��fi�ɢz� l�7%/�sc�`w/�e���w���8#�H�&��c�X�.B�Fqc�� N��:?:�(��t��	�j�d��$���K�f�����Q�!�|�͹��1{�'ܛ�&�����&4�oi�
\�>��Ü���ڴ�{�Ȍ���J���Q�5g\�ʥD�dݻ_u%�L�
gW���F/+7�i�nR��l�A���ϸ5��N�3�W,Ÿ�����������B�~k��jMN%韱�1�-z|� ��ͮ���SЊ��0�:�!��ƏH0��zș�tm9
���X���j��A<W�R��9�=���[0n��'uc�����Ă��1�2�S:X%�iߓ1�����ENU��2䝂��]}��w.��L�����+��������r�7J�9����6�︾~,�>ܸ�4 �A��<�y�%��d�7�M �џ|&\cb������9!4-������<eI/��d����-Y�Lݜ�4���d��_>��8nd���[�9ep\^:jw#�GgQ	*�«�g�3�L[!�b�\��!�1n� 	��F4�Ϧ��l��R�!BX����M?QjZ�h�g5�3�V�\�2������E��,W����O�p�9&��(/1\�8}<7x�*�$�<�S�4�۸q|CG-"o ���iP#��������#���@�J�Β�@��g4�D����b"��g�Wܔ�<੬�\7��:寀�t��g�!��e��K眹q�]l����~fJ:���p:�.�h�kD�����aB�v��7��܃�4�@���){�atm��.���o�q��dp������v8Q���
� ���ZC>�y�S�YwMW�Ã���"\����S3�A��d&�<E~P�fh�We����S����L�c5f%��W��=v~�����_ť1�� ���1����$�!\�D���P��_RM}��p>���`�����刮r	�c�\{����s+TsD�Xz0�~��7��8�퍌U�+�;��
g^��������w�IP���=�*p��@����=�zc�<�{��[\s��~��㬺��'�Y�hɛ�Υ샋mE�q����37��\�j�%q*?�a����i���l23,uw~�3;5=,�w��H�z6��n�5����p�2C��Z����_��_��-����9����5�9ĸ_|�wP��4�&��OZ)���l��>p�b�y�E��D(0l)�N++�H�܋�y3�R�ou}Z�7�q>>I��,D�S���%�І°u#�H���PyO�2h�(֫�=]d����ש��n4-�[���e����O�W!�Ѓ<��kY� �Ѿ������}�)aE$ʗ�v�b�5r�؀!ƯlV]0�i3P�{d.�F�7i�	f�\��o�mExm���=�Cqꔇ���2���@��s�=k�����I\���:�ÀGM�$��׹�ȧ�Û�4�5�l�y5�MaK?���;���C�^�f����C��
Pa	҃��(�?�YV����i(	�?�<��#���3��X���آ�v79k��(��5�{ՙ��?b�*�?���T�����=AR)�u�o�##1�H[Bi+�ꯌvⶋn�9*r
ҙ��b�PA�{��F�fCb)�rF a���\,�#5]V���\!k�t#ڎM��
߿ɽS�.�`̷�_������Z m���~H��i�o�֡�����%�Ax����C��X�P�zC�� �R�va �۳��ř��#��a%9-?�&�L?�@�t���ܜ�t�P6dp
�]�հ]����8貶C�S�yEokf�	�x�Q�uE�.�y^�rI�9���6d�ޭ��c��-�8&�G�;Σ_j/s�	��K��|i��>����W(r��}L Q����3n
����3��iY��=�-��F�@R��K����E)��c���ª�l�Rq�ùm�}	�����/�IE]�x��?����X�1 #E�~-��h�׶;Dbi��HZ�?nay�:�E�YќP~o�CQD3�$�R��Tav�:������[ H�%C�n�����\7�Q��[��{wD�/R�!<jGs�/�=%�K�h�y���F���nz�����G�͎aҗ@���4Xe��rt��>���k%��*��Y���,ϊ�o
;e*_�Q�Clb���/?��I2'p��AAcIGy6�����/'F,=����1��M~�9�HyV������8�~7�{|����!�/��a� MF0�d��R��r4%����������z����dA���Sz#ȰM�>2t�ܩ�NH;F�ֿ_�.�n����c)�or���*�`�*{��������R=���O�Ţ�͵�<�uV�#n���R ��3�<W܂�g ��ᓸp��/4�����>*9s�㡻���i	R��FY����!��j���`�ˌT�zyp<+H1#����SB��;���h�Y���ms�;~��W&�U��m��-T��܅蹀��n2%Gnc�sk��y�ft~:�.�G����XH�/;`f�B�EE�����X*j�Kk_�Ʀ�ٕ<\��F���^���<T�)�/�:��Y��ۑʯ�?k<]��Ei�����oM޼/�Slr�/���=+u�V��:ؑ�(7i�����K��~�&�A�4@8f~�!�d()��r?pJ>��ʮ��t�G�GE D�o�T*���8q�����袂q�?E�a�,l/��qJ�O@o��h�.$=���G{{�q\d����{��=G�*�L��Un%�����0jD�֍��ln�PDW�����C�"�kV�5�H�զD�̓a�(۠�o�EGnt��Ӟm��;���UjL�� �Ժ���A�L%���h0� ݒ�u%���U��[�$�k\QN������q����D�oqa8�qc�WX�n�H1������Oc�����`����O�2O,nj��yM:FdU�#b���p�v3��F��׍1�d�eF��A�F)|��� ��oxK�Pg��Be`�y�.�QRj����$~|x����s��V~8�x'N|���Gu@b����ly?Б"PeR����`Es�ܠ�h���A�y�MqJ�UoL�0��b�N��xW�'1�Ko�/r�e[�9�I�,�=���7����.�~:6
fj 	���"���)��7��&tON�Ƅ�Dx\&Rfi��m�����sf���h(����j�S� YÀ'�9�oO/�^��;�zC�d"��-�Ph�Y�Q��d��l�%�ZL�JԼ�S=�%�/��dy��˂�[RZ�7kfw��O�f�Y�9�C)��������48CZ���
l?1�����M�<���FL�[ ��}G|�{3=n���Jb![�������%�0�jt��:Īk�����'i�(5�X��m��G,}ɿ������D	9���֒���jtO1���-��٬~
z��f�S�qNa��©�I��K Lmd���w�:�WOu��;���>�y�!�r��4.W��/�\6֒�/$�K�M�kUe�v��|�2��j3Z+P�:`n��Sl���Ji'�/(�q.�������!��d�`F�䜫�u��E�T�~B��l��5�WY���A$��t�������E��W�BF뀲-�qr[����,k���o�F���؈�wLex�P�J�^�&��m�U���oa�Sl�u©��Ѕd���ߠ3�\�T���W�/���ӈ|�J�J'���8�����9��+4lr���1|�ͰDR�J�N�9+,1�3��1x}k}��v��<}O��jA���f����ĠͶ����K����vo�����0\,�_`.��:F��ĠY���j|��E�N;{r=M��چz��\0�a�A�n׷�ٙ(���e�ۧ���m|j��թ��BO��Σ�i+���/s���k؆�evT�;Șm�s���*�BQi��4%�V ~{��^����Ξ�E5��k1�҅ի�H�q�v��f �6�\��/���	�k2��js��f����^�u����7w]��J����1��2�-՞���*.ǙV��O�c���A�k1�=%
Ǒ�:�<��_vV�M�G�{���{K3��(8Y���
�a��-�$�Rx�zw_�����k	!9�V�����4:S�w0b8��j�e| b�e5��yj����G���~���8<�����{Y^76��B���F��2;��	�ð��T&�T�_�l�WV�r��ZH�E��2>+�����>�q6�6]���X���d^?��K�t	6-^kZ��:j�/�����D��zv�6���!u#+�1A�q{�k�����|��p� eB[�Kd�b��� >r��Nl�b��g`&Yŋ8���cEO�`y#IX��/�o��������f��)ۄ�����ͱ�ᔨ�=`D���_@��Ppq*hzx�Y������#hf�MG%k��'��b{�l�a��%fzB�j���mO�#�ê~���
�P��޸4H�"X�8O�,� 
��Y��+5��!�����fUV����+%�4�s(�4W��ͼ,7W�
�^Bq�3`�u��dR��X��.�$xHB_���� #���D܇��Ěj]�%��Y��I�� ;j�;�@�VN��c/	��n: A����;)Ӹ�-���;R=�@��6���C�:�ÿ%Lc����+3,<Z;�]$�A����A���ef	�%�u�k5�X�6�c��_dr)��B�R�>WAx�D�e���X��"�'��XRG��_do�Z�_�
����hMk�35�'����yp�,|����s�Ud(���ȋ�<�"$%
�g����/�8E��4H�pÒ>�zW>��p%Q��E�ylQ�Y���kt�w�F�P���`*G'qUY�m7h�[�<���f����7U��.�06u$mDL�(|8��ե��՘B��*1��4�?��j�W"\{�.����D�Y�A�w}�������SB�ҍCcO�wF*�ϗ� 4��#_��ݬ|P9iP�5'3��b޴;�V(G��T�1K�@aG�	�/� ��[̈᫃�nv�Ԭ�+Y$���p�\p�}$A��.���������^��$����ڍى�0����<iu8\_��<{��ԟp�$A=��c]YZ4�q��� �mF[BQ��`k&o�����[Qh��Pq%d�λh�[|�.%k\�U�	
%��>y$��B��Z��(?m�P�JI��{ލ�[��<{��@��z6(I��w;�9��b|)R��ԍs�C����Ą�*�����ZTŧ�=�tG��Db9��D��� R4�,4�9��Y�vLLVѺ7v.����&/$3���ޔpn�������/q�ʼ�:�\^�Y��^�?���Az�u��L
�ꅴ�\`
3��J�&���D.�z���B4{3#����$�B��"Ŷ��Gӓ�(p��b&��zh_���kWs�v&�2DTi��ܫ�R `;c]��tKR��B��}�(�!x�+��7�#Ĉmu�r�4d�1�+S6q�O=p������'8Ӈ圠�$���ǭ�4)�p�`�O��V�<�'ԙ�~f@�U�m�^>)h���qo@�c-甤�/�`v�2e4>̚{B�쫇�G/`X����1�U�s�j�a�'.�$�VoF}R�S�b���a�M8�G��|] k��ʗj!@�n���ȹ�M�)�ֹw���5���#n!��"?�j�.�]݁�M�z�/�F���`��X7����ѢS�''�-ȡȢ�ꋥXĥlEc"�{3��W�e�C[U�oS�
����j�*e�\����|�ˎ�>j��-�oG.��?�4sC�a���:�C��ʺ�c�h�D��˚z%N45�5tsl�̣YSwJ/]������N(o��d�O�9�;�>{w&���Ҳ��/*_oKO��ɭ@-#� ��.�@��*�Y���S�9��tfl5�)���x-z<^���vkx����w	_�'�$dJ3���W����`�����ف�V�K��`�أ����y mz�u��K�ѷ)��}R?f�j�B]�\ߑe�n��:+����=�
S�G�Y&�ݝNl��h�C��������Pf����[.l%��b�������d��N���n��x�![ h^�g��_Q�G��ł���;��$ Ha���'��C�SvzT����J~6��
2#o�:�I�F�(J"	(�yj\ؑX�^1� P����ί�J��}a��V 򍸅.��%o>��&��C��JY7��#�~��)�2Y[teR M�tQcJi���\��d�q�Pi~q�"�E��_s=��~5��E�&`�X7�Z��WWOVqA�;����W�P���"FG�G�t�|ܙ����ʜ�ק���o7�"RZF_���l:ƴ�̋�}�$O���+����Y>vV6�HgU���7mZ�� h3�nK�U�w[�[2ٚ�R/m~���Ċ`����Az�3��>�À�/���u�B���YL.��.��Z�8��P�����Hې�q�8�-�|����\k��,g��9�����M���|+�6b����5|>�V��'
�J�q�r���٫�ܗ�&�v��x���@�F�c6�L��)�e���l��)����`Ab��l�$���4�a���ˮ_�*����#bd��{8wMg� )��a����f�/�Ď:�R���Ո���<���Q%\���"�7�����U�'��%/L��n�?�Ev�����{�:+͡�0��!��G��U�d��}��qRuVi�0�C�u��;��:�~�.�Z����oX�x�y*��[KC+Asa���D��XV�������:����ۮ������<2Q��Yk����nɍ�Z��6�����#�&�Ԭ��	@������B��k���h�ޘ�{4��a2�!���G5c���������j(�y�Z�إ��}d���6�+��Hv���aI���^�[�����	��Y׫�a���ku�����-�����t�f�\���i�huLa���|:iH�z��;Or1Z:6�<���ث���=����	F
���%S�������;Y~[A�Px�R�� {�Y��▙�~�����_�˫�U��[�Y���R��߂�!=�BuQ�������af`�	+?�����k^�Pk��L�D�q�/�"�cyX)mQ��a��m��nKl;��#X ߱�=_	�V�Eík�����m؞�$�ܫ���	7)���i̝�|�u��㰔��E�\uu��I;�TA���џK��5�@L��-��L�xXǧԼ�D{��ǉ7�ҡΠm^��(�2o�x���eO������h�zy.���-q�;����Y�� �cϙ�Sf���ɀ��uF��x�A������KQr�F��I4�//���x�×n`%���KQ��%�(\����r�xs"g�)���/+�"f������^��G�|�9UA7o���u�����<���>��QX�_�����5U���W�q���4��mXߓP^�̨�&�бA�.�*�dO6"�ū��M	Y�6��c�<E�e��o�$ۖ��� �=�2�m_[yU )��jW*ß8;���ӌ��X�8b�ԩ���G���~K؃���b����K�Hs��i����u%��2�Ǥ�.(�_�q��$���Jy�B�M�3f�~;��hr���T�'�9�!��<��O��9�hm&�x�A?m	�w(kTd���n����sJ�"2
Sd��"��Fx:~��
	�I���������_�C��D����)���d��䏯��zħ�J�E�*>���v��7�@��]I�8�0������:�1�e:ˋ���^r��vU�٥����B��o�T~���%����A ǜ�Z�Q��s!�g3wu�}͐� ���8t��uF�� .1g<�����624�6fl��m�Hs�U�,J�զ3�����'Ӻ+ ����t
+������mX�/#�Q��^sr1��mӤgIO�j�LL&C���x�N���ݣ�t5���-_��$�k\[p����@K<��� Mxx0��������ǰ���;�w����H�"}3�vme�T;ݤ��٭���jnĢ��)�
�S��b���|�V6k�c���sɲ�[�>k������Q��i�z�(��nM��\���t%�"�m���Z&�4�g�SY-P����