��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2㨇VL�X�D��G�9�������y������HiGi�U�
�Td'	o�����~�K��M��6aH:���t�4����=�U���әڐ��Z�}WQ38�gzL~�2�������/��Y�S6=�IZY}�h5	�4��Szͺ�-8�E �mV�q=:!Gױ�f�*���_WP�������_������� �x
���^�lI� �:됖�YFa�+��Uh��T&�����*�j���uq{���i�LWW�fi�lU��خG,�o��?B�����??�����gW`��jp��~ �7���c���g����2@ �~&CA�K�dVD���P��������n?.�a�+��*�/?.����࿰$�K����a�(� ����wڰ2��h璇H��=t~��K�P�֔�N,R!s#ZB�10k��H�D����R�$�Ky�����k�=.�k�K����F]
-H_��ߤ���vʙv�L=XAs�~uu ���n�-�d5��u%��=������Vi8eĈ�Zl{�9O��V�%���XADDy[�!�,98��`d���(�y;4���f�im*��s�0� r��Ս�`����6��p7�ݞ(�=�ψ���_P�T��iB��M@�U�|�^,Sz)��ϭ�YI�"������t3����~Ȼ���dLݢ!F�|[5�.(�62W1�1�Y���W$K�Uݖъf��e�e~R�Z%�B;�8��S�f���=�}�����s����b�⟱�}���7�MIU�Zc� �Do;�����/fh��F�� ݳ��6v1��U\;�g�! ;��i������=U�sPw5�nw�����|	Fy�t4���b�?-���>�C����zL���m�Wmû�� ���ڠ@^!�*���-x�� ]sT1K��aP4Ϣ��-@<�@=d�k��}q����v��,��Dqd�^S�����i�H�]����	��R�"*z�G��M?^��d���Q2�6O	/�>7��A��${U�����V��t�h+�L��,m����_�A��.x"Gkm��T�V-�i��@C�U �F2�Ը1~}�Ap�l^%4a���y'�d�z�	"CG��6Q��ш�l	3#��a҉q�{ ?�%3-�_�	�h<�,[ �y���qa��"���z��2�];�P��(����x2*e\Jy�eZ��?��m���Dn�\@eµq��2�beM��G�*�=�����w	I� f�S�����}�P��o����"����`����\�ʐ
�;���ow��tѪy�^����O��v]?d����Ajd�u&*�U�ܨg�I���O|���������Z�
�p�^H���`�Dj�x��K���I�aߗ�B�l���y�X�|���I)Js�Bz~ ����מ�vkK
�fm9�"�j.U�Ҍ�Q�g?���СT�f��>�b=	\����Z(��XD�|~i�M/S9��;MD"9	�7l5��1�&�9��W�,F.�I��!���?s'S�����goW{QF������?2�m1�g<ee�c�uu޿�z+4_�JV���p�S�N�����C��#i_�8���@����1ޗ�Ҵ������&D��l�����V� \gf<} �W�Ү�T;�����>���r�M`f�E�d ��ʌ'w!q�_Qv�m�sb���+$!���N���j�k2�Se(@��ѲeUF��8u��t-H���pXh^����{6���?��j�
�Z�]m�k������U��#O$��TOL�n���T����!�4�3鐗�"��^}��+����k�۫��)��M�Wc���I��7�����D/��8�k�������<:�H�7�3̆� q��ʔ��,�J^�g�4!Y�}��HH����x-6���GО�h�08օ%=�������6��|	��rk������ږ%ŏ{�fR�ܝ9����@y��Rrw�I�й��3�C
�����(/�2��'��g���3����U�	؀���ǀ��'������xs*�Cr�c�M/'��=�Bx�������I��rd[-V~^oB�(������v�Y��Ņj�44'Zu�z�R�} \�� ��e�tS4xٕ�"n����Lm<DE.?�7?r��Ԭ8
�]c���Қ�x��Dϳ�L��[q��}��l,Z& ��Ǿ03��S5߃q���f��q�5Zj�25�ՀWU_t ��R|IK�VÐO3g��XڤSx s�������0\�UWx|Yɸi��5�ox}���w
o?�(]z�U�슖"������M��i%%]�eAe��Ьz���*[��������B>_�c3`yN�O�d�r~A��w��CAj�����4�$�Xs��t�w��O`��1v �&�OZ7/����L���+��K��$_i=���M��Wefl��o	)AY��;$g�]�u�ۀ����f���v+0Ȩ��[oܾ�-W�����$b��Q��=�ѧ�a>���_�Gz�N@�Z�Fy��g�����_��o2�~���[(`-��vT��ˎM���"��0���&BXd�zsE/P�S�5��>�a�"xhV�X�@ϐ���x�J�Y�]��UGd��Rc����$<UAp�knwW_�;m�=��GO-$�*
!���{��V,���Q�:�������Mm�8�@�����~����f�\ww.�J��S���W�cD�t	t��biٙ��b��L�E
��0�;��?�ka5��J�`p-;Ͽ%u6ܑ�"BC{Rr����@p�������Gmc�������t�y�6����_��b�u��"��U?Լ�T}m��m9��h�a5�OB���EW��t��q��ZD�_w�r�d�e��[�Ց� � ��D��nZ3<x�t�{	%�w�&�y?vG�/і2������h���S,�Q6k�`T��}��G�yZ*�2;��M�z*�/��AJ�RR�����R�k��,��nq�<J$J��I;QU��~�|T5<ڇ��o֢x 89�싇d�8�ډ6}0w���54 * ����d������f��J��E.Hk@ȫ�[d�D����^>����֋y�/�T�nN�u�����B�6kVI�����o1$��4ì���_�K���LA\._��q��O��o�bK�ւ����j�S��d�I�	�{$�[u=���L6_m�Q��ּUR�l�8� ���y�:#%����Irh�D\�\-_��4�����ϧ/p�n��ld�(�ˆW�Gے'����[#�cɠ�0��k�s�ɺ�K��4Y�|��=�x9����(�����5��IDf2�xp���i�R��S��37v_h*;B�a"�4�#N��I`
}�OG��Y��w�93~Md�غ��z���F�F5�%S�sUAl�U��x<�V���`���.;���}���Լ���,�E���@R�[)�h�آ�w��Z��	Q���"��fd�lB��J���DА\�D'������:��;8��{��%���n���t�0��q�{�����Gڜ���Gư���
.�����^�r��q���2���_����N}��m��V��\S����hм��n��%�������( �r��D�G�����e����q��~��T�(�ڟ��c:ݰ*Ɣ7�0�'�OjK{�Ԙ�˂�6b�]+����E��͙&#�Z��wt�t4�>��D�n�s��SfQD �F�g��[%)Nb��-�����d��7��L�?�w,D��N+����u�t�,,����Y�  V@G���M�݃p�A.�,����P���=��xi�G`�� �p�?���o��{�����+L��(лy��@�W�_���J��d����Pd�kbI0FV�'�h���)�s�T�K�uc�	Oޏ
֎Ѫ#2Ꚉ�6���;U��b8�~ �%k��!�>�#�ltrS
��}�rM��:�k�5��b��m�K��!%�Y�T����ws�h�9�W|�gl�m�8V~9���˨�E�>�Ѱ�V#k��=����H�|g����Q���q�-��J�uyJ�+��q��Z+�P(f-fŎ��š����d�C�v�Zo(���.L&d�*Ӛ�EW>5�22�:˷fWR~�{�֓�E�v[CCȶ/jN�����E�Ѐ`�\��:�CP,n~�-11�G�"' �%p�����q!B8~_n�1GQ"ɮ�!�pI���������H��u�M������c��s~����D��gr`\T�2��jb���^ġ�,���n��t��*�n�+��u�6�M�� ^<ney��.\�� �ϩs�'��_��I�0KV(����k�"�f�c�m�[�0{�S^�lO?��20B�[O��~o$������3��r�����J����@.����c��+QC)�V�4���R���cȃ�ӊ�}E>T�s�=u40�e���.�1I��$>h@p�B����G�gPz�Mѷ�ׁV����ߨ�^�l�Z�@\v�8����WҌ~��IѲ���PD:��%h|VO��d��"������u��h�΁�E��])�ylY�4�񪺀��ꊾ�·�a���cH� ��_���/�ѿ�^���c>��S�&�D�\s����JB��$���ʟk�x�=?3�⬾o=^|�� <��s�Xy�{���^��JB�z(���)�P��$��Љ��K�뻑�oI�Iԣ��NA#X��u�?�\k�=�IV~W�[�d|�WL�������;�Lo�9K~�H�3@����}j{j�#��"�N(��FQ0g��x��k����S��e3�~LfC(��5
��/��ٯ��zs�W��v���/H�p��X��Y��ù�iY�� Z�V?�����v��)P�Ӹ�YS"Ğ��]�f��l�֨�ƕ�r~�S���M�F0��X�����M�����H��W��	h�kЎOh=�@ #�s\^(�<�/K$�xМ���5�B>CZ�4��/���c�9������p���\I��i[����T��E�����St/U�8�^v�tW��Qǲ�+�e!U�GV�Vm�*K��	AsE࢘��Qw�L�E̎��N{C����S�>�6��C�67ye~XY_���Vq��I6�G�/��+S�i+:ujZ'��2�K�]��!�X���R�����h�y��(�zN��� ݛ��3y�B�/�`h��������l5������P��h��zΡ�����>��������w�锍���7�I�&49 u�ƣ�����g�叙 �<�	pS���@_���mkT �B-�Q��X��Y0f@&�dr�ޫ�1�C~�Ш`@�*rϝV0t��j���X��ڵ�35�&��.��>ͷ)�y.�:pMX�?�7�;���/2b,8�E��u�kg����m�h�b����5I�,�+V�00�̣cE�E ~�5�y|܋6R�G�m�g��bnB��(J5 bo1Vvh��y��nsP�\T(���!�|��콓	�&��1k@N����'t�87��8r ��rs[��"[�x+���t֖ Ne�-[�}њ0O|��&o΋7*b��I��0je}F���髇{�����>UsMl��"�[�4>�5)�0�肥�Ar�JQ�X�d|a�$�q�`�u�G K��;�+n+n�Y9ܳm3^�ڦ��U���k@�8җ�)��|��ȃ������6@���8>;pF��2��	�'j�)=�x$>���I����{����w�{� ��H����.I�P�L�ʍ�*;����ݖ�����MBW��<��ZZ��Ȟ�3���{"?�-�s�n���J����J�P{�~���`��T���G�N�e���[J8U+��G�f��e�Cq�aK!��k�#�Fx�~�s�f��ӌ��G�_�Rx����-�wT����U�73\�=~ԍ���a�: ;=;�7�L�d����:k�h�þn�i���Duby�y����C�qQ&I䚜7<|u�XOیN~6��P��;���q�@��!�|Jd;�r"C��`s���m7W���k��;��}b�3�a���[���֕+���Ռ��9���r9r�