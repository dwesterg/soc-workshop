��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,��}�$3p�������?^�n�~��:�ܘ�f8-K-R<�L��U�k�U�'\
��-@��LX��="��_X�`��B\Y`�y'2���S����nu4w�ip��k�\����`�1o���·��k��%����n�����P7� ���*�w�����!�d����.�	 h����4
U��[����m{���~�U����}�(�nQ��+���gֻa �Q�܂�J)�0����|�EﮫJ��i��w?%�ub�Ȧ=����U�kZ��3>e.��:�� ���TzR��S�6XZClLAL��m�*0ER����@-VS�gL%���2�Y'{�_i�J~�X��LY����G����0����0j=�����?0�K@�F}�7�>h����)×����1Tu?�����J������y鶈]��Zr��h�*��`t�R��BG ���м"�����N�<��R�qVy�l����gM�гb���eK�v�ܐ ��tf+�.��k�+�EH�mjܽ3��r��q��@��o`��8�IiEE�|	��	��ڧid�G���_�@6>�s~-�jI��Ls�x�p���o�U�`�3�y�PY���I9Uzش�o��|Ҥ�R�y���X ��.I+�2���c&[��{�r��s��]'t�q�NF���eN��	�df��d;��{?�$�Qn8��F�h��%x邼����J�cn� <�u���p��Ӧ�;�Ņ��%�(s�jc}��pOx�dk�o�C~�3��+���xZ�j�Tj������V	�x��v��b�q~�Y�P�PG��^S���1z�l��}m��`z�¹��X�"��r�ۧC}����!]]RљOH=;�&j<�O�r����R��E����რy�}�ˑr�4{�O�J��Է05�w�=#�X����U��N{�������qw�zk�_��xR��x���m\Oy}�l��m���P�n��H�ʠO%e���v/��Q�F3N���ȗq�w��ƕ�$Z��������$���^a�	��m��r�1�WAԗ��9n�����9�i��YuH~n�E�c?/q�u�'E��u͗�f�bΩp�R���J�G^���s��|�~��c������O�σ�1{�ShaZ�2cd�U�|�s���!r'��H�3�6C`��Q4-����L�?�lUJ�֎�G`˫�A��i��^�В�7�oHG����Y�@;oS�����N�i���o�yT�Q�
���r����D���G�Za=Yc���r��������11u�L�� 6S������ 4��T�w#ٿ��6$fI_�|��̶�V{1�n"��F�p��ę&���J{�_E
@��lU�0"��'�VK�S��S�Y��"��_�>##�M��/��pS8=����q{��༜aD���6�ȜwJ��=��ּ|��e��2�]��4