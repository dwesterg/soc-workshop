��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?����#P�S:;;]�f݈kk�l)Җ�e���1�ӝ���N6������d%KBS�ă���ܶ?r�@��]��-z�D��������<�c�70X�/H��"k>Iޣ���������E�I�1Z�p_X��l?�^�nm���<� �htb�hP(�����'�g�-Ԉ��-��|�K�T0Q�� ���b���S���0�1�ȏ�_qq�r7d_��Y�Pg�.>^�C�=jA�>��
�ep���T����KUni�u7�d�2��r��,��Y��
���t���:MY�~E�[��rr"D,�x�j���y�Z>�Y�ݲ��1*��Y>���6Qg(�?�%?�x���pt$�>��o57����F���E{%�z@��Q�6�������u� �Oir�2+�FR�^R��Y����Ic:b]BI�.8z��mE����58�o����.M��9@��<G��ʵ9_e��Tր/�kmz֨�wٗ몾�aO:� �g��.*�	�m����с��c:�O�=ہz�뫪����O����]F�n��]dO����SD�=����F+X�P8=�k�X�)��&�ֺ�W��Z��4�MgL�߰��x`�+��ݾ���`�O�,�j�G�gb/��]�:�x��t�5�oZD���R)]��Y0��{�����}��%8��������b_�����F��C�0��^�� TU"[E- �̖�*�z���ї���?��l�G�Z�N���#NhI��S�AVy���9��v@n�C>,�$�;��E�:~V4�d J�[�SP��c������k��mr���(78�T�+�H�;�qwq�A*w�ΓO�~���%��q�$��qk6Ab����*�Ae�q
λM�]��B.��Ǩ̠�Ŗ�i^����� D30��#�lH�AY�,lz.�-t;�����lQ���Lf$��2��]��38��aI47Ǉ�Zi�)������$�G�+���{�6H����f�{�{�ʊ��A�;�݄���CQ?�J+|qIe�?I���{�⤾�wq��O��T�z�5'*�l��R�0����E�x_Kb7�C���ֆ���9C������b8�@(Od�/?�pN:Ȧo�����	�6����lb���^Pƕ�#��؆�j����}*���:O���co�������|2=+�k���;��/�_L�̠�:����6��^
���s���fDz:g5^�����x¶��>����Fֶ[������uό�b�K�.��)��#�A�sw@5����ā��U2�r�5�͚'�Ul�������{�s���q&�
"��$�֡m�]����;O�>h<)qi�A�����[xSJ�+��%i�_�?����A��YXў�]fv�8�&,�=�v��J�R��pV�)����ܚ;��ZB���e�4Y]I�2o\/��pд��x�(� d�n��m��}UfU�
!�MnB����@3{J}�
�,�0� 2�%��GL�+�H9":�.X%�O_R�+��t��*� }��lmn�!���R���KӺLI���6�	rP��H����)�^F����6��L9>�3b���k��F�p��kL�I�Ab����J=�p��,���R���W�����U�n@\��p��U��U`�Ŀ�?���=J݄��Y�R�+�(N����I���Ku���//����POo�[ዓV^��$��!��t��(��VCҡ�)�;ka@�|Ȼ������9>����Ã�:���B�,i�т�5ĥ6��N���J����Z��%F��o酙�Bb��n��^r����y}@��7n���n
̨P��b7��9���7x�o�qo��@G�e��Ap��atg��[�GN�L�a�T��)�'��bK���Y&�{ZI4�7?MW���'M��Дc���@��_��oI|�J��q��LX9�R�9���wo~$��Ѷ!Fksp����- �#R��I>o#�U@�֍�4L	2���ir�zL��?��[g�[JĐ���l���6u���e���{���sS�]�M�����T���\_F \�4�h�t��U-{�t�;_������4���@P8��dA͔�J 0M��G~��WD8^��	^K��E��JIzz���H�!�qgJT<����>t��yǾ˄$���_eΊ�0-[�n�s��w�n�'�P�e�ak�UU^�l%���М�r��c�����$�1mݯ���<��l��R� ��h��O{����<KU�]&�0����Ҳ��j	�F�7��s>��M�xD�h
#0Z鋖�V}X`|�3U���x>a6�����n]-ڝ��:��#*�m1iF�a�#Q�9W*$S�����Nm@ߴpI���|�.��,�3`	U����!�.��#y����S�~�[�
J�VL�5�ͽ(�ә9�u_>��`�!#�W-�R��+>��4r�~В�P@����W��-A��6�R�b��4�&����WG����=�����G�2���5 �'D �r�Y!�rxr�ț��.�w�W�e�0}d����>����U�Yl�:����5Ne!?���p:*c�I�w~�#�A�<1 F3��rd��i<���?�� a�ҥ�/���y�Ε� +�F�({��enF���$XcT1j���vi���A!�x��c�-��27���J霸&�}������ߊ3�j^��%�^$�(�l�a�ڼ�|���h��2���GL���I>p~��Xͱ�A="�D�_� �i3,z�9���f�҅v������^	~ R�zƾ{�4j�ST[P�����D�u��(,sh����QIc�y|yx���|\���,����T����ȮUԭY|�P����&}m�v�Ͳ?��" ����\�چ�R��)�������<��C\֫J���ϞW"�G�>g&�:��\�mR����|�~\�y2�"��@4��Ξ���Ғ[r��q����w4D�B�Y�K��B9hm[|v� ��7�������k�Gߝ��Q�5�~��k�Er�G�"fW��ƟeCfH�O��7�?]�B�R�M"�>:�D�d��W뿴�����6M2��L�
F�=�f��3_3�k�,�����c�K��'���U�Fi�=6��~���I�LЮא2ץLB�Lף����'kcpV]0��>[e����w���!�U���:<<AQ'��d����s)��Β%���r,�ܒ\\�0�"K	C���;��F�*��g��
x�qD�X �F�����S8�ȱ�顰�Rw��[������@ �?k�@��/��O�;�U��d��Q?!���t�#�\��(�H���~�v	�RSA��X,���R� ]{�����7Y�X�br�Z��LKєwL�P�\�4�I3��}N~-fǝa���3�$�ݦ�oy4j�./;���1t�{}��!1kJ��u�0M��4N�r��亼��a����x숡-2o�Ƶ���͑
��B��<��<5�}�B�0��f�LX�vw(�����������:��ѹ�\Wn��s��¸ V �t*d��`t�����E'���A�!z2K'�ڃ���Ьb���q[k�U+��K��2&d����6d8؄S��5�b��T@%���d@�!���������pG�D�9��#4Ձͷ|�܉:�EuH�|,�v��u�I��'I��צϠ�ٚv��By__��6� $��k�_��;��G=�}T�"��t�%W�D�|��k�4��|GA����l�Nl*ED�o_{�X�,D#����a���_�.����s�!�ȼ�����ם|���(l}^���tҒ�j����4_�\��OVA��9��$~�p�άNu�����s?���� R��"��>d�ePHn?uP�k�9&�w��c��8��{�6	z�ڗ_��*�$"�������b�ֈ8��ʷ6G_/Ս��ߔ�؅i�Rm�;H�q�q�<Ki/��-�TD�{�yD�L��U�ç�,Q����ּ��o�@l�I����N;I�����,"]�epO�i	��F��]��U?0�kcl�qK�9�{�mN,(��T:+�}٥h�3��%y�Ha�p��)-�IQ����'�)#'�wEI
[�¼0��P��#�3(����p�^��2����xG�;OS�>Nʙ�\(S�%e�nh�`���ȟ���o$R* �4��7��N�OHd�閖�4,��S�.c$�eT@�A����є`D���&�ҍ=�y�#g�������/�+T������12
�h��4�z7��,�k0��?'���g�=��~�w�;}\<��iB�Uj�Ef����m���UD����b��%�},2A�5�����7��n�V��-L�%��Έ�Tܣ��rjc�J�s���7�8$|�մ�:�h0�� M�ZR;��u��M�J�E��U�&�9t�N ��Pb���
)u^ݩ	���5� �|2Tg������3CTu�u�*X=\V>�V���6���!��!�[)"�����Ʈ�������[>Z�
m����E�+�QFB��>���}���+��&{ ��`DQb�㏦ش�a�@y	��������.�'�Wu�S��u�W��O�v"/z��ݔ������'T�q�ӗ44��_��U4�yN0�s3��XV�d��c�z�!�|(����������?���NAep2�Ģr��Eǻ��Vu�>���S�//-Mj̺`PFSW�s�'���_��Dݓ �L�oW%,X�g;}%ր���d�-Gm?�G>Ĳ��%	�V4 �$^�o���4���H�&ő�	�3�g<����(��㥁��d�]ZF��[��є*�S(�&nQ�t�R�nh���f>��TM���}��6��0�����iG�'�U�R�#��7˲��c�Ԓ�HF��(C8�&T�F�8|/ y8bnq?�F%xR0�%U�%�oN��߂xT���v��5��^�}���D��?&�g���f�E�5-��ӟ�������e[C�"�n�xI
�b�њo��-�Ӽ��{㤟��h�j�9t�7�����+�7��<�E��DT�ރ�Om�u�f��c�������ҕ��3+�ڈ"kWpY�n&s�h�ً>�8�~e�b��������bH�6XPXJ�;�H��v=���R���C��U�=L�I�&����l��&�+�}�N��Hz���b��i��������)
--�ޖ$��;J�OO������� ��ApBh��$�nK�)ش�9��}ݯ�N�o-J�_o�h��o��bP�ăt�·a�������`?�c���q�`�K�!yl�Bo&]Y|}g�tQm���9.��_�%軲���&UY,�nd0mQy�S�9���b�F�P�A��ΤZ}ܚ�dTo�W�7�(�(�1;��Nh����`>�K C�k;�����RD�Ǧ��b��ҽ�.J��0f���{d)u9�5:��"�I^�S�f��D��bw���4��ՠ�LIG��8�X5^��U8L�y^������&V��,Q3��� a��+V�e�a�qν�O��1Q���.*�VB�W�$5�f�kӈ�������|�3��ѿ�傳��&xm�\���(�����H8�]�?��y�Һ|���$V�#T�$>=l
��֨Ԋ�����N�eUO��
|���Ӯ��΢��x�&2M2V��F�oe�x�\|���O'�^�J!�,N���vx�x�Q�lY.�\@@�cU��r����J͑���}}O?��۶҅o�^��4ݫ<�˖H�yP�Oo��QK�a��&�Do%��L9�w#d��=��z�bOYw��2�ې����JY��>�L�V]yg#��D�����pJ}��w�"P��>��h�x����0�0��a������_)cᣜ��~�~�;�V�r�)�����Z�P�۔�5�!�[Q�r�a������ڇuټ u��C1�)h,A&:�U�j:�xH\���~���#Ud��Lx@��<�1���3->�~��V���X��e�m���f��4^cRR��c�K�vO&VF�x-$�1Li+�FLT�KD���\��w0�v��lw:;���Zznr�O�v�LKڦw�AYnc�Z�gp�V{
��D�ٳ���,�p���8>XPi(��%�L�gtpn�%acH�Y6�l�3杯󘦄Uo��eA}�t�Gݏ�$�Y�G�
���S!����@C�A��W�n�j����;48E
X�-��xsMr��3)mgbh�O�LJJ���22�d�%��b�� aF2����p��:�EX�ヽ:ɭ�q�%S@��J�n�W�uEp��h�l�c�L�?��daYwhZ�z�����k����o�oVM����]��뢣�5���I��fV+�`w���ԅ/���}P#����Ī�{ii�)�t��,����₾�BOχ�E�յ�^�Wi��|v�>�y{&I�C����M$�_�x.���&�j29*f湥�g���_��j�2��^v���JL��ga�R����:�R�!�߅�_��s�m9"���迬�Y�_
�o�4K�JF��#a�"����eV����Kb�V����X�#�t�|��MVՇ�c�6�-��\3L�Xm��彴T��Ŝ����`C �PJ\�1y��C	�[l��U��^�8b�����"-n�sY��ɺ\�N�d�3�OPˇ;����7L��C W��G��fB:z.Y��v5�Y�?��H�X���%+e@I��8?���6���)d۩������AGg��<�v$���c�
�;���{��i�JB�79F����4����JË�@���w���Ÿ�=�">>P�&�鳶�i0��ԇ@V3��Ȉ��LuR��
�KNC��<�3w�n��p�G$+���lȡ�b��${����q����"$ǵmJO5f<Α�@v���u��s57������>3rD��+.�y�ؒ"�Ͷ���\�fz����8o
�b��.F8�i��mC����9�c��n�߱�t���R�Ps9^�2� G]Ֆi����=��\�ŗ��ma����lۡ�=���{$�eߘ6\�0rV���ӣz����<�>�X)�#\h�k�-I<�X�E�4l�Nx�&� �����M���ى�h�/l�)��DPT�P���"���󋣈x dq�O_�v-�Ts����G;9@O5@��+R���&'�T�� ���f<;AMR4�SM�B���摫��]?�2�B�_B�Bu���߀��Hl�\��U~�yGJ��v�Uӟd�R[�9���!��Φ���S�{���ܛ�V�x̬�>�k�D������=��źV�<�zI���1���w�t�Q.�eL:���4!�����[���Ԯ�P�%��:qZ��h��DR�Q���e՝�����h�
:F��6�+l���Ѵ+--�|��Y�
���ҀA JkD����L��bK�BH��iJ'����
1˭�.����"7�Z��A7IR�)�=~��7���[��A&@����� (��a��������;E��~m��^��>�%���Qd�F���nZ���Vݦ��m�L��幋K)�?2��*�i�xe*��T��R�"ץ+V�	�m��)��Z�����g���u�s�c����𥿃a�����
ݠ��E��#��W�m������w۹��tY{�Y�R���q��u-��-�
o�������zj$����j�Zr0�ovߨ����Y��J*h]"R��*`hR�O�>�Nk�\�-֊{ֲ
�	H�T\��c���7��>W��~��<DSa��'6Q���%$�8�k���#J��8N"�EA9�C�����^%H�D����
ʏ� u���?��!q�R.
�S)�SK63_�]O&�~��tDN�2�m����/���3회͟b#��@z����Y�pv9�:�D Vq�Sn/]M@|SI��:Ѐy�����la���vC�$�
��:="2�Z� �J��2�����e��~A^�T!�A|i�����EM���#\��[dS��Hyz�}��ب
�*�L��e���pE��.XD��³JG�f�cȥj�>��C0Tya@�Z�ؔZi�='�A*S֌¨$Lgz�r���é?ņioj�q��}R��b�	��
�~=f�½��'�|�4=�@�q��l<b���� �D����^O�e�a�_@�9�i�Y S�5.��mR�
)K�����eA`�o�{��g�p�wP#�u� �%�::9A�qȫ��"A���Y���-�������(8�w��E����mE{������V�
ٿy�>��U���Y8MN�b|x�-�Y1�w���vR�fC2;q����Ut��o����Ǚ� YOZК�1"����aΐ�S���H�-�����*�������)~�j|�L,_�!D�?=�UC޽B��t�o�i"��ߎ({�i��5fl]$��wo��`��Z�{��@\�dRs��ə����h����`�'�B����7���"��5r+�r<0Є�62
�2�\kP�IG��@���N�;��a��bQx=���+�hj"��j8%d���ҩG/��oN���r�P\����Dރ�@�jn��.=y%d����R?|��H���`���b�HQ0�'ꏪQ�/f�?}��-@�I=CW<�D>����C�C*zĕղ��2o	�e��v��_UO����l}yb��@�Z�A�jl�"S_(�O��5VIIl���(6;�F/�2\zA�B�n����Z�"h ²q�Ԩ�f��R��L�JO������f�~�F���p��ڪ�������x5[�CpI�WdM&�3����d-�Xq-�����|�QT����sj�����mwT�(����t-�F|��J�]ѾRGkdv�Q��w���]ӼY<��^Re�G��)"hBYV:�`Nb���<��~1���%}֭� j�k4��"����V��q���2u�����+�%7ۑ���s�pL"��?�^��P��:t{�h+� ���8J�_bw�����ؼ�n1յ	ҔԮ�����y~2��B�'�B,P�qAS�׃-�V?��Zy`�О���T�°K�'ݤ������pr��Wlް���*g���@�h��F��IMh OAMվ��eCO����WH�2|-���W����%2_�dwr�ߦ3Cm�it�u��{Zd,n�i.���sPCю&�f/�}��z�#�D��ؓ&���Ҭ�p�J\�����F��2b�{EɫZf���|Ú?Ds]�ZUҮ�Ǟ��gr�k��1� ��"\6��0�K�{��\:�r��T�5�r�x�%��T9�����)�ۮ�����%F���5��2C�:�����՞YVE��8�Ǵ��hI"�ܶ�~�t��F���R��l��<Ċ;Ɗ��فӴ`�U�Xт���� �)�!��@s[�Y����j$��!�	m�1�����F�ў�_]�#��f�:q7�D�J����Z��KW�W/����0�
�{�Ķ���>۫;�NH%Oa�u����C�˺q����
K���M���Jʅ��.}�;�u�%6��S4��eT��fD��Q��e.$c�b0]���b��5}�~���z�����Ga|Ui��&�,��/k�X���F���Ӝa	Y�6,�\�b� �du$��ף\�0+H]@��:a��&.�
�'�u��q� %4<s1���ݤ,Rj������>���顺��"������yF2��ߏ8*�`V��7�pN�ÃP�0gō�dv�u�����_�$b;NƩ��n�osxC��hn�H���4��-_��4��١!7S�z�
����^���E.�~�֤�o��Sv�}����h��<�Z&��[���m �g�F�wW�(���H�<nܯ+�̼2mY�Kr"��\β�(��{��k�#�pJ�A*��,��D�ظ<�`��H+�(Z�U����04L8E2����i�T��`�Hj\;;�O� &��\�;�1�f�ChÓ��^�b�{R/Ń���b~�P۠���-C�3�O��+���W2�WRk M����l���\��{��՚H�������k6>Mo���j�s�(4��=u�C}K=��*�L�`���9	�(���X���5�0��9�����.cű��(�'�����0�b��V73�c�'���!��7T:7a��|
����r�nĞ�(��>��b�>�@��C�h*���K��J5ɘ��P�*��pEFl�s�?�.%Q܁��*�:rgf&?���w�bi�)�T����,��d��)�2���Yk�o�FXR,4F�U%g�����+���8J���㷝G}�er3X�[*
��XA��6�8�1tz�`��>��N�H*{2��tMk���o�V������KQ&喇s�q%&��(��ju�:;r�P_�:����>9�0����>s���?c%x�w�1�O�I)Qpm���,�_s$��`��x���z�Η.�L��uys��}���>�|_�ⷪzx4$�;���?+GF-����`\H��������p
N	�X"ݶ�rd�R�+����>�����"j̥W�u�+���r���Q��2tX�����2`&[ܠ�Z��؞k�o�$�3'���̣�\���zL�l�=����j�^��b()s�DN�hG��v��?�"#�̗֋ɱ^��>Qp��0��D�Gl Y����s~)f7��5��4����=*� v,O�K���=�|�siI�Q�Mc@� �s޴�4�T�N�(�T���u�-?�� |��H+���`����[E�'���8T��x~�q���͗(��g�N�t�K�Z.�=i��ɡ�Ud�T�mX��+��ګ��w������|���J,e<�_`��M�e�W��?��i:w���}'��h�y�5��Ю��5;��D��1��zl\O�"ˎX��X�%���L��@����C)��Ҧ�nq��7�2|��v�m�$�jZ	�c������R����j�N"�u԰��?m����c�"�𧊮qT��Y�5��8�do<�M$\��N�X�=iR���7��J���Rcޟ}�(�x�#�I1*�0���$�618I��`:(.6�/��ΡM ��x۝����͏��0̗ug>x��r�\����ws���u�4|)'�)�6QtdHx��܋Ga�j��#"P4���ML�ʴ�>P��� ���Vs��箎|y�-p�������H�Z^���~�]BA���?æ�-2�Lp@D��<Wؕ�����r���������=<���Ekb��ŇѶ�X��*��;�-x��U��Yd�� �� �C/��|�e�<�b/�υUyn���K�7�m�r%	�[khoش4?���d�,����f��3�7#ޕˠ_-j"N�n�
^ϣ���@�܋���~gM��t�U1��3��U�I#��>����jXTʚ�3EFEb>EL���ȶ�����0a�Z�f�}Ҝ�f�5��za>5�p�Ҕ��x�~R�l3g���$�b!"cBS5�x;v�:��s�u@(p�T� ��4���繌~�;�Z.�a���F��N_z��(��a�+��+����Hm\�t6�;���:U��W����ύ���c������XP�D�4ن�?L��[+mE/k�]�~"�~qT��u��1^yҧ���a�s+s���)��+wy�� ��H���>�YᏁp�;g���`�n�<��e�0�{��:{q��%���"�9��>�$�I��-��*Uo�ϼ�X��+y	���c\�V��;����t:M�&gSx��yC���H%�l�nK�'�鬆���n#�AA&�i�It]��A��:ŕiP��\�vA�d�"�6|`ۋ�� �?�ou��Q�$��Y���� ���;�a~LP�����`!9I'#;�/�w������X�J�v7���ʯ��� ���͗��G�3
E) )�d4>G�~��c��M,~"��r(�~?һ�RO#��!g^�MP{,��D�O@�<V�k�SсG�a|Ô%q��j�up����(gX'���%
w�):{x+���� PK�vs��
�!�Vj!�@�FƥO9��:"�6RL�V�C�LݨL�\Im&�h���~���A���� 䃀��БS�d��e~=����ʋ
i��v�'onV�:z��jHӞ��+挼�D�c3��l�:��r~��-��1���T]6�a����B�I�+�ቭO����8q�I�G[�ή,�� �<�I�>���^�1砢�	�WPJ��od���Lg�&�
Kw�����D�G+���]��S�q��l>�p�]Q�I"�I�dh�V�F*�M���H޾�8s;�1������y�:�u��H���5�<����8�>4s��kT�Q��-��=�d� �^�{���?"��+��1*��m�����f;7�����m`}�v٧QH;�2�V\S_\"�%�����l�*�wf�9)�gǢ)ޔ�O�X݌�pRS�< O늱�"�����հC\�,#�S���H�wBbZ��k$���Lue�[������s�|�v|�t�� �6
��$j�nm�n*�+��*iۅ*��o�<sT��k�ڑTTD��W���gb+g�nt��}�;m�|��V�n(L����7.�J֯`�9]ڟ�[|��ߌ�H�`$800u_4��nH[cBO����N��o�M��I�2��}�� ��w6�:Q���BEA��0��\
�N���yh��=�.x-P���:�-wB��P�� .1l$�?{�Gd����J�ed-yp,�ri�wڧ����վ����v>�.'�.%~�"�1���`���n��~�����G�y�81LU�mh�|�1��Q�O��Y6�9dt�D�]:�s(R���C���a�\M���vu��a�ף<��73E9H�ӝ��e���O z�M�����Y����)��h<>��XD���+��;��b�=�-A75���a�29!���֣݉O͐D?q�ڢU�T�:y�Ȧ���v���D��e��@�����d��.y!2���7_^��Pr!C�@�.PM��b���MփXG��Q{Y����４�q��5�)�	�����<�����s�"�Y6!�P�xc��4%s$oX�zQ#�5#)'XC8�U?,�}������P�${�M$*m�J��޲k�W�5�כDc���D�9��z-�-z�S��c��ߩߞ�󋻮.
zG��Y�z��J
K /�An�Z'�F�`���9&V)ׅг5�����e_�aD�)� (iŏ$C���))�R��5��� ���٘b�U�ʏ��V�&�ګA�`�a�0]�BR�8ʙQ,86��	�!:��98"�|�qb��a�U��_��6���Z��t8��Q���C�@'/�)��0)%���=�$s����;NQQ������58ؾ^���w��^��S��%�°X	k+��Ƴ|���b�+�S�Ҩq/6�Zz��0������r�K��>W��T�՞-�1)����$pQ��@-��v|�_����Sm�Nןx���r�|�U�J	m�s�d�즢���F��O�ܛBA1}
�m*mR�0#+|j֕Ţć��
�[z�ȼ�]Kx��
��ԩ�a)~&�l�?G��Y�T��2 z�����n����#�C��������?��_w�k�<�1�k���E7�>X�M��u���~X��t^��U����0�_�f�9��tj�V�d�����B9Ւݘ�џ`;�Nҋ���&R��"k��B<(��qT�RZ<QE4@�z�'FC�?�>.�I=��VyfR� i�͵��atf���#s���4�� Q�A�+������StY=�����"wLv��w4t �y;���"ﾣ+��S�sQ#��x�Q���`S�����nQi̊�gm���ψ�7���c�;�Q�,B��M�]�Z�}���7"�w��=D�'E����i1h-p`N)�Q���D�C #�_-%��=�""�P���R���@]U�I�2}8�^uŌ��2�	�gI�=�)'���1�����$f�a:f�;A�s�':;��݇�E҅=ܧ
$�i9R�43����.��Hמ���y���f=�)����Q���,&
��8��/������kHOd�1��ƶ��K�\!�#� FO����T�(y6��e���R�޿	�����E���gO|FR�h�e�UU�m"�����Y@Em�[�z���~�Lbš���|�H�k�Q��ikM$�/Vwf����Q=��\�aA��#X������
�^��#%`�q�FO�$t�$��lr k�|4�d�pd����dQK�;Z�P��UF�͑��іp:����\zl�<$Uoi����^%�O�oa>:o�c�D���'3� ��	��,��.�}(��\�)?/���&;�xp��sU[�,(����0���܊�W���b��C̥��Eu����_̜Ҩ"�%�ݦ�(��eѬѪd*�����		���;����R�u0��(�8?N��e~���Fc����Y��f8�Y�D���@۝�m�0�qݫx��W�C:=�7h��#�Oc��� �$��~��<t[@cq+.-����1y-����ǐÕ�$�Ԟ�h�!�\�З�xrQ�ɨ`��'��RI����}�� f�#f�޲��:)������<�z��z�	[p�L�x�<����
����\��e{�@�|VU�G�������C3PH�''S>7�R7���I2����2v�*�#���|�kS�M�=`6����lp�� �����P_���lJ&'{(\�Կ}�B�79�w�����z!['ڽ�������1���A�m�I�Ũ�X��:z�Ťb�ʹBf��K(ov�0~���]��ݑ
x��lVg�Y���D(�Yi���᪳��J�\���nl�x2Ĭ�
�2�V���y�B��_��hzQ�?��v']��V\�:N�:�|JT��S͉�7�ȑ��Og�afI�),�y$��}ڇHxΕ���C[����/����֒}�����5�k��k
�[Y��y?|�c�]'�U k�	����r��H�r�PdQ'~C��Ov#��ggO�� ���en*kv��M�6���|��[J�q�'T㊂ߓ�tV�00�@@���L�FdZk�-�Gv�:�SP�������DQ 2Q�-�&�rS�n�>xM�]$ߔ���TY�#��-�������6/�;��!��waǨ(�׭������B� �3�ng��R�o�%�n�@n�x�z`\�vܞ�E����g���m&iۭr5z���>�~����2�k!��K�v�y�F�r5�-�&��:�
"��\Ɲۺ�ܗ=�Ҽ��`�iD]l\Y�/S�V��
Z+��n�\5�Y5ʾ+���3�}p?����o�r��@�c�Q� P�-o�"D�#�q~�Kg�jX��7����z�uC@�1�v�͓�o	!�9�%����n	S�vA8������<^~�t�f������Y+�c�a�;KK�Ѳ��[���sY��C�[¥<�E3��]� J^�}�D�X�EeF�P�̢�qh;Q�	bl�.4�Y���z��r/|�h�d�4����3��� � I�ENH��M�\�B0K?*�fK!�$���Rxט��_Q��U�r����y.ߦ[���c<bp��� g8Q4�E$�4$�M�<wЂ����P��G�A6�_X ��������N�hԲ��ָΘ		�Z☦�-=�`ZE���
�	@(�׌�2��l�@�0���a�l��	���ok���Oz
d�8�^6��O\�&��`�?K��AZ���5s�Yr\�� *�s�["�5`Ʒ��[��0�Ohqջ�=���^��1t}qRY�]�h�:�Q�~�����Pݣ�^�V�e��ٍ�34]�RC��VV�������CP��F^�U�m�$�}����$��e6P�0P��O�Ϲ*+t{q�66�J�n�V2����&'H��w��
�9T��h����ϔ����&(��Hh؏�;�uQ�ob�X
m�ɷb2K(��s#{�\*ڋ���<Lb�\��Mzn?pz�\�Yf�HRT���@�I�	Xa�Zd�h(���m���a;�ya���ħ6��e~>$h~�/�<������Q+r��O�{��$ΐ;Xy�imi~)Z�3�m��)!����c�����jw��4�id���o+-	��H=����'��Q�"J ;"��:jn��^�=}�������<�g��s������5�,��}ʥ���8YAݫ0Sm[��9I&�m������	҈��A��A۫����uL�I�'�5Q��\�s:�-	�g~ʛC��&�/�ā�(-�1�S��(0�<���!�����ŏ� ���vٕI�U]��n�ʌvs<<|0�Ȩ'�;�����f�I�����$+f�~1?=q�Ԝ����������z�e�Eq�ci �٭�{�Ĝf$��c�/�mᲖxlE�x�'����pǰ%�'>��T�ޞ��y)CP���� �,h�<[�' �Ne����X�2¢v �G�G�v�����8�`�/!�ޞ��ڲ��g�y� GN��9�g��-f���M��QR���#m�_��`:&ԫ�)�k�*����j�.S9���G��� ��&7(l",�]@�agRyC���R���dn�љ ��+�b�˦��gX����h�=ދ<��KS��_����j[G�`�}�!��K�2\����$s�LM|�v��!TNl��k���/�܇`q��Vt�/��c@|AH�����)LCu�/�Q~����Km·��Pq)OQ?a(��Ą��]�ǿ�ʒl������*u^(
Q��LqI''���E��+r��U7�t��7���9A.&�L����#���v�}QdMH���H8\ҏ�8N�y�\,����7-(��O�A8[�a��c.9��D���4r��޸|�Q�h}������i���ݨ�1qb��
S�Y����K��[�\�~��+���'���?C��V ���՜<}��v��7,�on�����U:�[�B�����q"oYoɏ�l�����I�^�n5?.5�y�407֤"�R7c=�U>I&D��z�Vq<T��H�%G6�*X	�����l���fٷB�
-�v$������z�mJ�H^S#�NcOD�Ѻk��*���֎�������̙	�i_�������1�l�� �u�3��v���HW�+������F�Qۈs}�:��
�&#�`O�s�h|ǉ��Zp�&	l~���`�r$�U$���k�3T*nO�(vPxG��d�g�CH���A�����
�L��f�0�`��tr�;1%�n)����h����ob`�CǄ�,����0����*j�t]��7�\h<��K�z�mˏI�_����Q�V���+ :ť��0�;؉][��nN~=�F1@豩]������߂+Lh~�jV�����pP�'���`U��RW����K�䛖e�s[�*%��cŎI1�Ἀ�ƫ�OY�~��[�"��TQD�7P�4����!�rsXͻ�^<��_�rm�x����ǻI�,��r�d
-��o(-<?����WN��a2��)?C�S���<��;��=6�<����nd�Z�r&�ϯĥ]^Ew#M�/N=I܈�K'�fE[W��nc�4(���E��G�V�!��^��q��]=#�U����=g��������:�Ʒ���Q]��$��u{�T��#��U�8x�h:�X���A���>O��pг�� nX.")��=���C�U��I�m�	��8�wjm�7�d�I3'h/;�M��R��#&�F̅�A0fG!�S�M�g����6���#�_r�p]tf]t:�`X���l��d�Qo��6KNq��D���Ԝ���G�]1���rڀ�`up;�x��&h9'�����c�h���q�N*������:�$ ~?�k1{nhSS�!.��>bkW,@?��q��Y�	[�k5���:��G��y:�Q�6��y������up����y�3�)�E���Μ�\O����ɱ
M?�D]�Y�Ͱ���vzWȭ�-��M�0�]� �5���Q�V:�x|h;#P�|i�[��x�Y�!����1�A�����i�C�pS�2��w�b�ܸu�
Ǆ~/9�� ���@����x�-db.@����L�&�/��
�^|���� ��E��_���@����g>���2g"�����9�����`dA���B=6ro��4�>��n<G�Y`�1q!k̵z�^(_S��f2h`�g/�bxb�W���AK7�&��M�`9�g�?@���y� �$�8;y�
���f)C��J�����-�_3]�IS���g����]qI�4�P$��>:�dfM�ƫ��!��bMBH�>��	5�Q�%ą�̕aL��:}��Tu;��KB�����g��[ñ�fw���(t�j� �H��"7VrҨwR����8}#u��K�ܭ���Q]�`-��U�&�?�)������blv�h�G,ٱ'�q_	�Kܡ�m�^vn��-�hL�����#]��TV>�5~��RԒ��DH�t����w~���؁l�剺M�x�
�P�H����%�_�+���Ӯtx�
�6�z��xmᐸd�����^��yVVr���,�/#��>P.x��^C�;�7��Q�d��/�΂�
e䡥��gI�,��s�쮌A���k��R��ދN.A�����̺�A
���Z=.g�2�]�����]EZh9��N����X'�>}@S�����lWX��x�x�������dd׉9L#	��+�s[�0�bh��nx�ϴ���+���w�A ���ȯ����W�����*��\V�}��҂��7!GjUȱ]#��7$�o����k:��w��0f3X����S�@Gݭ;�èl��
0u߁�0�ǀ�l�Ģ���G#���5���%"�Z<~X|2��ncD��j;�P��p[�U��+����[c&�d�c4A�&(�K�3����OǮ��mh�6��6��i�0*�	m�E y��8C�&.\���~�����u)^9�*�V�������m�����=��)8��6b�mj"���	R��>@/ҡ {oM�l�=�<�m�pA�J^Y�C�V�H��@rL솥�\C�(C_��u�ݛ�~��pl/B��Pƶ^G��hYN^��l^gE���l_ʏ.�� i��I���'��t�`�
����Y��r�����]��_�&�Q�O���c{�9k�.��_/��T�����H}��2�o�������pX��G7��xS���o�������U�H
�.�eqjC�,٦��W�e:FMdc,N$JM��zOg�HH�c���2���l�ڪ����`_R �U ��mm��t{���r�\)�$�*y�0�j0lK»��9kbĸ=0��!8q����l7�}�l�0�x:�Y��`Ն��X�fu�f3��"c@�fu!g���,� _.o����J��3_��	<�t��,͎;Z�XW�%9攡p_C�Ȟo�'#{��?�3 ;�J��Z ���V�b�/�f�<?#�#d���Ń0�ǀ����:��,���$�Xj�'yik,9Q킉�go����Y�\@����y�
z$!R�Ya$�T�p>g�֜)(��Qb�v.��8|�eZ���[�U!�\����Ȍ�b���$y�|�E�{���4�S��mz�_x>����TJo��皢"�*@�ͪH�6?�-��m-O٢,���|oh�=o�
�̀��j膦�Cou;��"����A��؇�E�$�
������0�ь�7�-��V'Y|�`�n���ɼ�43�O1^�!y:�!M'��wt�K{lU{��.M���\b���0���)�N����
炕�S�f��{v�?>�1�&�^^!���Ҕ���h��8��k4"'r����}�P�<�g�Wr<06�fy���݊��w��W#�rU/iڧ�}����C���U�c�)w�_E�zM�d�Hʖ%�
�U܄[���&�‍���U��(�p:�D�
aT'(��2|�n���P3~���4��4�L'��6�^�%��Dg-b��K�^�(��|����4Ck�56O����)o�K��gD��e!T�4W��y�
���2�כl6����w�DE��ۙ��@I�i�>�,+�b�/V�sƓl�b��N��rjc����@��ή�|%mt�K�������/��9�I%��/�&�������[E�@s���8���޳;>�(Kd}�'���N�N_���ب�a,�,�ײUal�X��C�`W@����D�\h
Tށ�jk�>�j����%Sy`�K�(���_O�}%"�Ԁ�R��I~��T�/�#��畁>":�g�����T�ۈ�ܼCê��?�Z,�M#`���x��N�>{�r�+b��cH
�S�@]H5�Δ����G�;L	�㝦*��������=s &���������g\L����ؒ� �p����=��T6��(�*� t��|�l��~~O���$� �A0���!����d�,^���a��k�D��:C����b�=ʵ�阰��]^F�1s߉�B���Э�8e@=#+���zL�	u��: �g%N�>�%ey�Y�n�%`ã١)��r��Ѣ6��+�畫|����N-�ڇ9zT;�Ј�RMR�ƍ���3�iC:���rR�����'�n��N]�a4�,��]��C����"�����0#+�A�-�h��Z�q)�(�՚�JÍ�EZ�D�dO�V̕7��s�s)1u ��-a�ߞ\�i��f����Wq0�̣ȞP1V�3��:�q��w�5���sq��{4�u��zH$x�x^�]�8B���%�҂�H-6%��P�*���Ӧ�jP�HA�!/�*2��h�΢.ޤ���)˽q�WD3y�w>����;��>5�Ĳ�u��X�K����(�q�|f��.�����s9!ȵ���0�A�B��8�y�9}���T��<%�rI9�D]�b���C��.�����BV�췫�,��kE� b��<��5%A�	���Oj	-ǹFu���=�2̔�uE�S����Z�_~�3*�f�F��q<�ͫ����e���I��(��ב�{��c˘D���t'�c��~+�k�'����÷���*Z}��n��<#��8pE�w�!{����y�:�?B|AI� �K���`��vR$E�y�v�Gs�����Z��n_^����x4�C�M�K:7 ����3�!�F�EQ���Rk��L{�o����ȽA��
�^e�l�*o�O�z��v�]���d��@���_�阎4w�	}-�ɣ3�Ve��{zܿm:{�F�o��'��P�7i�G�Z���p��x�G8�+�D�H�D���m�<Ŕh��*�c����k������	��Vm�U�I�C� �̣�� �O��Q�I�=Z��@	.W	\@b}��!��v��v0������Ni��f��$���h��E��e%2�YUj��`����H*\�>!�V�_
���5�#V-H�v�����o��^���<Z٤0I�"��,��E�7�k�� �SY9�������6^���,�o=�R�Z���ϋ�"�`G!o���p\rÚV����2�S���SJ��*�(v�o��vg�I�nfD����0��ҬWYĮM�7�EU�v�ȗл��Hݗ�(D �均]�۬�Fk�0W6�!�r�BΊ��9��+����� �:HH�wq̰k�Rk�W�yq)c$��ՠ�ԗs�)S��r(���N��Ę��Wv2�lhb���(�oq �i�Άr8xh����gt�=J��H�I]ju�/�.�9��0�������Kބn	��q��=��n1���E-J}���~H9~� ��_�Ր�D�w�`�ב\6�;;1�����6#z���jr���!�P���� `Z��ޝ��~�x���[�!��c�ŏ͐zgvDދhi�.?А��8	�	=���Q?m��T/�+,7�WA�$��j���c�
R`q~�|���wH�!�#�wr[����z���5�
8V\�ۚ`{Ilj�
XFq�� �0�D����[�F��쾶��J&�«���'��8�_��eK]���bSw�̝�V�����:cmd����8d{i��4�#A��]7z����K��Xt�戺���G	O^#Z����-nl��m�67*�����v(Yח�0�p�8�r��WY�/���i7�O��y�rE�l� �V�~X�p���W,+�x��h�%�B��꒲�A���ba��L�)�>�C)IAr'l6�5
r��(�n�x0���nt*H͒��hUx�g�G.:=�����\�� G��3��{%ɥ�'/;�Yӆ�eݲ�hh��ax)Z�!;.�L�!*������v	�ߘ�P{S?���V�r��[~ѽئ�N�rB���m����E�[���C�1�ٌ.�U2նY���4H0g�)�����-YK�:K�����A�RY�Nn,��8m��ꋹ�����/�n�iɄ�,@�G����-�}����7�p�ZvW*�3����@/ �vN��6���I�q�D��������/5���ďj��c	2}�����Ws_7H�O�z�G�<�u��H��f-rH֕Z���5�#Ai�Y zw��r��}�O �n���xQ!���$�$ Y(с���""���M�FMZ5���\��x�t�|���+Vv�e���e#�S-ꗿ���T�Nj6b��Sde�ͤ���+pR���ޓ���bLG>���(��/��l[��%_?,�� K9�b���i��;��L�6*���N7�L��_]�GQSsg�c��t��=A|�|n�>�J�7Φ«h&�|�������x���r'��yB[^�(E�l`Af~$��B��wͲγmɀ[�aYST0���J?5����#^w���ћ���q�'�7Pw6"��3�נm�i�}˫/D|/2�1��L ���C�e޶~�d\1Z�(.q;��6Ŀ�a�����x�v�yǽY�P9Ef���@k�E�J�'؊�۠��w@%:�{��US��SD�C� ����X�y9��c>7� >�+��r�3]�3�~�%!w�_^H��c@���#����Yv/pk�0�M���~���%Ƶ���,9a�^?X�N�h"Z�T��H�2ɮc��.��������H$c�,2�m�u��sK=cJ���F�MU�&މ�����)�=<�����5W�_��68`18��<���\��-�"����d���&�,;�^���