��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,�9���/���]N��E�]שF����1Z�#ߢ �d��o2����TS���(� ���3N����$�F5l�@
r9|~U����Q�d�ݮ��+�4%��C�Nx"n��<�.�����U��0T��'���w�Q�z�[��q0(w&���|6BP�4=�����ٴ3���t��W	�Aت�� ��a�͌�09�\�<\����� �f�v���%�z�M�7�:A�����k�;W�qNI&�Ǽ���Oj��PuS�ق�ӆ�k�>�N�ɔpe��$�t�1ĺǎkޫ�ΔZ��I�5�u9��D汁w�#h���,e��`���/k���ſï�&Ǎ����tX�.U)�yF�b(Ċtd�}�v��_mSFf�b$��j�ȺN�ŭ���՘�AH[Iђ��J���s�y\G4��Y^���̖� �r@*�I���t߾���ټ�g�R�=��G�j�y���r��o8��y���_�y-F�z��eә��	L� %y���r�m���c�"���H!%"�ǒ�$�TmP
T$�cx%/u(�#�,��s8 <�d6����W$���3��B�?A�2�5f!�Hk(w�I��S����5�i[7ݎ�5�G�������Lx��� )��y��t��3x[Y0��թ@!f�O����kG��w�V����ȖC+k�GB:��s��[1���Ĝ2��U�~*�trs���dZY�1�f��93h���/���D�k�3h��w���l�k�]Y��$&�
Q�hN���gOD�ql�56u��G�vI����w�Ů���'x]M��$��3"^n�`���`�}�DX�_݃/H��sVW�>��j�����@��7��]���3M��M�F�c�b�MO��#b5���]������eBn�)���R}�>�4z�/�`2j�5y��V
�p�Y�*$����/�����Yr�u�
�� �+����Ec&~1��S��mkv�3���:\1�я!�8�bD}jQ)9�V7C0� 񮆏�9�i@D�����R;�{�� �^���7�{ԃW��xX��qc	���{��B^���*i|�P�ͽbk1�ڝFf�Q{�&t
��X��p���Z*[�	MR���P��ƅ������+|�}�hvr7�7�Փ_����QxH@�����!��_6�(�a'ҹ*���O��k�յ�W{�#�@B{>�c氒��#�!߶��o�1��#;8���v�8%�-�x��R�D��$�"q-?c}��E�C|H��8<����7Z!�]���E/L~��G2��7B��n�"KKw����	#p���lb���E��9j0�'�Z�9�����,[1�-�T�d�3��Z.3|�+<�>�>����z��ݠ���] ������{�2��2����޲%�5O��~�x����Xʙ�	�c�(���3�<�KF �����Qn�S��p�kIg��M�]%���V�t����I��'4N%�H�����	���E@��i�ԫ�4N�
|��#�8�#�@:�!�]�O����[3P�$7�e���?�!KљZow��S�� !�8��m*F�([K,�Z�׆�}Kv�'Ƴ�(l9���DXl�p涭�.�Ř�A�a��9��AG���cGޢ�v�!���3Jq�Q�zY�u6 	q\�f�JГ�~ϻ/ᠨe�;��?��_[E3�4��'o>�q��%�t�^(�>��ZyC�rW��Vl��N���}�/ȵ�����"o|�u�ew��OSI~|n�7�eDm����+쯙��j��щ�ƴ�݀y���
�1ψ�Lw�phGn!w���ٺV9v��N�`��Y��T�f�hE˼��y(���Q_�F�
�':)A��cy��������uҝR�-�+���)x��kN�g6�����X3��n��}�eM}��Q1^�%��ޣ+l�|7��IaS�_�w�!���W��O�;1_`��s��,�}f�P�� ���lt�6E�t��C��ц��G7���s�O�ٗO�B��>�2>"Y��[ �qp��4���z���������$�pԊ.�/UvhH��}K�V�w1��>�^���C��~q*kdS踾ⵖR)Ȩ�q��%
�,#!����@B����p+��9s�{��~�X*ۣ+�3ٶ$�4��� I|��E���q9�S�-h0ȅ`�H��[�@�����'���8���C�Bu�7+-wX�	J9n�^C�^�[�����e��X}��L�L���Vo��!j��A[ݴ犺u�E	��^��O��WA��R��Y�����������u�"\n`pg�9����l%8G��Xm��JD��9V�]��s~ǰ9q"[�~��d�=[����~ρ�������t���ըd���13���q�u����#Z��|RXQ���fv�Xy(%�������_6���M�w�cw"ҁg{��?.�{�q��iW3yn����l�{�{�R�v���}�`4~Xd&8�>q��y�3�#�[�Qg����< �.�R�9�?}�l���ocS�zF,�'$����M�������q�w*ծ5��Jw>ker�����P�Ѳ{��*C���L̟�S�a�!�·-��\s���m_y��N���K4t��ީ�"l��ED��i��u�"%�=j{;�.�8�T#_>��1��2�Vj΅�@c�ĄʀJ���)����%�}]����˪:�ydL�;歂�& �(��}^�!�C+��}���_�n�2zJ2�B~D��i���̸���S������*D@f���1˿��4�7Yh)Ur�i�����@෶���9$#���-�3��b<&ߞ�I��|�p_�;�� `�Р#�(ԁ�k#�1�Bl�9\A���e��5�R���Q�̸Q��w3��{�\o14���?Yqg��Ԝs���:iX�%/��g�KK����+L��Gq4̖^�u$@v�6G:����Λ<7�b�N�950r1_��"D�;�>eλoΐ�ͼ���+d�K�>~�R9U��?W(����`<t�OͿ<ڨ݈|~;Kl�04�j�Htn��~���a��shQ��B4Ǥn&����Zݒ<��82�;2�b�04�ne6�]K%�u���M���\���X�Z��9ٔ�PM���'p���-/bZ�TC@XwL^^�W3@Z}�����F)r�����3G��G�o�O�v��T�O��>�B�d���є��#��8&IB�踅��ĳ^����;�����O���?��:v��-�T*�jR~'���h
����Bj^2b���!O"^Z���1������ǄI�}=� �������44=��UF��s�ŭ�X�t'���.َ����`͗x������t��U}�mm��R{P�z��w��_ȧ�=��kj4����7����!C�*T'���Y��He2S�1��n�(��Z6�������`�qDN�����I�H		�)?s����m ,Y�O�D1D�Rq��·#,��K4
�x���yJ1��N����D�G�~����ܾ'��A�P߯�%� ��^Z/n��٭�6���^T��OR,~.&�wk�+�ըL/A�Y�LsN��*��S�$|/	����If�k�����������A�'/�cT��p%��?�ul�BW.ӿ|�b��Ί�`"�("^�
Pp;��kiwq�H�9t�z����k��5]��q�r���&�襊�Y�t��8�o���Z#6p��̬D�_�-P���]f��xk&�m&�l����S����0S蛏Aǿm��0�~��,����g�|����L�эV�&��~�{�Ѫ������NB	�{���C5����o��Y�d� �5���2��PC�Q5��Ms2:*���[��s�����M*��#�Wax%s5T�'R�&�����:�+��i��]�"����g�- �bH�L�!Z�I�aD�g��p�N��K@�
��b((�t׃=�T��<cĩ;7�6��/,'Ɩ�*�D���v�Y�h�n�y5�t�k��|V��a�ǅ
��v�r6�]��7^��7p-�����p��~s���E�Ϻ!�*��&�Y�����p�J�3��\
v��Nsި]4u4��K E*�C�n�SJ�ׇG��v��ۥ�>5c/�a|��Pj.�R!}�/,o<`��� F�E�H�.~��wްQ��V#�����`���-YZ�7��������i�R�_%>yh���9�"k�Q��h���y#���L��u�p��~V!"��q�k�]����zl��U��~D^�`�Xd�q	V��4��\��vGj��/�[���b&�K>�yn�����~�Kļwlc����Z�A���b�E����4.3c�~F�ƌ�irkwllƐrPL.�lmF��b���p��o3�]b7�:JY�3�kb������ܽe�r/��;��S]�x� �;3z!^�}�z^[_��D��q$����i.��
!���!�xr�w"�_�A��!�����Į�?�� �O�Y���ٳ_Iq΍BA�;�G��Ĵ �
�mm�E{p%F͑�l���^�␐�䪃���ƶ��@���N��	g����	�Bx���VO�÷T*�C�����q6t����+��I����]�
�*>}&ՠHJ>�Y �d���9tYk~�Pp)�u��F*��[ �]+o5��S"њ��8�����ʆ�M�w\9�4!��T4\}_��hQ����`M�4����L5��q�i��@�0���I��?�I>E0�GD�-�>o%)��=E���6,A�?�ܛ.��K��D�l�W�l�`�*S~
�\��59�v����_j"�8�J���õ*&U�l�������)�['�߅h������R�ğ��޴�8�T�i���	.7$u$jq�������#��֍�>Q!OHc�E.h�qC�.ꦾ����@�8a��,ՒY���ǬVH��7q��뻇���\�/Y
�O[[RĠ�l�)�W�(QH�]��&]i9�7\�-<1'��Cڪ�J��B�m��Qf7�1��T'"oTWbԳPz����\y���(�x���#��^F��qnp� >�'�Nh��"Mމ�*�9%���.$���}��G�Nr�]�H���s�РLp�uT�Da�I��N�G���Xј9ƞ�x�;�V?E�.�Ņ?˦��0V!�iM����]��&b�?�0k 8b8��_і@��j{6"�6U8�x���ɼ�L�Q(�ٲ�n��y�)�w2���4�)�����f�?���,�ZO��Ck@�W���́H�y�%c��G����Lܨd��mh�����r:$����[]\�؇�]����k�bD���0]�Ag6]�'��/�ԯ��3�$�W��#{�Ӹ�8��(v1I�㒭��3~"�>A�鋟j�ǁ����n� F��uƋ�9�أ$��)~?O���0�?��I���uA ��i�A�&;l�DH��I�)�P�_$d��O��8�9�[$�����!������5�$�%YM ВJv͗�Hn��	��*7��W�ʿ�8\��͉ʏ>U8���Xbu���\�gqk�z�����Ϯ�~��¢]_څQ��}8�8B��:n��<��޳��D"�<�%�x��m�ܳA]��
�_�)�;�y��E#8{����C�2ˤu����cg�ּQ��홝���ٜ{^\A]rh���qT��k-}�@�-��$-��@�i&qꈞ�X���B�~>�T��8���[�-��/�gur@^ⵄz@�-��e ��8w��/9������?�P;�}{V�י�l�=��ٺ��[�o$���ۀz���
�V20=i̋g7۳t��*QD���X4v{���Z�D����+_0駮݃@�#R�NK��ts�5vY�O�ÎA#ؐ�ц�
'B�������U�7�1��NХ	qf�3��6A8�u�Zm�NX������e�y���l����Y���>���X�GRp�	:�N}��F+��}�FtP�0P���R<aw)~�F��C�eW��y�Њ�O��ѣ*�n�����^��6���}�kK�4o����H*��ۄ�����]�Vy!v��x/�ǣ�I?3�W���&�n&L�R����n�����L�ߨ�(��.uf�ͲV�#�֪]
��6���j�#����"K����*J���u�{� _ �v�EXRrΜ�r��2a��ܢ5'�o�&�ޥf�^���_k 0��"��������1�-D�˫E^Kk-,X��ۮ���{��ʫ&��F�;g��$6���!�m���$��_n�6Q�eKZ>7)ҡ]�V�B��� �S�\M2�=��|�c����O�*����o	����j|�1>�'EnR(�beo�?�L�?�=9��*���0��cU�$�I(+���b:DU�}�ل�L��d�XDO���p�6Ti��I�d���S!o�����(�f-�4���A>w:S-�D���f��}�z�ﳵ�l(j��X6M+�E$�s{�>H[*yN:[&�'�'x2�&?x�#f.ƬhN �C�/��ag�+�&b� ���Y�޳�M�Ӧ�/;�?���b�������9��d���B��d;�B���Я�rP�
kӹ�v��i 8���n�px��Lاt0 �Οy�RNԈG3���ݎ���A`��5̢��\Qs�T���櫫�\��M�7��&͵����J�Ts2L���,�c!(|x��!IR�V�ӫh >�f⌞{>��1�^�6�^�t��o�:�z%j[�^A��!~�L�5����j�m��êHE2ly���Й�z�b[g��k_P/��$���뷋��#�G!�z.����Ji���Q�q+��4�fc_#����j�E��4}'�o��Ŵ�?���S����ƕ`�ed��"*���>�i
m"����
�or�h�gU�J�Ƅ��U�y��*�(yn�#u� :�4�CTF^�-C 0Q��÷?���_��gc��7�s��^Q��M��3T���w����J�1 �c�[&�fy�Gg���M���Z��:�-��!����G��i�	|���+�6HNR'$rG5Ȧ�B�����mF|��%6B��"#�"z�A%r?���� ��_*e�q��>��6(dc�Q�U+��2�_*H��ٻ�xf�Ƴ��\���{h�N���D��,��E��˸[>
��<�",P�s��D:�B�����F��(��� �+�C9r�����W�cB 꿨���||�<Խ��PN��-��9��T��<�?1�����@��c�$<�����
�<A�L�����{K�J��i�����؟���F$�b������� �*��ʌ"�o��鮀!kp��>.�%s�s��и�et�a"���p�H<U�P�6�������c�֎>���Z��4��0�5��mA���Ң����Ȗ��]e~E#�����@��7:@X��W�!�����g"�ãˈ����C#���,�0q�X+ �;oY������w����Κ�f�K4�Q�H�nH���B�h����4_��7R��]��L�˖˞�)^[}��ڇhZo�0}[���ID1���X�}��؄C�W����������c��H��I����&��F�vEE�q��u��AO�鞭۱>��e�cL.Qp<���"--V�#��՞���4od[���,���mvM7�?�8�
�9[�ŶJ\3tm�_�]��Z���c��¸�Q��Jm�cɎ�V�N�K�36웆���nn K�P-f� у�B���X$L�+<�j(<��S�"j �[�������6��N{	~�,�Zo��a�cA��4������M2�]��_��|�K@���b�|�" ��#��
"��Ӡ����%� �uQf~-r%����dG@���*TC
����(���j��1���5z��_�/�b���C�՘�/_�<���{6٣9��%�e�����w�*������8��i�s��w�.����94,c̳��h�5Xa�5*X`�i�V���÷���Hu_�E,��
�_-2`$��r��sZw�HE��g}X6�Eu&r��6�0�ĦVx���wd���&Ƃ-���B�����l�+����2'���%�����H3��a�΅ݯ���o���Вsc���jo 9��{�|�,��'��!@���n8 � 3�����5�0�Jق�����Km�t�l��?�V�F��KtG���s����n��������.���,��D��>�B�\���H���lR��{��$��)*	�:��jnV^��.H���nc����R��e6���k�2��e)�g��)��q�*�-��������5܈�x�b�����'5��9�A�u��O.�ӿ������Ԫ��Zu^<�IL��_A��9��{,��y:>[�<��2#�ޔӖ����p��hٛ��<���Y�I���^b a�Ճ�A��q�H�11�8!�7�xⶹ��8�"P2p���V/�`�mm�$����c��
 O;>��w���?���L~��m�қ֯�!�Q��Dģ����*�Վ�Kđ����P�����P��\�������h/��.̠��E_0R�O �Պ�!���/M��B�,�_��ٸsI�YtF�:=��������T��`VJ(M���a�� IC�!�K�d�6�#A&6$y�X͠9*�7
/�Evn�����;3C]Gz�\%�E��)3{�MM�:�)�tK�����������-�:�_�k7嬧�.�>&��_�eԵ�=)�}����Joy�U�vd��u�˄8G���-!��5�p+���#ek!xyѭ�$f<5���H��C��K�WM�6J~�`	N:�L�{-�$��P����>﫩7V=���*�Q����bѣ
�G��Fq̀�WZ�c��1B#<�z�G�[� �.����e
���x�w\���wN�\$�;�4{xA>�~_~T�A��gE��y���`t{�(�ܯ�����vԑB8�Rߢ�n8^8�5��:�ҋ��G��/��O�^G��c��)��Q}5�#8�?N>�v�]�i?�5ܙ���%I��Gtw�{>��U��	�b�Ŀ�TD�3�T`4a�h�vB�1l?�JPLm��ށ9�}= ��Z����)F1`�E�?�x�~	�j�d�L��"���_�.300�0{��w,�N��S8�_�B527�Ԑ��V�� �G<Lixg�ߠ^yy�>�����x�K�:�4Hi�'m���oȜ*u�Y-��h�&�;y�.bc.�N";�mt�B��`c�D(�̏��e�̈���4p��3N2��-R~ኯ��zZ�3˶��N8�d�ب��c�	�)i�����7UHa����	~A`D��Zk�x�?�H�𞎟(zL���VCA?��e�ͯ��w���ie��V��eX�u�!��y�hk�2oI�^s��q].�Y�QE'dFz�$��L���Q%�oT��%�ް���ik�?����vH��l�$�ڂE�R�x���W���ڭ�)�%����
ʩ�����R讷*��������@�E`Y�C[F��\���3{|ڲW�<�?�(��3����=������O����1�R���Ac[�8X
I��I�(kgU�Qc8 )ގ]����T��ㄫ�

^���wE��,�f�G�H��f=�d��ߍ�̇�pb88W�@Yl;�n�l�}�A9�qK���S�o %�ɫ�C�9��I���X�Xt����`��D0m���
Q��O_ E���ȥ�^d���tD�Dڊ�?�C+��߄b�&8����y� V]���(B�H<��/����o9�Ŏ�mW��Ѫ���gN����!�C�\˳)��9�Ql��k^
��74zhY�~�F6���m�{��)���a�����z�Z����k��9` ^)�eGI���E@�5�7���[ZG/�x�s��^v��S4�kM;�P�e	젭:�ȩ�$7?&r�4=�����OxT�=�ǢG��2��z�m�Ǡ�d=<q(�S�������q�:���⑏#��7��~J�A�V��Ũ;S�*܉���!��_�2��Z%�P�f���
 ��S��W�6ZԳ��	���g�.��Q��ue~k�m,��A�g��3��Za��V�cڨ�Y�*��boE�>��ﵶ�"j��L;:x��_c�	ĉZ����4���3B���dS�V"r6��|�_�o0���Ԟ,���$�ᎈ����{w�щ�&B-Qx��+D4>��!�},��C�>�B������q)K��R�p|��0ԣөX���l�1D�;|Mkzs���Y�g]�Θ�,aW=�9'��m�Xp�����02��
���+\z%ěUX��3����듲BT`�I.����7���U��W~8ۗXg2�%�r7�$�%�MۛR�r��*B�	3�n��X��ܠZ�M��
%�قh4"�Cp��Q&
k0'\�$4��٣�5>Nmxv��M�TL9ZN���8Ż�b�2��XR�ZJ4H3�	t�&���X�#e���7JB�Bt��&EF�Y��>�Iz�d��`w�v��ӵɀ�j��{���e��ԑ����Z��Зd�h�N�0s*۹�1Qب^Ŏ'(�N�6� t�OEK�uT���6�;rxY���'@����ܰ�A-��LW	�kq`^:D��UTW����ŅyC�ŷ@71���L�j���C2=���?��h�{�@�HCo���.����t]h]G�2aS�pr֑tb-]&�3����;Pd���	��tz�Чm�82��=pH��	&��	�LIzk����h�2(F�{��ƹ��T�ho������mN�m��ə8:t�se��i� �8��|�>\]� w�ﲥ�tD�]�;)B��Ss�p��҃N�P�%,7	D`�*�|�E�"	�L�)��r��ʳ��x��!$�r8^"'.�ݽN���:�:��rn'Q�k�H,���
c^�����g�a	L}�L��V�Q��t���]Ov�����Ț���h�2�������1ʶ"��Co�\^����L�6�-��\p�d�>wO��◘M��c,w7�i���B �E���f1�Ά�-z?�b��\vB����zz%�XU]W�`N)� q��K��.,	:#��%��-����UȆF�G؀�5�>�m�~g���=��%�&I��0F�q�|?j��Dnݞ��?��E�Ki���d����,�H߃vh��[%+�f4-�&�,�P���ch]HZ��F��!M��uG�[H�T)&4���)�7D��C�{��v�_���%�8��_�R�˳��d(KB/l�v�/..�b�R��Ui7̩�?�F�d����b��)M�i����8_ �E���4��)/)���w�K�U�g �5���M׌�T>��g(��Z��3γ�ɡwoC(���D�6��&E��M�B|�N5�&q�,���l�B}^����R
��n�*���.��C}@G�UL�^�)�,o"j�6���?�f��B����2vϷ���3w��N�5X#��R��U⍌��lڜ�b&��"�|X;�
��?��jf�Zl���&��آ�dE�O4Q*p�fgA�f�Κ�31a�?����¤Q�⑊���r���$����2bʛj��Y�x'�{"f���&�!s���Q(L�n�\/����7�^�;c2�檘[�CF�
Le	#�P�,ͷ>9~�w���ϐ�8I��)Ͳ&6
�>so&�p��qH��(�_Z��?�A�l�dK���E��#�V�(�G�