��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v�����u|�K3���r-g���$
轤!Ӓk�������U��Ձ�]�ؿ�x�ɻO��6�N�D_|���9 ���PF�S�-�G��.kF��Q�7�E�Q�a�!zQP W�E�l�k�q�n�>;���x_nc�B�a�h��C�wK��Gt�D ֎D6�b��Ki���|�a�P�ns3l�p�jp�Y@GWD"�� ��u:��(\4�Ml�wT�y�$��f_��R�mQ+�6���(��"}X,,����1/�NߑrbD"!
����p}��7%B�xx-���P����5���A^)(�|�^Мp�;R[��E�6�V��� sq�<�qX31����u@+�D����� _-�'���"�#c�/�����%X
��j���72��DqT���8 ~w�d��;fK��Tj/)�(.��D����4 �|���YX
*;v���_O�z&̪7�x+�h�+ >0<��_���Hj����W �_�6� hm|'(��(pF�C����_�n`^�oMw�v9�d��&T^�.M�s�u���p>�a��t�9�`q��?W�]y�t�/��7(st�	�Ʉ���@L&��Si������a���! 9��#*�][�`�����&h����Ą��]������&���C����[��W�l�cU��&6t�̓��0I��F���u�:o%8	��r�ǵ3����	!"�v���ro?�{�:�����\���1@�<�wC��r7��+��(� �R�4��sp�� �MV�:^bL�ͱ�ԟQ�7=��K|,=�������	��p���i.�tpF ��KI�.�#�Zp`v �$�wO�d	$�.�aڈ�n:O>&'l-/HRաd�rv������>�-�ߔ��kr�6t��Z�b&��᝘B[���:1#ټ#5���t�Nz�&@��=�Z����Lͤ
���k�r/��B3�OM!���H)-�?G�9��
o��ߟZ�����gY�mS#���:�%�|�IG]�~�-��"��Vӕv��`ې��<�ʎ=�����xh2]j�yx?��#�<h�,��V�X�)�t�j6?�g~ IIWw=R�Ж��ԥ/���/(`�75zH��~���7��Aݠٵ�I�'9�m��r�fѾ� E�� AP�լ8�{�G7�8t��(F��}y��?���wc��|�>x���cr4�K�=,��VK�rPv��j��Q�<�2c�K6�0G�#�;�.Ҳ�6���u����9=��}�B*@�so����"#��� ���pSQ�X�B1qft�6){�A�ga���M�sސ�ˣ,�A���SA����@�ZW�P�y��~��kH��^KKչv%g6��ڡ$'��3M2M@�C۶�`�ˍm��i4�Z���d�v_�l������˃:uE�Y�[#�s�y�f��C�uK ڇ=*HSڐ���KsaRo[�˫
�(��mi�U�èl%�c�C��xɏ��?֬:�#��$�à�L�
�骙5L#���M��r�'��R0���0��j�'�!�>�˔KhB0#Ս���8p���!ͩ��\?O�1~�}^ӛ�G�j��L��-�m]�����d�$G^ғ<��v˃c�v�
�M.�CH6�>�+E���h6|g��* /�q0���n�^�N��ojM���e�[Y�p�e�s�����!h�o�]�m��C�����k�z�w�*H��:��[XT,Q|pHS+U���Z�=�����;�4�ۏ��� ��Ta�hEɪK��k��FNɊ��b�RFLP"�ҍWd�������X�"��
d�i�N�}��%\��.O4�Ze�Mh���	bݻ��Y��T�2��E���c� ��w+
���~� ��uj�1ⵝ�B9*�����o%,.w?oCm�F����|�H�8̨�m�	o��t�;Wښ�U���CGuG� .rg ֜׺�6�2�}d6� ����~^�t�:�������r�5�}O`jÉ8ᥕQ����dbu,��޷$cG���UEh�a�2�y�y�P�o]3I5o-�g=�̤�3r�Eϝr��U�Q-+B64G�1<Q�j#���Je�\N�ܫ���>�D�l�z��W5E*V��	��@缧�4!���\p�t�D@��j"Ŏ��\� �5: -�l�q��:��VmN�>>8<Pfu=,5��㿛�V�w��9D=eR`�pR!m��VC�q�q�c��v�k1�/��0���I�R�o�����[[��r��/��i�� ��?C]9��@�M	Vu~��E`\�f���v���ZT\�W2�������/��B��W6Ҙ�?)��Q�`@�M�e�ߛ��L#���P%��#���L!��R*p������l����57v��r��Z�4Z��02M��iO��x0x[�^$�6^�|39-�󈆤#zl�	
h�������c�_���}�)#��֎ب����´@<�r��!k�LV;��n�ȴHP�m��;�����ɧ��1glcb@.<T��<D&P��+�/΀6��A7�!UW�*��M��a�^5Ŏ�.x}�6SȴK���Mϣ�_���e��a4#��"r=6�=�JҪs�F�qJV��\�@Ƴ�
��	M���̼���M��%<��}E>�Q&�F���A8Rͥ'��2�I5��e��y&K������p ���rO<����>j8�S��xI&W��@Z,�v�I�-��,:��ޙ�h��4����4�d�V���̊~�g��f�Ժ�����EkOCQ7��M��Y�c����^f�w����*�5/�6�-z�s��O=jv����!���@����%x4+�h�gl @f~X2ɮͅ"8��+�x �V��.DSMϣ���̔v���v��"w�}�.<O�"����Q��ԓ)��zn���Rd���h��g��t�%�vŧ]�Ҷx	������A�3�)f���?�Ɋ�Ȩ0���n�}�kB�z8 ��ai��,�H�{�r�.T����wfx�%�R7���?²���*�q�Fz	Ebb�&��p���$p����U!qEN���n��1{����r<`�Z�ݣ6Ӧ^>wJ+�0(ma���s�i!i������{�c�7:Q����6R�a��V��"4m��N���~Q�Bmb[�m����|s�at���J~yd;����TZXEK0�Y��&�9@��u=��C��_�@��?WD��"���.�!��pQ��i�v��Կs�"�����_r�Y(�p��f�+�1����KUk���e��Ul�6�
�"~K*�<����`c�Qpw�U�Z"�G�A6!���%�8�q��?�W|~�����j>Sx�i�c�t9��	�S�vO���j�~�j��H�'Ho�{X֕n�1|��~�Yye#�)���@���PG��z�Y�P�� f��-YR� �U�<��+��X�I��6E����(�&�pJ��\jHD��8f�ւ(~v4��o�&�fy+ߚ�_2</:Bu�e:�3�įb���R����WC