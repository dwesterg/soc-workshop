��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�G�'��"w�$���9}=���	�����N6!��Y�f�c� �>&تi���3ǝ������7��21ʸ!E:?Q<a)�sͥ��0/p�7��7��v���T��$X�f�B*��K���6\�Z���w��PL3��ޜ>�!�y?05�v����V�.��U\���O��L+���~}
��k�Ry!���r��,Wr)�m�![�^B��ln���~�rG�yRQ���G���F�_C/]��:�,bm�|�v�G9�2m�'��!$�VB�s�ÓBCy��{����+�z.R����K8vVF>�� ��y��M�Ӆ�.��kz���'�R��"9�W��Z�Fz��|\'l���B��֢�T.ڞq���3�L�C'�q-�Ԥ�A���sm%F��h��h��%w�+��t�8n�x�݉.ΆM���T��; \(�rY#��Xɲ�Q"VSE�����"�����,k&�L���0�~�3��S��W�iG�ݪ����Y	nʝFHX}�n^6��%�7ֈ� �s��&y�?���X��_�������>T�z@6�eS�z"ӳ�WJ����H�T�eU�� $�z���EO0#M�.U�L8�1��x!����{�����]��M4&�CZ�v7R�+��$�;-*0�7��N��$��|Q�
�L��!�w��ubj�8�jG����	S<���H��c���n��f��13����f��s_`�*�u��>L�E���ZOT"�8P���Dvao�D�1ؗ�__Z�Z/�Zp�s�LYwME�3_9��Μ�����'��c�� l��yKb� ��J�?��0�����$ ��+��j`7>�x#$������7*7��&{IaApwa:��jG�"<K[��TK2������z���%6Ƨ::��t"F>ލ�ˍ�Z]OT�d��,�Xk�Mx����[�����Ẑ&��3��k7��4D"g2���٬a���N%6�^�h4Q��P���)[�������n	~"?s���Z[O�������/%�CMV�!�!�(���k������ņ'|�Hk}����A��@0�dc����V��?_����.䁠�.��_ϗ���i[yΞ�Q�����^�<��A�/�<U0�p�h)mPϫ��Ƈn?9����^�R�Kv�j�UK���}߆��k��#����DU�8�Ïxb�r���p��,���S��Io'}�%���������8Er�1sGs%��xM3f��Y��r� H��"����.�!�"�|O�ݽ�.N�C��q$6$)jJ�zV�jz�L��'
ʖ4�#%��Ǧ��i�rqg�Nla�O8����;G��N��ˆ��V�#��o@ 4�=)�;︰���1$� ���%ͥ�Z����/ ���e����uN4��1�7�9�t��߻��iȐ�i	�ϓ��d�B���Kk��������B�Wμ8���[��K�o<h�5��]
�t�`���$"�+`K�D����Ɛ	Ҿ��.^�K���̘�0g�d���jت;lW~��Z)��h�C���=K{�Y��_����FA O%���ވk���l�����+1����M�����y���Cg�T-�m0�x<�M�/{F���Ɓ�a��}��og�M�7� 2�54{<>àmRF8yP����փli7��Uu��G���Vǚ��%���(�xh�c?�� �����һ������W�g9<�I�s`�X��0�f�c=I�6��˲�0znG�@�A?�C2
O���U��ϸGK�����*���������.YD�,M2�Gh��JY P�g-�jM.�z�JW��חT��UJ$��z��$�;��&��GI��5W9�D�����U�.,��}i��n(<�M҃˚�&��<��{�z����Q�XRH��][��V%6ha`�Jh̢��T��֘�R�����	�O�f��6�|sY@�4�t�-l���g�Q.*��\=}�9]��1��c*��w�В�OO	����sRi�o�7S�H���,���^���,O^���/��#ۯ��B�2�D2J*���k'�Hit�%V�'�~���A��)�#������8;V�xI��[����C�8"w��6�e�5N�펊��[(6m<��Ă��g`����$Dw��_ˍ	���D�2��a}V�X��GaU���>^"3w����6ik�6�t&��G��(�:�R$:�#�|ԫ���N�Z ��g�4�nnu�o�+�N�8�,�%�o�c�4n���"�E��4��F�L#ck�!O�ec��j��*��B�nDXpC��E�g�ԳM���h	l�L��+���i��d�!�Ơ7.�{-o(_C6��r���Up)q�p>�V�lCI�� -,�aA_aA��sfxL��sق��_4Y�Kt������gq���@�/�+.m�-��`����m]������g���.Ǎ?VOx�웛��[G�_.2��jC�
�6��%$MᦂML5y:zu���LC(~�!�<����j�UD��&i���|���l麺�����&r'�<�RJ$�[k��܆7:`m/���g驀�h��*�tO�$�8a=Z��ʛ���*�F詛"�D� ���F�b�/{1;��0�[��'�����\�tH��~�o�Bu{X��֒�	k}w,V�_Rb>�4R�ے��L��U�������&d�/l�ȷ�o�ҠѬN0�w�A��E�\�T�s��"x�N�_�3c��,��d^a�Rk��]��Ֆ���/�C2C?vcq��νO�J��9�aB4�q�P���c�F�]e��;2���v���u��cЂ@f[ә��P�j�4�֔����P҃Ck�]R�=֧�Otތ��[��z���2Z0x��g�� ����>nF}u �	�P��->�W���갵j�cH߀â�����!�^���끉���m�I����_��[��
�
�E��k����K 	�QAVϸ�Ƴ7�8T��7�jѓZ�N����Z$gJ�Ma4R���%C,�N�Q��R=�nݨB|��y�۷��x� r|8Ɯ��0)�y�Ø �St�r��"΋c�B�]��m�w�Ds^I�&^��F�p�0X��!>��٥�03��xF$a��S� 0̋�,sj��a��I%���e`xI��YS��v�� v7������NOi��Gv�7��Gv?�\V ü�ChK<r~Vp���q��^�I�F�,�p����)mDF�.T8�1ߎ��ɂz��k�Kٱ33̸4����1�p!��o���D_�� �?���V9�1�<�9�b��{��Ql��t�̌�o�w�O���Z�V��{���#��s
\�%p��F�����\7�^��mn�Ӿ"1����e��P���V�It���#�I��4��Y���1<�*Ix�!���R���tTbM�!ڵ��-�r48��6_�#ڋ��$��]�F�N�͌Vk*��8�`��-��[+�,�	�Q�]\Z;=��k"��TþP�Ҟ����W�p���qL���ĻLhMe�]�[Z hh�}Su��uo+�q�,q�P�����2�A,:�_��]y�6ھ������������
�6}Xk>gO��Ʋ���\%�W�;�*���~ݼ�'�u��{�B7)x��|q
�5��/+4���Z��c���<��81���d�����*���̭RH���H+w�+)�zR�#��;Z9��
yt�Φ}�r(�d���֜�N��x��Zj���Im-/�C!���������rI��A
l���\x���8@^Q���3������Qd/�]��*�}�ⵈ{��T�_3�����睲�dʒ0��AЧ�碥�>C[����*:�z1G������+� ��h\g��4K�H�!Fǝ�_6��_�R��kߓb�E]ٛ V��v�cC7(�C����U����-,��ެ��%�&0�b
a�O��-��b���J�	4(��������q�0���|{��
��:'�Tt� vp�͢k��<���9�u�F���ץո���9��iT��'zCt�D$"�Ck�qw��v��h'v���U�dG�b�0�$<�1u�E5C�'�Y����`�����Qh�e;VJ���;�aG���.y72���á������G^�~���B��QuϪ��Dr���9���D�\�p�=�]@[�����"͉�ZU��w�]���uG��Bs��T��+x�򔡪�p[ǻ�^P�e�tѐ�ar2)��ȳ�z���O�����P-�v69/\�ł]�V��9Miج~K"u�s2=�](_/����N>��W|�gU<c����=��D]�٨�gJu����<&�K�yE4�:��K� C3��ݕ��9E�)�gp�krd��<����x��BY����˱���b)��Ѵ��'NV�!'��E���Xc�-�+�4R�΄�+g6�3���?R�SZ��R|��M���]՜)�	���i��[�@�4���}�r@��``�J�9���L�Jg˦�xb�]ut��-m���@�{���h�a�y��N�J�����:�b"�9��W�5Z���e5�r�\L�)E"���2��rV{'м]]0�uxI���X`�z\��D';�Lѐ�����!=��D�-�J�<��HЇA[�`��&V�E|���i>VV@