��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��˲�|U�eu2���P�1����J�2�@y=܆��X�n��t���+-1#Հ�B�H�b�~"�{����;GH��Y9�QR��c��ׯ�b�i�j��Ñ"(Y y�AG��) lW;#��2��rn n�c��n����dӻ��4q���狙e};�e�h����ήr���[�̉���Y~
�-�ʙ�d`�d�Y��8���N����j�B��M��tI na��#B�`��f�v����+�~X�<�V���~�����p��ӕ�i�:[�<!n$
��������2�%��A���IP:�0_*w�C�����t�q�x��A�Sh�GTo9�������j�.~��x>�W�fyN��즄)t-cWy6)����ݸGdj1��!���s
Z����YN�O��ʾ�s5��;)���X��S��=qye�ܿs a��Go�DFSg����v��%��w�u��@��&�N@8���/�C��[ ޛ�{�g��λs:�q;\���8��,�ZW��"��RDkO#�|ة�C��:�hэK�Iq��R�p����SU�Xj�	R#bJ����|���E7��H��8���s(����]��ɟ3�4��M�`S�v�Su�DӲ��˩ ���bSʽ��\R�
E�� Y��M��p0��h�$�O�a �����Mv�;��i�ȯӝ�2���:�ܵy���edD@
�aDs�u^8���c,J�[H�e�j=�mP�P9ǹ�ϼ;�Ҧ):L+�ŷ
�A~	�� ����������^��7�'VƤlM�5�ct�d��훔5�T�8ڸ�/H[8�ݣ�vR����'p╎	Ӊ#<�Lo�t-L��K�Ǐ����q��yY��½���v-�X��(I`�'�G{Ջo����S��@<	���؞��T��G�_C�3ތ�h�\`�g��S����V#�{J]�i/�@"Xc�m�S��*/�ӈ[�no����2��C=	-��{�^���ڪ�:���g~'�.�s�-�GIXAB���>_RQ�!�D��bf�M%�ǆT_m4�����[@�K�Iڙ4b�¢c�_�YBvOH2m�k�� �`�ߤ���{9ԢO��0�L�W]hZ�oc��#�>)!�!�S���y�{P�O�~�N�M?)���e���sI�d�k%�����Դ����2�b@Y�ac���c�r�M��e�b��p��]��NR��j�|I�7`��D3<?�U��K���Ֆf�J�&��d����d�hMʃ����B|b�ā8N���q�9�hj�����O�%�.35 ������=׭H2���^^R.�pa���oևP�����u���mt b���7�Ƶ���80]M]���Yyi���R�':�ٰ�tg���Q���%�"��*FD&1vbv:�ZT�{9���A���Ӗ�e�Ѩ�m�B֜=#Sv�g^������K��Xf����C1�p�C�������O�8$#��h��7#����x\M!�L�4�����Gm�U]�8��HA]����z������)'&f��Q)���&?	j�Z%ߊ.�o�wA�|��oY�5��EnX�P#���m
'jN��򘼴h';�!��k=�0���G̓��0\@�8Bz���Ͷ�� ��B�X �i����~091���r7/s5LI>�S��q�ܞ7T�w�o��	�Gs�,cװ ��LΌ�p��c�V���VHo�v��+�w�
�����/�,�W���I4�n�1�R�*����JHW�vU{�H��q�2@
@H���2(���))�b���O�G�,����+	�Ad��+2}�a�5�����Ucz���Qnr�x�M�
$���uJ��Ϳ>fh��d刐q�gTJv�=f�{^*��Iy��H7����T����B�@"�Ā�����\�&(_.倢s���,�q-N3��㚱"�W-�aRo�?�f���3��d�l7�~fc$��:$�֊�SK�c�_�C7�L��Bz�{�h�]�Y	§X��E�`yYl�v'�I���~yښj��)��=��l2ML	���7�`b�]��a���#��`}�w`���Z�UZI@�ئE�����A�-Й�z��(��j4�=�S���'�<yq1���c�O�������E[�J��z8wfDD��g�nT���	LaP�˩����q&�%��~���(�.	�sꯝ����mT��/��Ĥ�����P������E���-}��*��L�HE:��Ne��F��T�سMqƦ�y%�.��TH��bG��139Hrp��?ۄ�%X�����RE�i{!-bG�mp�g5ԸA��"z���y=�J�������ఘ*�E�`
�j��B�������X�auH���x8�^����2�؎Kִ-\|;,�۸���d+m�ü����j+#T1�rb�ImB�5�w��������;���Cߩ�0\�i�K�^�I1$��&�����~X�!e~
Ru`��:Q�q�k
W:~��^�
p*RK8`�����_���>|;�uYK,%-�5n��_ቁ��}�~-�>��6��a4iis��;�g�_z#3c5yK����y[�IHF��+�\'�IW��y���\""4a+�T^y�?N�I��qTt6<\I����,� S+�31�8�kat}S�_���v�>�xN����	��0 �T���Bz������ҷ_����Mg�9�3�l�'<J@�aɱ����L%���=V�\盟�EN��d����䐇z*���c��(�z�|eyFC�^�y9�I���{=bN���;�Ќ �>�y=`�� �y�H�{����tR�xUܹ�b�.�C�� u`(?ں
<�B�-�l*�Zj���d��r�[�/����2b;��M��5�5;�2��R�b������R�5�����=�_���M�/�!jF�l�dU���i�*�Qqv�U��U�"}{d8_5 �nx�%���g)3v�	�n�Sae�z���2��1���k�&����g��3]reK���.j�f�N�t�6���(� ��ǆP��N׭�<o D�C��G���s�@8	��C� I�8�<s�;xBJ�]�[zx�;s�
%�%|�7%����f��B�s��Ph�߹1c�i'�,��vQ�k�0��/l�o�!��v��bb�����!�W�zQ����xWr��D�$�r���HfQJGM��1O�b_$���@wi蘡7�����aK@ג�����EB������A�ɣ -�)O����yFf���{��K���R�`}O"��cu��A	��K��\�FS��~�Q'��O���`�n�0�QG}�.��$�a!+9#/k���|=(�h<GT4��s/�yŅ�)J+r��&���u����Clٙ��g����?�������F�O�t�������8x��	�?C����Sd2v1���v�0�鏏��A������g�鿹��x�
='�I�>��Ól*�����#LA3b�q͖�V�p�`�k�q�/�>^w_���5������������gBi��ƞ�CE5����R��GÀo�[��}�!:e�pIi�[�V�F��yQ��.��paDj?[��W49��|A �I�2(���:����4k��#��!�YU����N��I���;~G������S��x���2o��t��y#�0C+-�l�c����*��A��/�Nʢ�F�l��V�`>l��&
��Z��=
�2���/�jvm3Ƭ*:������@���QD:T{TIG\�F�.1� �����?c�k@�e��-�e��F
�|ᎈVp��b+U9��-|�dNH?�M����*�2��N����+'9��ҷ1�\�
ߥ|���&���:���x�ő|���y�b��Tk�+����Ɔ`gC��እYr��O�q�H&DF�p�)�C��Gm?J�����%�1�]|�0�s��^���P��t0���\�������-���h��D����BQز��B��RM���$U��Z�=�e�����o�y%G��p�!�ֈ.k�c*�b��}�����o�ϊ����-]p^�m���=����^���rs��:s�6X��!�E@,�E�Z���Qn���57د�oxӑ�ƍ=��������X�L^������8lI����.�P�;ӰMb1���9<3a����1)c��<�M`ByS�Y/Z:�D���3�x�"���O�O�;�����/�p;�1��=�� }ҹ�n��٬ÿn������⹉q-FBw�����,�d�@'z�p�4�~�f��=��{qN����Rr�~����1j2�
�. �>�r?5yR>ˇ�ȵ�R�dʘ���
�ή;��8]R�&ݴ�į4Ej�����v䥶������sh<+��N�rW��#Q��$2������ZO�7�+�k�"��)� P���n`��Kt���{uP;���^7k,7�,�:"5��f�0:۩���k��֦��J��19@�H��Θ��� �Q-��"~�_����.��Py/2���4iUlN��1*����95}��h��/�l8��W�_D8ju��L����b�i�_.f�%l�K�7�RU�����X���g���-Av`��^d���;��M�&���
�x������飳���F�uA�Y]r��㡙B�j &&sͬE�Ib��c���Lƨ��T�3T$�����[�ןV���΁��IX�o���E�;Q��;;�.^�A�fP�P���>��^�a#�Z���/Z]�^�ѝs�9�'U�_�R�l������!�tz]w�{������qNMFaT18�"�i�w��6W�A���kJ|6@�� -��gQϾ,]����C�㜡�41|Q��>4����aи�M��Wvn�߫��8���:�����e/E�"w�s�|�6�n�e����3QgV�J{xB$i�
�q���e���j�o��yR�]��v���s�pT��K�t7_�^����c-r��<��DXo�$��A�R�HG�Z���.i�+?�y���A���1����wr`]6�)�rI�-�I���U��]\,��uϑۖWR
�ϧ� ��7$f�@T��k�9m$�{�$�l?[�;�=���hgҏɻ`!�k���3؇���.�P���L;q��%���R~�|�����~�����!�d��Rѝ���Ey��?ݜ�s+���/��YzBJ�K�����*6�;m7d�g;t�V���ɍL��cb8E�.X4�?g��P4+�� �(Uڞ�eK��^�<ۛ��� ��\4v:iY��-�q�v��kY�d�6"ǝZ�����k�z�Ԓa����qf�	�̜媑9� �*�5ep��-Ĵn���
���|��m��3Z����(m��K����B�]�$ј:�_�rvB+��4( RQaD+x�w����Y�D%3��U$�I�j�Ih����]� �B�e�v���M�0Jb\-!�ޛ���3c���?>��	��Y�BՍwp�Nq%��
Xͱ�����d���;�����qx��� v�U1O�zg�3���-�'6���h��F���#���P��&j/��w|o[@,Ru�v����J�S?��n墋|�4~ �A3շ�W�b�g��L�%��Ț�����xޘ�:J�%�$/�C � $������F)'&�ȅ�0��QF*�Nf h
�N����ʙ1��5����۱;���T쥬�P�~�<8�7y�P��:�� �ܟs�"��D��A� EڈxB���X�ӛ{aao�J,�@ۊ�ٹ>/e��Zn�7=y���
�G.?�	S��SM�Ga���m)���n	
�-BcC�\��Cv>F[�5V��Sr+�,���J�3�>��w�U7j���_u��:��Y�)�ȥ#��ሂg���q9�N��{؛�l[�Y/���S�~��<E�H������~����$F�M�s��O���v���ۜT��� ��>�e�!4
9��q��N��F�WM�c�Ƶ�
o�qD��N�Hn�����H6D,U��Hw�(Y�;H��)nV��L�rw7�EՆ+�t�&PMN����]˄��WMi��X
�ĎCN҈��-h.�-]2c���{M�=�'î:�Ac<k'��b
�I�Pa� s�@*�a�_B�Q��K�5�ȆV�� w��V��<���]5�kp" F���(�M�U<o��g��\5�� ��z��Wn3`�ޏ���&]�2e�Tߺ)o�\" �6~�Ѵ�_���͘���OL*��W���M,G��`����mШg�2P��S�GL/�[�z�DL��^"+���L����e��bۅ;�(}���b�'�2)�Z�_��L��虎*%ru�6��R�j���Z�ð���e���#���W��8;���ј�]Aަ�w�?�Bs���y;ꦤ ����L�ѓ����,��aw��6�_�a����T�xmw���_�ɓl�S�s}�I���i�J�t�J�\Et8�2�"⏓;��	�e��Vf.^��6؛-9e��bs�jJ!:�%lWi�Z��	+� ��=g߆P���P����$P��z�+��i��$7��	���_H�̶�o�:�B�M�3Jh���U>��at��*��oo��I�8��l�ۛ��g���%k��X��1 �h"�@6��|�W`��-Op�K��H'(�х���me]��l֟7zZ����/]���
1-�������w�������؟�7i 
��՘=S���qtf�l]�h7�Q�9����%=������:�>/٫�~<#!�`y:6IF�AJ�� �ʟ礄��1}�Xa ��4hI{(.���!H�,͂��%70��t��*�&�M�rzG�� �;�@�	 _`��r�d�}�Eg�$�.��FT��c��j�v�Ǆ�����͌�t��>;U�{`�ȉ��|]��g�
m$�f��;������.y`#b�0tA��#~_���՝��s�h�qy侳g9���l9�Q.Mz���Jf$�T]CUA,�QU���@$���?��C���R�,�+2\>E�MU�0O�q:_���剆�m�[J��oi���;g�J0"�L�ָuD�wX�p/��(��Tscy��q���V���|��\���@���������d+�5/*3u2�d��9�R�@%d�V�i�H���A���ר�ωS5+�bC|Q�]��V��_��l�YRļ�
��Y���g��{�Q%Yi�-�o�:����f�s�W���7h�W5�"v��V(�Ɵ��
Ϲ��s��6m	&��@�r��`��h��73qȳx�xs�ٖl���(v�av�gա�Z�H��B��fW,j[a����+5���oJ�;hN�c`��H�:���S4h��o��.Y�9�A`:�!~�2+��Ƚ���<ƴB�/#*8�e\F|o�	�L��|������N�Ts�0�bp����	
2{5�&�!���)�|�<o"eXZ�I�4�/Y��y~�vYea�����h=+�K_+�1�l=]J,�ɤҎ�V>���~��6�Ԕ���")�?&0X�A!v$��fhp'P%60��}H-:w�+�w=Z{�����ޒjhaC�j7���N�R{uK�%ܸ�6x�#s�тN|R�k��Q~������&�A5�pčQ/΀�=j�P�W$+M����.��44��ɅG��A��Wg骟D�hN��Ꮋקё%ee
B�p��� @�
j05����qqe�Ģ���_�.�J-�>�T��a7<NZ��2}j�i���˒~��
`����8�!��^#I���^n&lvF;5�.}�l\>�m[�1��D��=n��"K��(��Y��f�h�Ć�*U�uk��؁y��ie;��2D/���8o��	�.`�߆S��ϫ�x��'��ױ����4X��@<��'�����HE���p����K��?ʱX�ҍs�9��E�g&x)�U��B���q`�N��Y�ro��*����-��Җ��t��[^�jRBFjP��/�<�=6*�j`H��=�f	t#���=	>U7�k�W6�r�D�z�N��Eo�t0?�Ôm
�B22Y��o-��`W9�R��(�(�8Yf_����`ӟ�ٱ���@h&x�<�҇���TG=������skb�0��=��1��}/���a`�\Y�嵎E�P�b[�X���H�29E�ut܏ ,�9��_g�����tW�g���z^���E�V��i���J~R��� ��F·��^P�Ӈ����35�LxJô�Ǚ�$y�ݵ��}��$�5����3�f*���&��]���J���)��-�����6N��W����3�:�����T�Ա�Bog��P���l�yR��Ҷ8�#�V��%����֠��9%G���4�oO�� m),v͚�o#�����6�Bn4,�#ø��&Ր�){�d��6�&A߈�8���;�n&����[�*jƧ@k��}�O��Y�ْ	$R�Ɛ3�E<�p�_ZBm�]A�n�h�Qc( �᳤P��<�@���a��� �pp�F�ܤ��IkK��mʝ�X�xc�X�%w����aSu�µ�󦌁����i�פ�x�<� ���Od�-��*i�B��,n���^����bG�(�j�P�:�[Pp�q���H���7��V���{�q+췇�r�1xkdE��h�Bh�d|Xԏ�����*q�N�m��[��"��_���u+��-o�>�P������ŧ�G��� UN��"]=@����)���ǵ3ձ�@����bQ�����v�)����Z\�(����]�����vݓ���ڽ=�~�]�S��nrvj	+�l���Jo�=�<�v��>�i�W����۽��@+�wb�$a7�=��w�W�:����a��vG5������?�~Kx�q��F	+m�<�7D��M���G/��� �pv��d�oC�qk�T:Q�q�fi&9��x��Wj���}��q��Y�M®�߫�~x,�w�x�@kP���ؔN؈��JZ<t�)P�dS�t&(1���b�c��S�G�2x)�"��݅�f+�G��յ�bu��*�*Z���Y���G`W�[y��՞��H����ƙ���k#��7�10�DF����M�	�3�;`�b~5� �y�u�v=>�p�.H�uŧ�Ad�N�E��C�9�J�\�.�ZE�츳��~��/ �gn������+mz��׌~�d�q���~��-�����]����\��,�����%U If7Ow�2�Q]_�1��1��-��.ϠWI�md͈kH,"�a�tܪ,ue�-�С�"��Ǒ�5??��Lɨqk഑���7Ll����7�'�'llX	VRj��-��%z�b��"��蓫��)�(�B͸W������v�Uj�ꬓ�4����6Jv���!˖�0c�ru �B���+H��q�0�Y��v����EϨ9l�i�:����7![Ӳu�h�1d;0���OEĚHC���XyB(f��z6�����ɉ���(�����*Ra�~���׀7�i�Ը��-��飾@�L���m1ll\�{�,˦�Wf�y<�u�W���b�N�~ޥ@FV�6|X&�V��Y�@��q���� ��5�W�p�F�e�\`�~�m_��\��`�Z�{�B.���E�E�׺v� 3�H�2�Ľ�َ����WJQ~�M�ٚ~aq��B��
צ
��D/=$���	���%?��E4OQ�Hb�z��qxԇ��wq ����_n�k�[n�p:��@+!�#��utz��&�if��xʒ�=?J�kJ.��/��0kPR`w,�)�{.d5��W�����[.�cge(��Y�-�X��.�����[c�G�.������6�%���Ϋu\�aeU��e}�^�?��;�/`�W�u�PG룧)�ځRLk��2��+����8)G��4`�?�-(DNp��
���L�$�;Zt�^�嘭�u!٫�L���M��.�;��n_�+�ȴ[_X�J�ךZ~B�������,����?�/t��xFU#vO�	4���-~��ph&��䒑h�fdơ��������: ��/�e'ti�vٰ�C=�
��
(0���ɪ
C�w<h;ō�O��ђ���M��O)JwԆ�)�x9�_U!L��L�`3/!	���Yp��<��B] ��y���oB�n%�%�F����{+�6�vϒZ��͉�C1���X\$��א�y�ŀ��?j�����T0��|mI�B|�W^qQsg�绤����폒�|�n��V6:/B1`X(�x��r�xH���p�4���I�Da'�����m^�T}���'�������V+#T�b$!5C._�͈�䶎�M���Y5�e�n��zw�J2kx�h���a���&`N~�_XͣC�Cxd�l���GF�"�8��O=���)X��+"��G�5I{�I�];�o�c|v�{�~�S��k���(Ҿ��Q�A|r��KX�� ���\
L��mae9�NQa�0�ҩ�Tu]ߒ3�,��Μ~l�R�̎�/�L���Oi����B$@�X�z7���j6����,��aw�oG~��w١�Xwh(@��Zy��OɊ�:z�~�y�7�v�<�]9g���~��b��T[Ṕ��7@�dF��|���ݍ<�j�i
�#��>��<ކ,��o1����k�����Д��(�3&kpj�A���s��E�Z����.���I���;�(���X"1���~gW5��J��b+�;x�g�P�������([�ϯ~Le&����r*�N�5(��I
��ꓮ��#<~�m�]v%�1b{�{ oU��S.�9�S�M����K��Ѽ�9���
�xC)��|��!5|�6(�I 
S��Ը+�q���O�L�~�G�y�h5r#Yx?�0�q��c���[����<���A��5�[�1)��PP����� �L7���!�;�]����{B��\�ڔ��&��Ǒ:�;#{�T�)���q���Сd�q)I�'J��Z�����II����$��6�X]Vh�� ��-�"���'���0TC�Y�0��E��_�R�p�=��*�����n�h]�v#CN�:-�CO��A�}&�d�'�ks
1-b�p�}��~yXl���!ۯ�1�2X,[y3�`�o��P��4�)A^��e��Q�I�?=��y�(y-T��	�A� _޾�\�4�>p��ʽ����a5���� �~��B'����L������&�ą�NV�V.��t�e���G"\��R��l�(I�Ք��s�!_'������t�L����O7��I���S�3s�Jm�]=lӰEɋs�#c��g[; ��4�_���y���������q�X�[�w�u��q��%�$�L�*.�UZ�L�N�3��^�go":��*���>g��h��^[�,� ���v�F�Q�M�oI�*�1�*�r׬�tv���0�%��{x	�	~��\��a�����J�i���f��`��8�.�- ߽��x�n�,1�����*x�x�\@/�aer�^���g�O-`#8	�e�/G6��u>P�wd�p�x�r5㞻�����b_��˲z��q����5�_�r��վA�?ȴ�pD�X�q�Ŧ�yؑ@�=Yx�.��+lHE�zW�ˌF����)��I��n"�� �X��������\�������{@���Sj��}�\�f�tx�h�&�	oB� >��ƈ{g�ݹ�C������R �S�r����f��Ϝ�6�m_Q;�w���2voc2I:��I�z�FY��Co^�Β_:*,���r��6�$tm�'�^�=�{�XGQu�k��3x**flN�mw<�~%p��f�i+�v+x�. ���-/���S��}�@�<Z*4��Ĝ7Dl�)L� �3&~�v�	Z��Kү9�"���J:0pXMv�Ag\�Ͳ��qb�E���o���}l���n)�Įp��V6q��O�vD�X�0lpǣ�O�:�_�C5�}��n��?�V�QO���[¸J�V@�Z��'�)}\�
��eO����&���I4oN�7�S��Ɛ�q�g���+�H�u�^Z���O̦
W�5q��ԝ�?�DJ�7��&�a��a��O_�zU�L�%?�����E���i�qD@C#=!A"���:S�)����S��Ldh0�q�����~�R�o�2����]�?ׄ��|��z��ֆ�c����­�C����RZ�!v��I�b"DqqpTv�~k�l^OO��C���<�G5i���ź\�	s���	lp&`z���la��������w�Yph9�;����fia���\���E��͙�.lɤ�W�%^ �m�\XJ�Ϭ�U��XVEUش+ r�OYm�r{�Ǩ0�*�
A�;gMm'؟��V����H_��^�\�'=�"2�j����.ޢc�{ʸ��(k�/��F��8_'�J���nŐ,���ˤ�"�@�U)�\�(Q�#�z�t��QB�|�R�.EA�a6gt�Zߎ�T��xzZ�j���TR�ĖG�˘wBÓD���<�ֱǟ��蒑lYA��Uy��!�*��.*�ӛS!;d���_�����X����GE�Y�
��%\]�6
1���J`�>�t��C[�1��G��c��v�8�����ehC�JKp&7"r4�k�%�OzE|.��5ĵ���r8LŭH%[G�$����$~ҍat)�e3�]m�P�
kbY҂�����!�������n�m�ӄ)�Cr,al
��<���>/FT�����<S��x��!��.��{ ����A�|��~��-��E���|gd���~b؋+��o���7��C�L�C�붤��ԋt- ǫ�C��y�娼�V��&|�(��x�(>ɻ�KY�^�\�M2�����T�/~AE�6��~�<�1y2����$�p�
9�>�'Ԩ`|�J	xB)�A�ܸ�{�ǚ������椐�SnVc�)k՜e�G�h�٨wE\�G
)�m�q���{�6<�&��`~�e�YӤ��hI[Ȕ�v���@��+%��p����hU3�_l4:w��~�c���m#� ��q�(X�!�P�U�(�6��K�_�ͬ[�����Ȝ;G#0�\%�{�M��y'�`���U�J�V�����a"���֠����
�cs"T��[�i.\ӹ�+gʜP��p�������lf���V�y�6�8R �*�T�?|V
���+�\`r=��u&＠[y��1E���V4ä*a��*�荎5o�S�CMM	n�׳!G�{'�4Ku����ܙs��F1~d[L܂l�29���)X��!h<l�,����6]�#�߱a�@/�x~��2�|�K��ZGP�R���:b�UZT����b����1b��@ I�������8��M�F$�o�%�e��I���b���g�A��,=w83+o�����?>&)n���@d7�w��%>Fn��-i����i)Ku���K��<�agR.�_�&��2�Z)Zk)�  pK��c`�;Lݒ}���*6%�c�7�ج���rA��q>�Cʏ-CTxf3h�3��5鼉�j�x�x1X�##��f�����;����*�!���pvő��Xh����V��e`�jʕi(�~��Py�Q/	���N���[�S\�e��Gٲ�Z�� ��p��{��Cʥ
�c��5sx�)�))�H������)�}�7����H\�j�,k=l<���Пn�[)S&m��>��	t����\���X�g�LC9�ྒ@��z�!W#D�'cc�o��������*㝄��c0jR�cPs�
h�џ?rׄ]KQh�ڟ��?�.��R�������^��5���*�_ߦ�h�d�|7�VmO�/�����dh���}c���0� ����bԠjbg����v�f��raG[���v�֕����7 ��1�,ftA�_/+�PkS�O��B[A��SFT�PQ�4~�iT�t��f�����5�:V�FHq�
F��?��9̟&b�ͬ@͓��R�W�03:S�����Qp*/%1�{�q������:n좹��	o����si��g�6tj�h6
�Хq�q]Cl��~v�}ק�s�X�j������-c��$���=�t�	<Ŋr�t��Z�t�Eq�,=��v�Fx�ZtR�X	����}Z�����3����ojywJ!�,�O�W��;���C�|�>�����瑛�k�	G�j�v���5Nܥ�涓@��UˮnA��V�q�E)G���B��s�tQOi}!�+T���҅�N��עt���w\������c��?��N)&�v��ee����Z�Fʐm�+�{G�S%��9GP�tE���^j�h��f�/�I�������X-9�I��^�h��Ü�#��� .��I�v5�E�!�(��������;*EԹ\�˿"����nfV2��`1��3M�C�Շ�H�JrP U+ȃ��s��}�-����l�ߚr:A�s)8@n��:������8�(�/!�!�#j�kppk�����Nt�8� liW�f�eˠ?q�xL�hu�<�
"�*��'��7�����ޣ��`Y+R{�ꜻ�4+�ǁ{0H+���*։a/7t�e]�L��gw�T�Z;�a�9��F�W�&f.D&��6D�̕inp h8�)ώ��I�[��)�J�rӡ�4u��^�d}��5:�(���C:����O�]lv�M~�v����Xq~Y	�������i�B����B��r��pm�4��-����?V<f�UD�&[nO�9`�w�{�p�IUЪq=��ɱ��XDW�q.���N�Bz�\�����s�/(��D6|��Z:�S�9Bڀ�/JerayT����F�V=[�߉��Ó�Kd��`�|a�/ۼ���jh�ϒ|]��������`c
��d`�D�S����+]�O ��\(��^�Ȟ@o_�i����i���� ����P�hn��������5�Ҷ�&�iͿx�cc���/O���	t���s��P��S���^E���ld�e�C������<~�-0^;`��}�)�Ʉ���ڈu-;�r� ���24��,�g���|���D}���N�;��\	A���%{&��`�U(��ZQ��E���Z[��=L@�.3R�Y�	�x��.T��{���i*�zMxF��r�����g�����a��ds��Eo���V�Tl�"�&v� ��Q�HϹ_X�f�'9��h�r}��ݽV1Ok]�( v�x�F��M�8��"����)��S����҅0q�'s�[f�n���J���&�s�@I�p��S喩M���t9��#�>��
B��Gl�h���P�}��#����8���*'*��W��
���|��g�0ﯙ���C帵p���V���� �U�0�bo���E�P�%�1q��Jw��Z�^q�l���詾\w�I�S�"}�p	�;|������A���1��>�NA�l��$Y\̯<�W�i�mR�g��O��ˈ�~كg���#���a�w������cY��yߣ�e��eHs(w�^2u+ϰ��c���C�"�s5�+]$���:,��.���&}����YH��M��˧��Z��X۴dV��h0�2]�$x�kQ|CN�B�Y�O��.2�T����rh��&��]I�U����J��,�e0%e��u��TXl4�#Cz�N����62�@�	��	PU��t�F��(J#�P�����
��N�D���.�t���H� M�����W*�nd���,�ͫ�<�+��m��#��鼮.^�f!4u�J>��u��n����d�e��[T�Z�P���v�M(P#��o�|a��M�?ղ�z3�*��M TL�o)&�:�f�`��-���q;��k?}Hb��(�T����N��۝�M�ۇ�Aо�����Ik=����c�н�s�����'�]�sE�9۽���h���Z��ݏ@{S���nۆ!��Xe�T u�b��e�X�ua���ՙ��]U�fCHH�F���ϒ���p��cJ��RZ!m���:�Y]��z)�p�q��T"��%u�ձ��*Z+��oҰ1~�0��D�N��W��\Y(����:O�흘�y3! ��EX�<47�YP��n$�q�Y������6;�W��s+p�G���bIN�%荕Ce��zV㐓p��ñ�s+�24zEV�4��>���� �2�9ř}�2�X$y7+�EZ04Weێ���I�)�G��a$W'��i@��Ø��O������ �wakU�F�2w*���)Mcw{ejK�Mz8B-2�t(��{]t���2Eԇ$���H����{2½��x��F��%�	�+̔N>1c#@&��^�����|1'�HC�	a����c~7���5r�}+|+e�wg̓�kF���pJ'Z�,$\t����N��p�! �M
�|#۰\���}��8�L����-�gt>/gW��Jيc��W�������|���1W������x�������wʳ�]�$��֤�d�ϟ��8OI�V��Y�K-���>{�A�of�}�]��ɲ#!]Iq�I�&̖��-���-�h:J�v��o��ɘ�1y������2���q�L���urt�m�dd�*��%�)��x�Ͱ4F���a �
xSG�(�O�h������^�j~��}�oN�$��0f���ᄉ˙�t��7~\���Z�zf~��=�d^kH���6�ڕc�߭�������Ԭ��7c��p����W�����P!�?�%Ԭ����c̴��i���b��܈�CA�Y?DK�>�_D�T�lRJ���4ךU�S�Q���ۢ����P�����r�AV��B�������#<��+��a��㰸���k��_��_�ZIo�鹩���0N��z�g�5�^b/�D����%�:�Pg#"�d�x��y���
3�'���Z���JD��@�IO�P��s��Kp.�o�YxC��-�d�r����RP�Z[������S-���a���C�Nϰc��ײ�j��a�X{�.upK����phs�����Q�z5���q�,6%_�����M�>D:Zi/p�$�]\��dEO�I7��ݭq�͉���,�Ï63�X�~{�� ��-�?�:��Eܽ	�E6>��{q�*OlNM�����%j�>���f|�Y���+�:��`0ë�>��,�ߺ�J%U��#�6�[���bD�C��4{�,�ԫpX)$�1�S�"x���|9��av���'����� j��]#q��I��|f���F+�*�X��`e�jD���ǺG��f�UF�GE��J���c[s[�(��P��}�,�[d!,y��
�v<Z+�����ܥ(~�<���I�4�i��B��yԽ�h@n�C ހ�&RsX/m(���ֻ�֍�a�h{���9	M3죺Y����H���bΨ��͆{�Ƒ��΄g�͑�-24��9�i���	�xfc�X��v�U���fR�Nc�}��֒���փZ�^������B$�*�V4V�1�7�I�-
)& �o���+kx�O�(���-���=�2���^�U��(J�Q4�橜.P*w��An��İٜ���Oi���N)6�,��n�<#L�>'�+�e?� �s���p�Op�t��3��΀�(�����r���N�i0�{
C���?%4�ݏL����Lu��F�����gZൖдC>�Q:����d�PAٝ)}����zdW�Y�z�.1���DY㋵�/)�m�ͨ�˥���;�M*���H3c�D�3_�n�Tn߸���8��W{���_{��r�������>!b�﹉����KPgP_�,�y�9�R��zhKP��nzs�ї��	 @yi���Ux����zo�(o~cPI1�{ݦ��0I�T��Ss���8DT�PŬ��C�/~��F�y���-%�o�����CKJ��Up#�p+���dG~7z�]aD�f�Ε�$Ԋ(%�snc,`	<D&�:G_�*���2����dI�L��Я��]"��࣠0h�X����t�D�<,R~鞠_ZJG�Γ#��zr7/�I&�w��s����sm֟�:6^���i�%��r펋��"��� {����i�0����\ISlCׁ����\w�*�7r���Q�O�7Ѯ��@�������Ψ���<��X�$���m䓵s�1�Q���_,�z����Ҳ(=r*m��q��75�i��$pCd�_{8M�f^����VI�~l���Cߩ �p9l[-��A�|T��!�e��'�S�����.06�B�U���ɴտҐ�����&����#���.�E*�R(�
+�\3�
��)�B_k}J�8��Xda{������u$��D�L� ����h�y{x��T<���{�&�#ud�ps�i;�K �c���`�%;z�4�A�Y�V��N�f�`�b{n��y�:0���O�jGu�k���]�q���do$���W�c������D9qL�^��:���Йb\��W��e���	���7�S�|=Ov7��BAN��!\lM�F�(n�a-s��wlR턙���u\��� �]����״��_z1T����Xa�O$���o3�J�%.����-��%bN���?$���3�
o�^���[��V�1�G��D���QOY!U����}2�+7`�>�T��6��0C��?�@Y,��e��8�i*l`���.:U,���:�`���d� P�9%�C�{�r l8ZKJ�H��ǣp{Y|�nK4����9s�"vI��%���������i��o>M�6�oߢ��x�pԸ��"�&��W�cgJ�y��E]n�P#n�&�n�b�y8�Wےuv��Cn �{�̦������΄��)�mX�i,ќ�}�iT�U�RTɅT��,V�*�*D�C{y�Fk ��&ݙ�u�oh� �<�1>�h�����*!
�%������t���#5E�s�4�Z�?�/��#�|��2�@wEa�l	9@�d>y��;��f#�;ύ�5LGe��-���<;5N��w�X�vo e�ھnj��s�4��b�צ�u�J��O�֬�� w��D�T�=R�Ǝcc;0>�9�fwIإſ��P!3�W�R�����-����n��^�&�/	դ�6��M���d������/Q�7�ft�$&�أu1�J��jv(���8��|�62�[G\7xU{����y1��9rii�����3<�<x)��O�l�X�`��j��*%(1��$(����f�,X�c���7\P3� ~��N˩.�	���]�Òz��m<�1m�R%︯�1�)�C��s�\,�D��� [7_����R�H' ��Fc�f�_�}���,@�Q�O|���M
�:���R������湨:Ӻ~��1��F���2���}� ���M̚��V�M�m������i�óB���g2�vdt������ln�Y��Ⱥ��C"N���;��F��;;�F�����)K'z9\9���e� � u�V*5�/ZC� �ݷ��Pp9A-��2�-�<�6��Lz�8�`P�zS8��K�9�� ��@� ��?�_�>�0u�`ky!���̅�q���8pBx�.w��UKbn�q6����VR�9��cg�f����R��z`A+\t.[>������`�fh��q+�ȉ�#��'��%W?� %�6����2��#o{���`��df��uZ���U\&ϟ��P�񣈮(n���:�V�'��Y���09f��<m��6��Q��caͶƃ�m��R��@F�n�I�!�px{�|�sW� ��4z�#�-�כ����!�.d�)*u,Λ�լ"
gje�B>���a�F�x"��(���׳�_��C��!Ϧ��wo��܁�(�{Ȗn3�KV�J��b�����T���{�zD:�����-"Fڽ����ėä�O��e�;��l���S���^�w#Dܦ,sĮ��>�<?Bv��� ^5���E ui�V ���CW5�0���J-�=�\[N�8#�~pN;������}fn�]&���O%��o�!�M��1��c?6i1��I����'�۶s)�,6���IST/�!����f�K����Ut] �yw�[܃�3�x���Њ��d��w��.O]����dq�r4� � +(?��GQ��|L���yf�n��Ҧ7C�eƒQ�9��@:��Nn���/<fm�����=�>@�����y��X��V���K��+*,��K�����y�D����L�bW�d�x����§��֣J�r	}� ��ij8&��Э`_E�e���Y$�ލ�C8�$lh�_�㔔k�T�wI�g8t�4F�ͻ�席k��0���g�0�9;�N!�`
<|��ѕ��(�z�Z�H5a�Z��m�r,�H̝ c�te�����ٶx�B"/���:`�z�ۤ��%��z��(B2j�������%1�u�
��#������X�xЇ61\�f:V����������z _-�	�j��?M������Ҳ����p�U�X�]~���!f���eK)�8���t�[�4a��I�����i$��R�UZ�ŕh�����P��#6����
X�t�ԖV���/`���\��,�E�	�U	��X�i�@_d'�0�;x[&pL���Ғ������=r�˾�M6(y>��e�I�1����czF�E�	���FP @5}`K~L#|ú�#�:A� �ơP4�t$or[,����4p�>v�tPe�0��݃�ur	�qN<_Rg���U�G[0l���`ѹc���kb�o±�ͤ�wɛ�m��H&_�T�V`.�䄾��ܪ��S/���2*�=��b��[	���s��@�H�q�F�א��UO{֙��a����5tE#M>Y�}n}��%w�q!��e~mqI	��@	y��b�g��fO���5g\�����s�����g��DU�wX����^sX�O��pluɃW%#5��}��̼��M��=e���T��գ��;axz����3���Iߌ?fFA��4��(�HPc;�(�K:����P�)0S�x�B,Df��Љ>�!J�sス���G1�i�u0�rNNi�����
�B4�s�HK]f�\:a�ԗ���b[�s�"h���Ѩ?Ď���U{��z�S�|PL���q�[Rӆ@�o��]�@f�0��6�o߽����uÙ��+�Dd�pU�B�m]�Xb#o�!�8M���d����f�^G㝌Ε�m-������^��[���O��/D	g��%�����e���5���aU ��qu�����Fx��O�\�,+o��5~!X�Z�B}c�'ۼe�?�d;2�ҭ0����wn�Y���.���q�����^"��{���#�~|��*���3��yu6�^��b{�Ct��]zW 4�/]u��O�����&���vb���LѶ��Lj��+L�麍��t���߆W���z���_�[ފ�M�e�֚{,ҧ���7%�O#�b�,K+���Y�V=c�A���XP{�v����1	�zQ�N���i$R+>���`�CXO�0�$uԱS,!��g�� no�-�s�����Fe�{õN���Q32*����ZKi������D?��H��%��\Щ�طW/<	Ҧ;�u�����7�O�c��_'!���m
�� ���I�qh,NI�3�і��}����W��O��s|�5�/?�VÓDD���n-n��j$�N�
�n���VmT++<<�?��i�N�q�<�S&�l���E',���4Xuٸ����P� .� <+�֚*���H*��6�f�9)L!��d���Qͅ�eg��|54[��y�m�g��l�c������NklRJ���K���ӌQA�3�s^P�=4��*� �ѧ%	2�Fý��]�:�hޚI箘?yR��ЀӜ!KP������vy�e��Ah�p��X�u���8��+�P?@� ��P�E�}������V��A��*`b%����j�`���d`�s��U	U^��ռ&I�Ɍ��>�ve׎x��V��g�&�J��|\N�l�b�>c���b�f[uG��-.����}�:4MЫ�I|�����G�+�[� ���(	3�q2����
G'���C �:���Kd�0]p�
t>� ��7�l젶�'�st+��#\�!���	u^�b*t�T+���}6ĩ��*���х�!�%���>���K�yDu����W?��\����0�T	����S�:�H}�|^r�U	,�	�mB��(,,�� h�%����䗈l��
x��^���p{vMӷ�,yƋ�Mę=�_;]B��O5����P�@��5�a�/��hVk��� [Oz���v���|��>}���S���Z`�W���`h��J,MeQ<�}>}$<��#�߬�3g������:3[�U׭�36}IX�^��z��t��{z���/߻V����]ώz�٣I9L��ճ�o��Be�(��H��\��r�G��(����,��5�]+��f<)�K�7�8R��2p+X�@=�bd�?���l�y����^2�18u��f����Y���(����8܄ЗVb�V���������'TNߟ �l�(b7��ۛV)l�7��V&�~��^3��0�M�$��q������FG_���#o�^������cl�4�g�|�Z�q��蔘rYuA�K���I����4hA*oJt�����Ĺ�83'�{pE���T˕�G��7��ں��ܓ���>�
F��MD<�f9k�~�R�7�]��4�@�J� ~D@�Z������Ř�Vj" ��o������-ЫzkP�4�	U�d�k|+�ah ��9��>��hqԀ���yg]��;������ ��/u�1�f���-����2���]��L��H}oT��L?V�2�k��ٹ��k���9����J`U�՗1�u���jӹw)���u�</%K��sX���)���99�L��ɗ��\�ԙ�2 0H�`mln�sk2w�������g��j�g�y$;��q��q��T�ͭ���&�R$�<�D�O\���%�m�K6��`l�hr�<�dl�E)�U@{O�R	�΋k�F���(L��PA�W4ٹ���M=4}l�p�L����㡩	�ɴ#n1�;�/}<7Z���3W���X~^������O
-�k�WB�Y}�$�N2&��]R�]�u����*��S�a0sY�:o>g;!�mV=�$/^Z^$g�F����d{��l~�6T��YLc&R\�ܥ�B�r�ai3���J�*"·�%<� 8`>B)�-5~��	�ѥf��oYT�Q%����ή�u��jq��S���zx\3c���e@�mt�m�;"���<�gA&^ݫPq׉�e?m�lCz���Kƙ�B�ϳ�9���(�>�f|��N�*��2�r�#�����z,��ң'|�l���n�%���~A­�\LX�&��d��g,g����C�#��_7�Ӆ�4�o�=O�⃥)��?9ڜ��b�F7 *s�Guက�d�/I2���fc5��0���1�d�ox~���h��@g(-����26��cz�T�%���4�ׇ��`���f�9���@H���R �nGk1�j?dHQ�H������D�	<��� =�yZ�0� ��/��W�Δ���,���gB�݉ۦ� �d$ ��D��ѱ}�>�֏Kݧ[��KP��F������0�����a6�F�
[�V���4�ᆋ���UL")��	C���\��7@H�dy>�b��J�3�U�5`����\�95�F��䫡S
ԉ��B�8ҡ��V-�	��k�o���tp�}����v^|��ʚ���2�4;���=o���iб��T���x��D��u�C�E�����c�u��|'�菞B����('-NV�d�<�@}�Ka�oZ�S�H���������sO�w���p���h�����;��$�U�O��vߪ��齰�����&�mH�k̟㢖xn�X����2��#0Q�(�؄}x�d+�id/gIMy��Fs�����I��f:�(�\x&N��=n�$^�$56DQp�]�kx�����-1(��&`._�������~�脍�Qɠ>e�ێ��G�Ւ֡oB��K�4�����` 7i�<��}!p��*Ep�v��8@
̛�9-�U�����!��q멇E��܁W"��et�6%2�(���z����i�c���o��p�n�;;^<������ۉ2�ܸ�C��c_�;��J���aH�F�2���Vcd��i�~!(��ݰpb-�xI%�����L!����s��L�ټM��6$�L!ˮ[��kwCw�!p�"UJQ�ī�Or$�[`�1����"�M�:����$V�Ō�����c����a`V�,�a�\A\� �GirҤ��M���	e�1|8\]V�JCm�wݑr��n?�����o ����&�iH$���9S��'�����%�{�nP�㳃WP�Cx�%���7�ӣ����H5c;o|��I��NP��'�W��^_I�]R=�x�<���V���1����oe\���=	`�O�#&z�_pr3�������z���OJ&���g߮n�te����Lhg���]ST��DM��
d��������8#DN��x�Xv.�@�9�o�A5�!��MXP�V��O:&��d��2�3H5`�%B������I+h�_ѻc5������
~��W�S��I`T����3mc�+����	&��`��%a���η8�鰭�W$x���xU�u�3��1W*��ݠ!|D����m@nrK`�	��ϛgp!1̱)�0im�ٞ��DV���?�2�2?����i ��)��i��0��Q�i���d�&�v���Oۅ��j��M�P�`����w�`PsdM�H!>2���,��1aR ��y[��o⟞����=��B��Y��Z(���=߫���&�����[ǝ~��w`��٣W�kS]�d82�o�{Ǖ1:��R؀�{�༈��_���;ԅ��O�=',��5�P�+���Ez��l^	ې�����G��ăG�\ۥ@�z��9��z��_����,�+��oT�E�9]�l7:�9�P&�w�Z; �8\��1�S�8�[�6~>q�kP_�vH�ZX�h�F*�Į����\�,�3z`�(j��8'�L�iU.S�0Sf���%f�#O�X��=���Ͽ�<�@��\"؊8cm/�X��\9��=6�"�j'Ƃm��A�����̒�X�I�<��k-��va����q�����(u4�o"(�b��@��+9�y@�q6��0o?��C�y������ ���Ϲ�UC������c��=wY�1/x!�͸��c�������7��Ch��'c(u��&��Y��9����Op鹆2��͑��K��w{r�^Y@���4�� J���)گ�GOeg�}c�]q�"�X*�W�)�������]��"�P[����ͪ,�ې�O_~��U�ȩ\`���A��K�������N٘���1�Bng&��6Q J��FP����3(N��̣M�$��)j��}!����2���\�?����]Iq����[@C-z�Ebf5+61�4NJ���/%�}��+�S]�ئvK��6#f�j�f���R��q��"�@)Y�s�r��K�"K]��kTE��p�������d�2���Ǵ~ҔSJԗ�����9H1���/�L����9$x�jx.���	?����rx-��s0��g�_���"�`!Gc�ٓ�ɥ{����E�bOGjK��si�tC2�tS��������?�G�����ֵ��ZX��W6�i{�58��@�V��!�4�L���O�����&��/���="_I�t�4�4t	p���Z�bgb��G��	��j��:\>s�e#�D� � 3��s�Ը,a��Dk����ib¹�J	��un���Uu�	Q6�Z��q�2XCl�b��$V]ul
�$-k��#2�u
G�q�&� ��OW�ǻ��z����<+��6���Lq>mzH�Zϵ)˞c2�7�A�������;��d2�8C����s�e���<8�Π�BY���)�(|JFu��J�!�@iv�W��ՃM*B$I���ܬ�LN`�D���<�j�ڟ'hw8��ݯ��_�3n�
a�ҍv���v��3:���"IYQ���Ȉ����g|��W��G�?��ouM'�G@$1��O�ȅU��.I��k��H+�F5N�=���ms�� (�|��>}�0���x�7�U�x��_$��U5IL#KEN,��G�)�R��,˦���v�fr������c��8 c�-��K����C���xf����X�-�:�WEʣ@¨vp���tȁ!��;���4���1�Z��V�PS�"q����ϛ������u����޵%_AJ��e���1�����̀��:G�Y8m���aߪ��
6��"��=��z$�����S%������.����\��"���X|D���&LF��������jb��+Oq�?�(84��r��Ք�-j��ct�!��/�t��τ�u�Ń#�ݿ��g���	(�ƧH��f����hJ��G�/�J���6�������4�G4�^��L��v��p�>����~��/f��q��J�v�����@~�Q���_�`�<l�ɍn\y��!��DM�C[�%Q�q��a5Z� ��` ������uZ^Z�ew ��*!(�(�oυ��oR�`I�R7V�^g�Q�Uo��}�\���������xk�����x���X��'޳���k8w���9�?՜�j���\���D!�r30�rA����e$�Iy�ή���b�c����89y�L�	J�^��]������,�Ơ��� ��afI���\e �����a������D-�6wٗG֖���S�,!d[/��dÔ,�.��+�(��ʠ�ɛu�J'�I����S�q��<�ߧP"�T�X� ����P��`)�	;mQ9y,�{֏�휇{]"��m�O]��/����U��Ӽ��`�j�Xn`;Tˁš�T�!���i���1?w��fnb%X%��^UᔏyoK�d���p��Y�U��r��S%�T�E�`>Pգ�ؽ,��a�\!�,Hä�$�(�@��v�=�Yr�@�o�:f�����
�[���(D�
��r|�W����e\Ĳ�짳М{8-��ew��t�U�\M���b�GR�a�^�k�:��A'�n�<}j��f������L#�`N2^AǨ�2Ŗ7O����%i����&5ҕz��GRS�������4��r��Ȟ,��xFx}F�2B�Qs��
�IC�yzӒ���dx�$e����F���^�?�;��i����} ��I����ɖ����1ܣpշ�����f+_q��7ǘq��c�oB��^��8F�g��<�\J��7H�$����4�������	�c营"����˔�}X��=��2�(��RXҾ4	�n��P��nɔFaL�i�g��1�z��Yq���0iyꅨ}r#���n�s� 7�{8��nR1'�G�dv�x����y�w9�v�-�1��ȭ�V{?���Q'⿰MS���h��mrؗ�I��b/"[k��U��u?�	X6�vx̛�H�0�FӪ�;ft�e�J#��]�6n5�%	Di1�f=[8.�-3EUV�|�#HI�p9�\���U����ڊ�Y5�K�x*�Uv�s�̳�	v�"��M�?1��y�_n�hjJC<`l���G�{}jyT��I��9X]�N��Q_�� �LvyB�+��X��;
�s���Z�A�+/�W�o�6���q�d��'��?wX��D�C�4��ꎷO����mN��au<[-�tȥ�4o*&,�ZpF���x�������R�~�Z�w�K;&I��Ϟ�ȇL�xڙ�F�������<a7|,�Q>�\R`U�x,�C�e���4�K�!H��M��xE�^�,�E\ɾ��S�H�uė�t(;�G����t�O]OGn[���$��&� P2;v��9U�f��y�A"��g�Tr�j��[ƃ�\S��@���A��}�����2h�+�/~�� �/���9��{_���͙�AʖO?�����1��ʉN�ӡ���1=���D�ɉ���$�X|6��ŵf(S1�������`;��:�tU_g�	N2����
�.؜4,�H}O�����bI��!.�//�~}KI�S[$!����c��=d�(�E�D�C�P7	{�iӴh>��7�@��������D���z���c�Y<�X˴��.�-����^��ʰa)��z�.�7�e��.����aX�Y�1T�iת́��^5��*��mZ�C�5����	����&١���:��KU���h
^����5���`%{�2hJ�񡦖�"���Z
�M@a�^�X���<۪�j�6�2a;L��݊Qw� .]�����.�+����t�4�s/K�+��d����(օN�������E�0��K�ģ#�6\��5�gT��C�+��t!�'f����s"�7��#j�W!&VN������ӋY����i��c�nl�ՊX����g5�^.���:bιw�9#Ũ��QrJ5��d��);%�s�q�A7l5�۔�jt(�m ��
Y�r���~�,Ӧ�3q.2B���v�F�r�V�a��@�3�j���������,z����x�*�Zʳ<�B;�*r��R�K��A�e��֫��mj�r�:�S�A�L�=}��]4.�ꮬ�9�����[#��F*���/�W?���ubj�y��a�s���p% �ª�Z�Lbf��(��]��s��ϯ~X�o���!؂��?>��D2MW����Mh����>��$�H�S6�,XE�$��H)�9�a�5tu�dB��$h�a]N�-[A��Him���V%�!�X�K�����F��?8�$_�b�S�׵� �R�Y>x>��5����z��)��z�\�����w�T�̶ˠy���JƩ�����
T�.`V�\��y>���GvZWå������Q|�w����L .���� "`�kqNt`.Y�	5>��h��jz�)�ռQ�֫q|�Yg#�,@hF�+���\L���Zܘ�Y�l5o[.N���5��n{,V��h|s�	&_!ä۾H�2����3Z��,��;5a����Pd4>�k���L(-!��,ǂ2��X-�F&|t���Ro���|�s#�	
H;ΙD��[�t�?�L�qd
y�e|�@Լ,4��&l�=G���%�/T��f���8�����H�ˬ��lHT[�V���&F�p�,�j��4��@�-���E$��E���e� �/|tC��b��7�T�?��S
'ς�
d���4&_��:^�ӫ��˾�{F N*����|��0�OlǨ)��wZ�[Z�ʒ��V�B��9�t*����M�W�0\2���◮!����E�%�p�G�����Y49H���W��F#k�2t���A}r�{�-���LGi��j�x�Q�C-1Jlr�A�|	�w�	�Z��އQ�{Ǯb<u�uU?΄^E2�{^�����R���4݆Ed�o�;���~�;��\��lLE�ƒ�������p�fƽ.����]f&YNN�0D�csӍ�2}@�ZH+܈1��`2����]�n.����<%���n�	�?J�Z���� �E]��:��t�l����Z���m�D� ��l�EpY00&v��)�I$�
�{��~0&�~����SY�RW;�z>���v.�>tfW3/�S�GB���� ��2�r#S[����YkT���j>O�$�-od���/tC�\Wj~- �2��Z���f�3У"V��F�R�ӦOĮ]�Ü�f���ժ�DO�Ǆ<tUja�P��U'J8H����ed�
��0�X�+i�Z�"O����԰�z ��ß�����Q'�����YF����y��=Y?�KKaPH��h��5�A"Qj!H��:g�Ei��[�3�E�{|#�:���W�4�X/�P9)�O��)Z0�A�X�U<��v�#)8�߃Jѷ���B.�c�D!*j$�U����:%	�9Q��*ݹiH�(B�o?�<�}�������A�r8���^�\ZՏ:�C|Z}���x#?-�0ƸX� ~k{SR�t���l���E��QAn��n��|ϣ�����B Ω\S��������»�fYivE���L��jvM�N�u�b�^,�"��5�FϢC;���d����l��Z�
֐�����@3g/1���}��β�u���4���Eq���3�RI���-�/p�JZҍ�Hu�e"����I�Nl���!}��n������f"aa�rF6	20e"g)P�e�g��)9Ŀ���?��ܪ���}�-Yf�|�x��ⴚ�(�l��Pq0;����[W��G�ԝeU��h��[|C�v2G���v|v��fqX	�"�9)����D'����W���E�{���d�TN�5P8��+kg[8T&��.�e���8&J-U6'��@��o;y��:�i�4�Iv�>�YO�<��N/���糤�J�W����x��9a�ǝ�N�l�Э�����c�Osvll/�k	?�<> ��#��rxQⲯ!:!,���'5��I��hO�dV0tJu�&���n��u�I�`m�J6�ʶ���C�ĺUKm�L�2U%x}���	b����������&U9xh9��<�'?<G�q�ꅖ{us{p]?E��-I?ʄ��G�����;^-��N$�F1Q�h��hŏ;`�.�g���%��x�!u�>��{�6�m��P��>$���Z8`,jo�����]�ǻ���gh77��|���`�3n��� H�)�'줘H�Լ��@�\CT
����jj���٫�!�/8[���Q(LW�(#;( r 	!w�\�yDD���\�I�[��ZR�J�ns2쿁������@����Cب�a�́Ȝ88����X���!�kV\�ҿ��kRFi��*u��s��;�'���M�3[����";��u��x�!	�t�^�q1N&ח����E;z�m<	��h�b�,���b�gF�쭊8��g��A�!U��3�*
���|��'맔�܇�t>2����[$R�?�U�eF�O��H�i���m��"�'1.��XCG��v�)�x���H,���V ч[6�y�E�������2�(E߫om�mA�c͠��-��#ۮ���PS�����CQQ����LG.�I@ۂ�wO4����u���&+\�x���������4u�Fp\�}
�I�]���=LO�k� 
ܫw(K����L8����z��35��,A7�,}���xR<������c�̪m��8��[�5�? Q�cܦ����$�cx:��A���C�7�н�eh���d��MI'j�@��4���"����v!���"�P��r���x���no���-�8 8�PO���� �*:m��zn�6���<��j����᠂?��� �o���A�p���~>a㌖��/`��1OE��I\�@�>^zQ���Nfǿ"+��1sgRz�r����5e_0��䳞Q����6j)�c����sv!��Ѓw!�b���N:�%�H�O6ѡ��%&@ho�;\6��]9�5�mFT�k:M��N�;N�뺩��m7�?'�p����&�3e���p��II�V$�����-A(t�b�	S�Q���[%HT��jH��e�����L_��?Pqp �E�TD�8!�>�&&d�s%c����Zh�8%��<��b%��l�r��Q���f��i��!��jD�O��T�@�^�wJ=��0+���2�Ύ�=E������O4����0f�M�O@�����{�o2��>baK�u-�\�
2O\-���T����LQ�?U2T��ro}$il�s
���@iu��۟�&�Z�@�}��C��%��i/��a��6�������~3y|U}%�s��V+j�_X��q��)����I7@P���9�&�e�m�ޓ����6��Rqfo�S�Tx�2��{���̓i���74[��;����h��fes:U��B�%��e3�>�3~×���๟ƹ�_��p�)��k���Dٺ�׃�b���'�G莬��_�ş�y���q����#� �a*u���sb<r�Pڿp��*����}���l�݆��i�~X�u����m��%��_t�Bɞ�chϙ���a��_�n�G?X��w��Ģ��5��0�Rp���ͽ�\��[��)'�P��9���b}����ps����<1܈��)]���ia�4v��d��s}$p��M���(�1�vb1�_�A1��vl�ӏԔ��|cC��7|��n� �?��ٵ�_%��,�O1oȬ�?��+��g3�%H�3!���$#k���&�d,��ĺV�nc�`�ƪn#��F����\^�9|����6����������u���Ƨ[S^�7�w��F��)��L�ڀ�mNϽ��ż-m����p ף�j?:��8�?��J���YgL@��5�cF�h!3����UB��q����ӎ6x�SP6d ��oG�xߵfj��5����)F���#�f��w#qQY"�6��g����M�a�A۟7DB0��hI�s\�K��������N({I��4��جX�{�T�=��c-�,�]�G�j�XcU�jϥ��6{��5p~��5��*�2O��Y���P��|�����%�J���d~�`)�|e�<��пd�ь�Z��C�Y4/LJ��%��8@�X-����a�b� ��c-^!?)U"�c�]HV7m8K��(1}Љ=�Z!��,l���ưI��M����E<���D	��B3\�_,�ݚ�ѐ����V�L�(aI��|)S�Ya���&�~@��(���s�
���;#;o��W�(��g���~�3��I|����h��D��Н�y>@o�?��!i$M���BQ�j��ĿuE�wAoC̶����g�<ۖp[�C��ƥ�J��@|�D�k�E�+R��AOS��.eUf���b��!2��Dv��
�]d.�-I��F��癣�噘p�f���2��C��y��*�/���i�K7d��ٻed����QY��SI����v��u��UE���
�4'_E=9���ܖW"0�A���Ѷ�����0qzhVH/���T�C��|C	���##��U��&��, �vLw1�Ss-���Lv5.4��%#��A�eܫ��IjmFmi�wV�`9�yZ���R��o�h��e�o��(�~���=�6�&��<i.x��1���J`�|ӕ���D��r{T%� ꭛�Q�w���qPZ;3�D�tyEpo�L6�!�
˫�w��w춧<����J�U��H�ǿ�� �tQse�Z��� �[ǳ��%J�7(�!��� Q<]w.�<�!k��(I��X����ź?y����EpR�2Z2��e�����\TӐ�ݠ_#^��ڨ Ǻ�ϸ6�0vdըTA�OĤ�66�V����+���tb0<��v�{���m���X�8i��w�f\�Gj͌�Q�/�z�] I�.�/4����b�y�ݢ��rH��	����0� 35l^������z�a�����iNM��nH�������q�zYj�a�N���ߙqs�Cc�F����}6{3hS�Ca����T�8��G���H���qpw��M�ͦ�R,�*m9�2U%�B�ϖȭ����#�m+ܖJ���p�O@�� "�l��r�^J��k2{��_�',��Sw\�{d!Q�@��x�;㜏�����k)���[[]��|�A�=�T{'�%��M?4�w��g��֡�2��= IE�ݟ\v`Q��yFZ�]���/�hBz��@8Hj�J&V[O�li�x�p�h�Z�W�E`x2C��'��(�b��\@C6�HZ�i��W��-�\�c�,9��eP1'�|����Nͬdj��<X*
W"n5&�{�+������d�$-Jh-�a�).���U��v
]KIP�����!�����2B<�n��n_��mj�豟�^HxB5iI_�?`�w�	���]<s��2�8��YS�$Ǯ����nph��nh�Y�.3�O_�toL��07cK�옞���a��>@�>��0�lQz�/<�d]�G��d?�/�Ӛ^�� ���Aw����"=qH���c�����m;�
H�Y�n�|�y;���]�NÕ���FF�1��L�` ��s��4��:{�nz�F]4��L�_0ꕁa?
�w
g�&�1f��n��l�M�~�	ܫnI3���Rw3
��<��P:wS�.׊+'cf�P��Ohz@��|�:�dO|�z��r�+*wC�� n�2f>�L[�+�_̴]\�zHqZ7dC�����a�Y��^��0s��:�E�����O�1Nq~���ڨS�U�Iyt�\�V�@���[fw���6_�$�$|J�={�S�3�G�tz�����g�e����0+��.�%=$��&Ḛ�uE�R�O�ۡD��a����!���v���~���T�ڱ�$��R�Q.]b�MQ@% ~5?h6�L4��|\�?e�۳��3m�t�����$"i�tG��]B�� �]%Xw�k���@ܑ���f1��[��M�������yB��'���@��#� �e�d��3鱲����	�h�O� ���wb&����%?dl�*jE���H��7�G�и�"	������4p�����Ó���<d@ur���ҳ��=֗�Tr}Tx7ULF�1 �i��+�n�����𑝤�tV&
7˜��r���
27�=���_\�Ḣ�2-�,��+e�e���/�aE>����]K�;{6~Q��d�e�i!,��5�Cι���f�v���$�`�;���;�Q��.�/��g�X�����v�k�
*��У�<�js����� )Sc7}���+If��3�%�$r3���=�g�._��2�
� t�+?�����B�)�h�fF�11�87@_�)e���	�/�vZ�����L,C0g�R�C���gu6[4��!��I�O�(����.�#��\��w�T���?