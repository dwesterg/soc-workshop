��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�Ǖ��[�K�S�%J�L�7�@qM��M[�ߎ(��.��8�M,�t�e�r����n�9>���E�Fjo��g����ȋ��T���\H|%-���?"ӎ_؝dwƺq��[��7'��P�t!G�3R��Ϻ�<���j�L_g�z�ݝJ7�ATD�cs�⦼CXXjي�v*��Y�n�"���P9����E�<��d��Q��7{[E-ý0������^,K��i1�]�q��:�(��U����^�d��)�i�݁`���"�~��D(qav�buZʍ��@���8Y�1�v�)�����������N��*o���w �w��y��P>���'^^9����fz�<�
�??�+�{����E��-�g��������)�2UJR�x�z_����;����b��~�ڴ!��n:�Ո?6��rZ�g�i�b���빛ѳ.���p�:��p{�0��̈ʵ���SCF�݌������:rK�j���up���NȲ
kn���B[�#���_.�"����H���o4�0r�����y뎗+$6�@k�֨�D�V�w��*Y�"�v%,�f�^o+�+��m�Ql�EB߶�e�� ��G��Nq�g�w9Wnr�,'7��W�]v�7xkNӞXs)C�o���v�]"+{�J�f	U�e�t��f��iN�;RX9����|{+�1
;�-1��`gxz��j)l�Vy:R69��≰�=�B#���L2E,;J�˫~��[� _SCU���S0P�UP��;k�b�
�������2Ty�?��aNmZ˨���D*\}!Yh�Q$���B�!���;��g�N�=[���Vkhh�O���9�(')���k�v�ߏIB��ĭ�j-N�oʶ|~<���X �k^�(��E��?�d��`p��μ�{f��Y+�T�U'X�5y;�a��Z{i?\�5�/�z'\DՈ�e�3��J�r�Vz���`��*�WY��ؓ�+���t��w�Y#�XM�{�\��)�	�i]�?�S��CA����>��o�R1.�μ���}�b�!����Erj�%TP듸�l��<���>���hS��#{�m��w�Gj��9F�����u2�/U ����#�s�.Znl:�����y�^��Ɣ���i�%���R��Ҏ1{.W+Q�_V<�Qńy%���+F� �{��u��-�v.���?�����Y����ԑ�i���6.	߯����z$`�+=A�+��_M��!��1����"�\�	�4C�7S_o���L�g����>��`F�y`1Zw��)-4}n�hj)���r���Q?{�c�ܡ�T�����´��u����$C`��@����_�
{��t߹�T�DQ�|P��8�>�M���1�b���hU��),w���τ�JD�,p�{�ySya����4��FG��hQ�F糀�\�
�>�)m�5�}�^MU����C '�����^Rgi��=&em~�dQ�S�5�m��N9zI뽣��O�[�1&O�l��ҳ��j�FK�
�1��.�����^$:=�U���E��;x/9]��4_N�g~H�g�Z��U�7�*���t�QH���tȿ��1�
�E��)�RT�W�r�� ��t�l��]h0�g��ȍ�U��"�r,��n��(��ި_��1+m���8k�݈��k�Hf��Ђz�@`=����n%�T�cZ2۽�X�ޭKU�B$��d7|��!����T;�ba}����B�i�w�t(
=T��K�!j�|bˢ(3��+^�&e��Z�E�۹R�v[�PӀe��R�G��ET�����³�W*ϱ
��H�,g��!`��c���R����s��9Rb-�^����87$&�o��s�����MO����6�}O)]*����?bD�(��
n�R��y��e��Fn7`�?U[N^��"u�8��h�E������2�Q���D�W\�*׆<G��: �����(��3�S_�JP��@ei�Ƶh9��d.h��Ѩ^��2�簆��RH3[��#rD�@��a�vU&)��)Z�9Ć�r^W�ʇ���h�G�t��h�q�|2�����d�M��_��G>ftS�I�(T�L�!�j ���Y��5�7�'��O�hU�AF�:o�3��K���h?S'5/|n)'��ĺet�-�j ��%���	$��Bq-�:Ŕ�boj%�ތ,�u���-i�8Pm7j7LsE�ֱ�;2�s�d*�Sq�Q�Ft���U�y$�_���S	w�L9�!g5�y�7���9����'�Ԥi߶a(��ď3d����65o�"M�>�\)1t7|Ė��O��QR�
��x��H_0��^�=O����Ý�$���~�'�K�C����0M��p���6�xd���ߑr`�Ȩ�3L�9�Il��Q�r)����֘�pk0��A<�t�2n�H0��-�#ː�-s��7�_JO[����5�@����1��?�
��a���:5�E�5&�J:7Ю:���(�!$�:]z4xpF`'$yG���\.T� \(;Ȳp.��K"�j�L��d�xFch��D����y��E&�OS����p�&`S4&�V���3C`]!���Y=����$	����m�A�|���3�'���r,�M�l*B�fy��=���6[����8�����8�u��+1��p�,�V=�c	m��&`d��?�Em�T�2�^8C�5�$���Pv��g�6��tҹJ�]�w��F����5TA���o+�d4�ꁆaCtaM�-�`�5R@���v�Ʒ`��P��˓`�E�Uq���Kgũ�WU��B�	\�A$�B~+3_,�F�l� ��-!��1�V#\Y,��v��X7XG=���?�9d�6o/x�hr��+��{7��Ɇ	�N*Q�=uٟ�H!sF�Sy{�`oJ����5�5���͔��H0��R�'�p�H�iSI�5Y������}Ng�p�p.~��F!�h'��CJ^����\�ˠ��;�|�	��2�ZP]�ڍ�֫ؽ��Pw�B���� ���>0
ԩ��=�~�">�V��O�O�>�Y�5�Y��>�LWl{NY�⬃"��	��Rl[��(�L��]��,��#3�ArJ��=}~�Յj#������kc���+wY�����շ�3�wa�~�#V'����1�8��ܩe�ϣ���>��y�Y�0�������~��,I��!|z��/�E����F��N˜W��}��j�"��ᢝG<N����E����A�鏊���zvSN10@����/��0�nbv�le��9ް~�@�����ĊE��~r|�j�/R�ѐ6��2���,���G4�c�#t�E�S����Di$��Wahځ��󛡓��h�qV������s�2�v!�y���b��fdT��g�y�9����I�pQJ_W������I}F�f�8�����Q��*U]��}=P��ZJp�:b�+���8b{=�{�~�9��Q�r��da���B�,�r/3�CS��Xv�T���A�Hl�.t,�r6G�)$^�F%��f��|�l�S2�I���""͊u+_�!�9n¿֘V�3L���q�|��a^%�HGL����ۊA����O�C]4�Va�A_5��K�瀒C蒠�#��a��S�	���6~�l�TU0.+�{������#c���1�;�j��=g�`�f��x��ngfh:�����A��o��{� N�eۊ���P������iO�z��ҋr*�d����>�o`��o��"�!y�7��9�?L�m�[ �*v�X��q�OΒ�!����l�r=~��p���ZZ�49h@7Ѷ�H�%z~zjdr\���Y�Ck��#:~/�@T�`(<��.k��4�`(��������yK�P��/T��;mOw
%V����p�A�1�[nB��s~�#��*nc`�v٢����I�º'�e��#c(7��E 
�Z����8h}�hV�{,�)�����LP��筰�G���pʙ?w�����"�����:⭒�o#���t`>���U�\XSSK�O�OQW�#p&�_��8��id6Oi��q����y�?��\�ۻcv���gS��B������,ñ�\7����(��3-{Ns��X��nDV0�y�ǒ��4��_4���3|��o�!`,@��A�q��{���C����\������j�/)z��CG~�E֤�@�Q�L������>��Ӧ�<H%�g�{+���nF�I��Ke�Xk�̛+ �=�ٿ���1b��3:|ؙ�L�H�n,ǉ]��:��w��S���2h֥��j��B]��Y\'�{���DP�޳������H㓸H�)$�{s�xZ,�+��=���u=�?I�]��i����;0ro<�5v
x�!�T�X��Y�Φ�<Μ�����Sq�����ZX���()�E��Ջ���	B��{Gʌ|�C[�o�X����5���i v�����jN�O%�6�|�-V���xc4�ab�T��5���{7��
nJ�һ���W-^���	Jr��I(=��y��܍�}��U�6p��!o�]��r<�`m�X<b+�8�kzt�Ĳ0)��ʡc���7��7Ѻ�{�Y��"�h����!����?R���F	�iZ��*������u�x�R�K&馩�)jh�\Fݢn����.��ۛw�+�b�}xW�]��������Q\���oV�2��Ov���<�f
�'c��m��H�2̣Ϝ^SO�zͲ���y2u��W9+Ս>���E��:�b�ܣ���.�~/�z	����}����}ef[�+x��P�qj���Q!�����e���g�X[`�'Mn	���������^�D��c��f)�Z`]����=篼U��"#94A�:��
���+d�o۷���l���q�wF
;/�n��m�>^@�E��H����Խ����&O\v2Y�fQ)Dz�.X���Ui�E����"�@R/е����z��,�k��GR��n�Y4�(�|�D��b�
����}%P�'I����Bh���L�,�r_ Z2`��qO,�!�kw���[}id�*a(��{t�*��K��At��'���~J�F�{"O�F�@/��J�|���6��D�_\�:�^4�xvl�a&�ny�W(��d���oX:'��*JC(�2��Њ^�o�>m���di��Ou:����v� xN)�}f��N��,���4P$.@�dM��?����
Ay�ԑ���֦�d����p�������+��v�j�m^���#�Wc`�Yk��� ���?�	\l��xʂL��0���5��;;\�v�1T�p=V�z�Lj�g�~�zV��u��F$z���)5�B	?�k�'x��w��׺���#rBR�p��++VF^����۶�?!
-V���B��}�-�8YP�׌(\�����ӌK��?�!p8�RP�M��q��4+6�Nh� Nʳi
�S�p��1�R�i��SE��.���nd#,G���q��h���
^��8�LI�� ��ߪ������v�H"?��<V���4�(aǧ�3`��5�8��M�ì],����B:��w����]�z�pҵ�n�'wP�!�w,O�Fh0b;3	��i1T>+%��f���{��*�ā2NޕKqw��Ǘ���+Z�T�y�tE�3�A')���Y��>x�[|t��\5��y�G<:MQ��Q�iIn��x"����j@
@ݗNa����8˚�Ţ�����Pȯk
-�����2[捊|����*3��(KޖUn�����\!�\���]^�:H�����&�!ķN��0�㑬��MĿ �1P����Tِ���?��|	���9~_2)����q���Cy�E�4�m�)���~v�r�]h���i=Ť֖�<W��H���T�,o�Y���AӃ�*���Rb!hq��d�������.~��a3�ǌ��Q��j�����KlX�,T"4� ����jI�U9A�Z��pL'(!�S
�^�3�����m.]#ǌn�/7}��lC9TS��l�����n�N��*�59k $ X����NRl))_r�D�m����P�_h��@�tbyS��bi���,��wō����	
kX[�W]��B#��ԃ���j�y��8��%9���5��Ǒ�;�3T�����<��Ez�c�m�DQ�d��a<�T�������ܯ�l����*��
!ջ��mG����<����E�M��a<ۏ<,+|��W�<k�=�"?$�u�����=P}-���}�<jE��Ô%�W�C�N1��L��X�-_ˠ%B���'[�K�/�~�3c(髪��N箜g����q����_�㜬2D46g�ݴ#�M��<t6j�SЌȑcp�0T�/TaAwxr���ŰD�Y��[hMw�[7�CI����jح��`���m��] V��Y���Ҙ���{u�Mz'�<�H���	C��C�T�!�h�*q�l��:R
����+���m�O��*�*��Y������� 
�ʜ�?�Ӳs�A���pL�'��H�R��-�-��I훥`k0�/ɦ��E87�+&m��(�\Ӝ!$)���߅�#��r��~)W�N�vR�қB����%�ΜJD��<���4)�'é��g��[�r�kwe�J�)+���4��&���*9`-�:0�&��d�����(%�<��E~]"�����pZ��.P��Ԡ�xfGfw�5�~zj���:uK���ɤPs�����U�PM�+.��?�)��N�#Ĭ�� L�m8���T]��)��I�8���5�S`�v k��+���^��穿��uZ�T�l�`^��.#{�����V}�~����UAT
0v,3�F���
G��
����	���ߞ-4���n�ܺj?�⩯�ߩf]�8�a.Dc��E��Xy�ڢ����$���V �n�b�[L�N?�c�`�