��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��� WЇ�<�$.��E=����6�E� _��'$��&9�eibHu�W&�!��ϴ��N�/� '�g�nMJЙ/r�h9����
�3�9�4FnZRV����G�m�>|��}��/k#{ß��}|�SE}�v�RiH. %�I��':�7 yY���MݙU���N@�#1P���[R�w�JP��4��g����zKb��Gd�R�B-�w��f�&�����X���c��H˶����GB���.@Z\�\ h]��=��٢M�ţ�������?),�<�+?򘕦+A4��F�:O�./:��@0��o�~��a�py�k���E7\q�HD��ĳjSY�gOr�i��0NE���29�)J��}�u/�f�}~�*[�o/��n�ƍ�?M/0�P���U�aP5	J�!��D��;F��u�-�]~#��Yαq?�	�55�7q�F�pO�C���~SA`��WuĹg��;��	`|�;q��#�\������jYژ"ZF��%�Ripw�9#���$���%�G�IWd_�)C>-�q�����������}�
�@�꘼���o�L��,�k��d��6����K8�F�'�B�6������2�Y�Av�r�w!\��zT�������K��]r�>H��)07x�M_�x�;$xy)�e����t���SUD����t�EL������l �"�8���Մ���C���|#�W��4"
������$׎�ou�D�h��&SZr;?�QE�]ZD��z!�0n݋n^�F��Sc#q��zG4�T9��E��-QIƙe�7&0Mm�tښ�2�
9,[������y`�T8K���T��K9 Ms4j0Éd��*(�1;.<���n��9c����� ��kS��n��������ʑ� 㣶��+qp���V�q�9�j��ˤ��ؙ3�`������Oo��Z��qVu��"���Q"�]H+�-��f��nd�%e��*�����>���p����^"�Qp9r50l�b�&(�RV嶍����f������SE�{�|%7�W?1��4¦+�X���	d�q�8Hs���>b:m�+z�yzvC��*�RAs05�JF�gf
bC�x�ś̒����"�K�OQ�"�M���-��dE�	�C�s�������e�{�#�����|.s�O￰��csT�R�b^�w��M1�o>pw�w,�@�r"�#��^D��U�L�~ݯ@���ۮ@����(�<��� �E����{.�r)��$�vI]m.���*�x;�X+O�Or"�f�F�͙��ӑ"Z-tt���5�v��n�<����"�~�����#35��rbI2�;�ph���E�~︝1��r���5�q�
�I��]Y�C���y���T��/�4���೉�̌��e�R�� ~�*����Uߧ�(,�J���^���;O�&�<�)��u��X��P[�H)�vh�W��+k�0'��V�DT��Œh��A&Ií1�X!!VF���^�<�E󦣗ȧk��mi��HmD�۝و�_5,��#�:�ū�H����.���g�vS�♫}M��t���G��nc@ZHk��,m(H������"��8���^�3rB��PeCj�*�r�����^����r~���]��V����\��'��{C�:V�쮙'c*jj��)�!��N�0��{��t�y�ےX+O�$�п�犯>h<���2��!������P�������+��v��^
�ƦꐞX\u�Y(�OxK�X�7�¦,�h�LB[~b	X�f��q6������Y�$.��׳�,��}�;4q��7�r76$֗je;��>�ً�t^F��/%&����(��7չ"g,�m��iY��_���[�i��/�k�Z��0�L>���1�uq\�`�^a�Zwܓry��&��_F�]6^콗ܗ�R�`�7�'�<��pW��Tl!Ԑ@��� ��Ae�$���SsOge?&*�@�Ω)�p	��q������"f�ۓv�ƶ� ���T��G�-�56SH�4��D)�K�tmN�6]��� �-��隊�_���_u�*G��$4��דXV���}N��]S��ŷYNu��.�!]X���A�
��Xlkq�����e����쳯F��0�r��h��:L���[�\k3�'+����*�I/<����Խݞ��{���g��h���9�-2� �[4Q�Q�v#Wr���5�ֽ ə=������岔�_���{!WX=�{��ԙH�I�vZ�D/p�1I�K����P��OLX]#�vC�:T�/7�T��5�l�Go"^�|�zLՋYQ��`��kłַ:H�>C`?��H���.m҈qMS���@?N��p� [�c���1s�(�E�İc��zZ436.�49�"(��o��c�"(�/���`Rv߆\�mu�@u�e�uo��&���o.���K�U�䧳�%�H�r��p_���g�и�(	��Ć��ƫ��t��ro��z���u�k��2۳#�٫�(�.ft5��� 4Y��1��P0��!p^�k��LaI�A;��:_��o�KC�T)��Z0@��{$J���l2�F4&Y�5�9�}��s۞j��p$�KCb��vӲr�ﮩ��/����v��W�Ĉad���>�w��*�aU!tÛiO�sJ���(��p~���q�G8��9i��[�U.v���E���֔[\��{u���jS� �#�0�B�-ɀ�Q�A3;��$B@8V�U�.��6
�Q8���$�l��6�x}'F\�q���5�_�%���Fu��B�C�cB���r[7ӷAs�_�0�3�]��(��"ڭ�f�4 Tn�Y���ihx�ڿ�'�-�,&��>���\'c��%+�5���۵;�E�B�I�(���Q��dE����I�!�e��U�L-�z+�����란��1��p�f��Ϻ��"�
���y.|��r�4|qߚ�t�����_�?���N�Ƒ#^w➣��B��5��={+\Jj�L�F9Kb@����zp�(jr�	D�������B}�Tdk.#��mq`Da��3Y�N��Q��V�Tc�wI�����\^?��7��5I|X��*RR���qAM�/<N�i�7�J �I]�g3��賂�c��H=�kJ�Pd����@�*��@�ӭ5!���ok"��u��_"c�����瑘���αy��y�����xw�u�^��ʡ��}���5EE_|h!t�x�ĕ���
���f�z�  F��p­�q�j�Ta6��L��8nZ�Z@5���I� m���^6V\�s���\�e��H���]L�Wﱴ��;z����Fk�쟤�C�$��չn,W6}��r�\����CR
DK�!=����Gp\����V9Y��iZ[-�Ն�D���j0h��D�Q�>5�muJB��{[�]�K8� u��Y�o���dq"K)�}��W�s�2q<7�����OXٞ��&m�D�5$�*ߊH���r?����}6ـ���u�Z��|9Ɣ4�����_2����.ٌF� 0�� �����@�SS	]��1MX��ަ&�O!)|�v��9!G �)�e0��d7�{
u�6�e
A�"JJ9�|��`s+L�'�<��f���[0����&�>H�ӡ�{EX�w�ٿ0[�K=/�ܑ��~��S|^��Y�٧��9�E��t�Z�NΫ��s�_o�)F2��Vxt�}��jrw����G�ɣ�b�m���`�v76kr_YI�;	��Ig@�H4��hI�t3�Z]�@�O\%�h��qLG�-��yh8,j��u<�:2�s��╃~Uw�] @��?b��(�f�7����@�Y�B��&��\I���Y۵��2Z��6	k�8a5��L��C�z�$&$4`<Yhɀ�d"8�X�����Ã�tO��s� �X��l��"|^Z{K�faP�|�_E�񳿞�ޕ����K�bn��Vw*8JE���?�k#]A)T�7\|Oz?�މG�Bf44�l+?����41�)0��:1E���J(0�8�{��wmp#��T~t�g6�'�������*ct�"B�)X��J���VU7��=��R�}��c�.����_�:,�H� #���*B�'�����^��O�Z�iu��Z��w��V4~��4yRt���jv͛����.��vJ�v&�T��	���f�ǣR����F5o�;��C��<�\l�Bf�$�����Nbn��A��� +W�&��%���8�k[F �o�(�)�uA�l�#���h�v!kE�C��U7�w���������a�� ��0AM�JXt�_�Q�<&ZOt�9�.j7�N��r��ٚ,�&O���.�{��G�|��������Z�QJ�]��Į�!Y�O���?�
չ�	�ykՕTO���$E���������w�e��%��|��o�aeT�G���'Z7�--ɦ�C����" q�����v���������3\��i���M���Z��p��(m[�0��u،�G���At0��Y���n���j�"fc����BCJ�!�x N�
*蕯�V�8ڍ�g	���Q&MUd�����l)�t� }��oE���E��o���g(~h����Xy�GtN��EC����"�n=#��� M���|j� �;io�Y���`���"%ّ���k������V)i��^��(wB�V9���L�T��+B���1?!��;�']�
�:����l©g#��me!�qh6������<�'�2��[>�p&�a`{3��7�HiGX�]LN�L�]��3���E���c7�WV�	>��*'�:�,�����B��%7���'~E�j��ߍ"'c�BG�������n��4�� ��qx���PG#�t5�|g_2��O��?�h���6Z@�]`��Z�Yi9u����\T�?"�H��|�V����^`NUl�WA�Q.޶�;�:4����Ma��٤޳�1?� b��Bt`�7}��aIf�)�r���{
�9c��Q����QlcC<o���>T��jB��4�ݫ��q�v.s_5��&��NU-[��5M���h��I/�S� �m�K�Q���e$1�B�d*�g7 }�?_'�k�Ӻ���{���2�(⤒��=#x�%���n8z�U2��;1?�ZA�Y��e�C|�g�T�2zF\��5fc�5.������9��: ��*�U)̰��KO�G!���^Ww��U���+�g{%�Ї��wb���#���
+Ǯ+�<�6�x��:x�&_ǲ�gi#�����Hk��n����.]S�IZ�!��Sm��$@o�I��ٹR��e���c��IE���Z	ΰC //�)���a�j	�Q���������	�D�A֙����BwJ��G�q'rS6��&�E��{_����q�ͨ��5�E��Z5�oܞnXT����0�oYD�����}lS?�0n@��KQ�BgnӤF
Ɛv"�r�(J=��e��h�y5�;]w���+SH�b@�B$��/��ZSD�Ȁ�P�TG��]g����)���bQ�`"�N�����J�4�G]������l�j;��A2B����M=Ѭ���y�I̝h��֡��Uȁy��@����x
! ���/�6�n�E{D¯�_^�¹�(Ok+�W9���/ȓ��Z�r����f��o�S��l������3�-�_Jl��������.�Y0��$��Τ�2Ԩ�	�wb1��?C΃�n����.�2�AUm_��A�@�OJ��!w�e'��%��s�5���o����k|���rd�9X
�+&���帖��o갋^G#��"�����:�	k�ؙ�)�HہA���l�=�P2� i����P��qw�D��BB�%S��v���x��u�.�i����guhZ�ȼ3=p�`Z�����)����ko� �H
r�Ldΐ����=���C"��ā�2��?~y�3��|wG�*�Y>Ez/� �/ލj�ɞ����O���,��V�t�w&��ȑJ�xkbQ���8����(,�s�X0�!I�6�����01)��*o� vD��Z}��A�ݭ���y�%ގ����QֈW�NT�PO�-��r��q�_��5(�s$}��/�I�U��V�К����t��>SnIH��e���i�>F��1���2�?�JӬ6�� �_�A�S.�Jo�hJp3�����QG͖w�N(����ٜ�#
 {_*p�c��#7�F�,�-�Q^/�3q�#�Ca�S�ъo @����$Ӡo\Č[aW���@�D����+rR���5���F0U�W�{�7�I��nه�>ͣ��!��;7�gf�.MNҋ˲f䕹Qג�{�g��é5 &��l��YK���2���:��d�p���]�U�ft(F�؃|cd����^Fe�����6b�Z�T����[�ch'���RVd���
�a
A>�Ą��������/L7Ǻ�ك��9 A?$xzOk8m�������|��"Uoh.�!��/�#&���]f�c�[��""�W�P*ȗFF�
UL����H.��]I�>k��T�Q�Z�����(�Һ"6����qdZ�^���tB�ֱd)���v�BW��Tq��}j�X�)P���FI����z����hK���������MU�%fؿlX9��;ȁC�.�ӆ�~�<�4m�Ϸ2��u�������-9+���I,����%	��d�5��:,ʋ�������!��I�t�so�u���G��YGb�摔1[V�cֵ}���)�����z��i�M��Չ�3K�~��#↫z����j59�洊}�b<�=O�Z�[U3X�ё�RG��6��D��T$��IX�>���0�ߒ��|붶�Z֧9���%x���7,���9��=��WKZA x!��{6�f���]�VؒEY��&*�WaB���Q��d��h̢ ��I)�R���p\��Jpye=���8��v�\.ב+�@)�������#��� K�v(_�A��3�H"�5��]�o~^>��,bHԌ�B@+R	k�v�k�e�օ`J�C�*u'�!e��-?Dfx�dڱ!���Y���Ĺ����*a�L��A��"%��`�)��g`a�Vŋ��.�Ac�<[���m�C���N�\੪�_7�;���bZ
��+��%���9[� I��QL�#&B�S��]RF��R�}�ߵ|�����q-�᥽i脈oh���,�/`��VP@h��Y8AG�RCv�����wj�Ɠ�AX��*�������	�� �&1����ȋ���/g��@39�m���C��y�&�������!�"��iG��mz��a�,DԤ�k�����	C,#��Oj	~E�0��N4tyT��6<�O3�[@/���z~}Z��`_K��Y:s=���͐�p/��Q�0k&�J�޺+;���"�hMrtl���T%�����.���B��5f<�2>���{qUN�~�C�;U�Ӭx`jf?X����D�zh����*`$�h��*
�G���=�f`��_�1�E�MXN�b��ޡzfm[��l[)7�G�M����J;]JE��2����͙L��j��-����q�?���`=D(8Mf�G�>a�NS�>��� ����hH�,����Am�_�	N>2�B�q;_�U�R�`0�C��v8n�j7 ��]C��*����m�V�1�� Ii`��wGN��7�A`�	I�M0��.����6��>@�t�M6Jң�@�~�K���'�$��!�6��p��6*NщA�N�?]q]<G�ȆkZ�3�޽�g���)��/����yϛ��f �kL����&�čY�)�
+JZ��0v�l��E����ᇇ�$d��ZIEPe�O�J� 7��bm��6zqg!
`T�I?u�H\��0{����j�Y�L0QA[Bْ���_�KD��^@�H�]�}�ʒ������/6R�[G6vK���f�6?�>A�1o`�V�jc��5L�5_ml/<�jfK��_�_Y�8�R�X�c}�#���$n�%�m;��:B𾄩��Pu��Kh�
����u���7XQ9°m������\���=S� C؍�%��ɑiiyj=ԋj�=}�ޝ����N������#f2|2���&�s=����*(<_}z8�	�yt��z�|0M�����h�T�|e���q!(7����e�l�r�U���k���}"�R�s��D��/�c���.]6�p{��CO�,�l�p��xi�x�����z�TC�+v�H�q���A]�M������\�.�
�k��K6o�����Hϒ@�y#n�<�n�ii-�_c9;��������AM�;���3% �O<}j�>3`1q�=�N�ޢ��q��g"k!��Zj+�N�s'�f��p�eW�]*��zأ�[2��"K?݊P<"��I�r�/2�M�`m���Ji��^�Q�q�!�v9��PҎw�\ �$'AR�Wh!;My�r�4����L�Cd "��@hg�G�Ոz��L��n�F�7~+���K^F�V��J)�a��X�k����s� ^P���l-��ₛ%V?�~�Q������r����Ci����¯,/�?%�^#2o8#v����	����09���Y�a1�E�H)�z�o��[@�S�@I�U�+�����s��:�d���=_��W�C��\�$���A��{�o��%W;��/�?hh��ҋ� ���ޅ�r���(�|�Ҭ9�Ŷ����w>�¦�^׮:��5�Q
g��J����;, ��+��ـ�i�w�G�c���A�nvD��B}P&��w�Zz]��$ɚ�>O#o6x��`9��Ÿ���T����3$n+��n�yl�%X5�C�v2g�/��sLJM��H��b?����w�wp�!�� �`�y���j$�0��#�>IF�|ʁ�8�!{��������n�q a�G wI��!��{Zb�<	�7*�`2({;#��)�F��-���K���w3���	B����9�C����Q$?�U�\�����K����%^�D�:�RZ�xe�	�TƮ^&�L2��#Q�P ��Ru� ��YʭN�0�"����32z�j4���-^�K��@��&�m+(GAp��l��D�����K��P0�ְ!5�N[�`�İ����vOrZZÛE4�9��^�a�&�B*�Ͽ6�*��˱=��^�L�͕�
��$�s�X@Δ<��u&V;���N�۷�
6�z{!���f��,)����÷����/�B��6���ɯ�kQ���T�
3�/L�v��0)��6A`�$��%��`M0ag� 
�N�	��Oӹ��f�Z4OD~Yww��x��=�xe��U6�Y�5��W��[�n��m�KH�EG�&f���]�%B��*���FKXa��߾���	MU�9s������5�~�VV�m�!edOOȐy}A�+����c�l���9�S��^u�h�9�2\��8�6s�#�����1e��{�{A�lo�pP.�)��P�7$YK��[�5���\d+	�z����aUu��U�)*U�����fw]����^�$��N�5�+x�N�S����ݜ��w�Y&��e����ٺ��2��K�hM�q��a��*ӓ憪�AbY�D�2$f��A^ks�Ag�1��g-���.�ϧ�8_[�qJ``W�2=�!���I\��/^�.�}���,�
��:Ό�C��S�������D)hq �j��!}i�^(]7��Ĝ�j{������5�D5�����5�#Eh�}��	�H`�v��.�lQa��t@ �_��3�>���84¦X��,+Em��=��
b\u�(���)�(f�:{][�#W�s䆟 E��4�g0*D��J^7��I�w�@e�>ݨ�����L�?<�'z
��U1��8�H�1)O��(��m�����\l��J��6U�+����,��D� �A4�"$ތ���ݼW����M_ؕ��s0��-o���Ji �pF���B8�iW[%��Ŝ�IނT�S����3��������h���0~P���!�$�(�s�c��?{a��q�	��w�@4p���0����~G�8_9���e��2T�@a��#�jK#� �����[l�ߢ�:�������o�݂S"G[�<N/���Q
	TzJL�\K����#)���֝5Ʒ�'(��j�H�@W��z��� 
��n�����tJ N48<ԊgT���v�=� �51`b6�������i��[��x��^p�5�B�J�l
�8�Py�<��@.���#	J5I)������y�Lӵgz]?�Έ
���W|��[��:C����{�P�m�Bqߙ@8��H= ��&ԗ�k�7GA=MC���=u�g޵���(j�ۓ�b�Ԗ�ҡ��9$����3;��e������`�Fn+M���N��Y�$o��#�I(m��������3�T�����7r*�܅�f�C{��c�7��e�a��%�Q�)�	�*��"R&X�2e��z�6��UR�2��H�&�˺���>� ��E^��H�Y�x�7
 p;�=�c�X!v`w§<�~���'z�Y�,�xf�̃ >��S��gY��,F(*{nK����_���+�/��ɦ��lJ3���	�;P�s�fra�C�d�o)j��u����3��8�<]	���)��:�~J���P�����.���c�+Ǌ�Q�&��W�����^�fy{<��er���H>�}�&�޳��):`���S�Gޠ�(]�t<.�%��5����0�=� O��6��|�;��B�R�S��P"q�ʾ���R%Dꫤ��:�;B��m� DVY�8y	��4}%�M�:d<�%��I��

zqpv�;i���H���蚚%��v���9B���Zs}�)�a<�K��QG�]��LiyY^(('��*p@2E��nz���Kd^&�n�X��S{��2�G�]�3פO��������f݋�^�DⲤ���v��n-������-ї���W{%3q�|MSأy�'���嶁X4"�8h�[J��{�J%�P+�1.C�Տ�	�GyD�/	�rI��{pro��4�3YT f���x���U�Ǜ���]^̚��Dt�bI��ԺE��ol�дc1�I����D�H0�I���Ol�a��e��HcA�ED�Llpp���T��I��Mv�F��tP2�9)'tL��H�������F�p:��kR�����.�&��b�Wb�Vi@j�U�Z.��,ٹ�܅ـQY����>/�ġ��ܱ�Z�T�R��.$#eυ��"�mr�A���:�b5��W���b�pn+m�-�}�❘�� �t$�Hl=A��H���1|�I%��b�^�O�s�D����-q]��)�b������W���ߙ$9iKm[�tV����,�xF����HZ����U�d&�>�O�U�Uo�������Z+�M�A�i�����qїݣh$ր��p���������*���8�+�ɭ�s�k�f��&���H����qO׭���o�/B|a'�Ԋ5���L��K��SOX@�d����"Z�6KX��7V��J�� ���F1��)�N$ ��wl��r��Gͨ�����,��y��I�"��@{v
u��ޝ��^>�����H��m����ǜ�[FL�Z�ߨ��c�ʫ'UC��CV,��u�*�.Ai$P�]�����O���$��-�f�UNc����%Qt��T�VG���C1�fuN%���Gq�r+"-����6�lq�!�F�l��;�
sc��[ϝ�N�>�gg���f�I0��
�
�����Y��G�v�;�H�8�E	o��'愒�p��H,h�g�=�=]�ցZi>�k'#Jˈ�D��Ʈ5��f������xA�%��mf���m<@�|h�{�-��f�\U
]���=�"�W�Be�7_��B�{İ���F!��
���02!$���<{ও39D��$�=1ӻ� f�7W��ZwI#��O>��;�>^I���
�Px[Î���Ek����z�x��,a�îST`���C~�$�\/�"F�Q�+�W2fxR�ZJ�#�'��l-v��r2̧@A�U�,q��\��&�Ց��U�pYv�T,�YP�3�_>�Þ���Xڐtp�L
=��K.GAɋ�Kk�
i�y#���#x�F�SJ�����6|K��N�GXkd9c]G}O���Q���TK�1��o�U$����>�u�%��]�%nQ+يF�|O�| ���\W����GQ����rc����3�����b��T{7 ����ԬV/X�d̆�l+5���m�d�N����Mp��F
�Q�,�P3�|�;�axPZ��k�2������;��N/�X��b6�r���T��JVe�m�H�3��R ��G@�kx�����;3Q�O�l#,�"݌k�\F�&����5"�Tm*�(�����z]�3��~���:���Wۘ�b��$m����)g/�G��4�c8�͗��t5�/���o�b4�X�i��Ki�C+g��r�_�_��\+�/q�k[��ҝ���H9��dH��&��b�Ņ�JB}�p2dP�:���K|�a�,7ӁR#���	
�jݨ��a9m��8��1��3-�\>l�g�& �h���E9�(;�47��d�_[Wy����&2��_�����k5q�X�L��-�ml��VA���c(~�#rzb���J��UlS^����ւ����q��R���b�O1_ۄX����0NG[1��G��?��Y#�4/���y�f��q	K:��i4X��?g7��[���d,yv������k��#WL��:P�z@"#�H�0\���Q�`�����Y���g1%Oj��\�R/�;�oG��_������i7{a�%�E^��g��+2�q���{���>�g�A�:�	A�*0OwJĸ)�1�<��ʸ�Q1f��5��H��b��sB�~�/#ٯkMaSg�yn~b�	��(�L%��4z��LM����`�qt^S_,�������j�K+���j�܏� �Fù4*�S\5��UҪ�B�z.[3,xb2�Ʒ�;�Xc�5������g��[����H�!�Z)
�I�sg�n29�ց<bTW��YѺ�ا2�t6ފ
'A��61��G[��ϙ�Lf����E�3��*#���,q[�@�b����=z#�u�����~S�&=f�`_�5{��O�tAD��D�.T��I�@�1��{���J|���	�!+��>�P/N(&Y�)��."ߙ���K�/&�bk�%�S�E��D�fۿ�qa�4u��2-��⾡�䋁�{�����uJ�n�åCw;x�#�X���ET���:J�'n�a��hPA�N<���&i�!|lg<H'��xO���R��N:�R�kI{��-<�G7�J�=%k1�P� ���l��d��5�����d�����,����<�؊�o�̩j�W��xC천�N}8��y7"�N�A��e����(#2�n�d(,�j�~�HĶ���z�&�n騑����2.!��qV��겷7�k�����K�B OefR6t�A3H�/q���E�^� �	,"������}���7d/[�L\��|�wI�4�����q������G@��(�@�ʶ�&!4���g,y�����;v��+������ziӐfq�6�����/W�XK�7��5��8����)@SD:��XǺN,E�3���+7!�Â�â-�i�q��������}�Y����a��c���p3m.��ӭY\�;���#"g��AN����#|��-�Oc"�˧�<��QĻB�R��#��{g��s��H�F�"N� ���^�/d���`Q�,y��(�ݐ�-�-�M������O^-��:7���\�8�i�!��`�n^,ݦ���
J�-�/�$D{L�G�N
��z�
[Z��"u��e����n�Q�f�VԎ�W��/�M$�I���mj����L'ut�pR��>�Ox�Ψ� �"��!�F�@��'d-�ޱ5^����B��6�-���H�)�5�Wt��Լ��H���T�c�c��!쀂w���&_���㯮)��t$qS�rp��W�� �r�c���E/gA**���U�x!gN�/�K��jk9�)d'�ʕ2���u+n잺��٣3N�>�Hp�ŋuټ��Iٙu׭b�F��a�v 듎w�G艤���W�<T�a�󡡪:�2��!�;�
]{�����i�$'�v�xQ����{�b��� �+�[�ȳ�;���XeI�]����8�zg�Y��IT�h�=r�v����0V�J�%�:��i46�mQ{�4�i����`n���C 	�U$���M(A�ש�"����?2�g1���[ɥ%��we�[F/Fݱ�)X�-N��Ǘ|��1�V=�nvk�4�t��0C�j�P;p��s*�R���^Q|��ԡ�\��-���xo��sP�@��D��M��i ���<�p�]a첹n�*`����=���K&F���p���¦��|R��Q9���uf
ʚ ˉ[�iQ�ɋ��B�嘕�mTG+�R�������t�U�S|>J��H�צ��f�I�"����1*����]��6i�RPMmq��Yi��D&�����pwY L�AO�a��Ҧ�|wW�#�oA�-�h}��=X����t��1j�-g�no��s��<b�|������F����!�ji�R.9�|[+�bn �?��P�ا��J��@AA��	�AAҺ��^
D_�ޅ3�[�Ay"���U܉�uf�p�q�7�Qf��@|�$J�E��TC��f�I�Vb��b�M:^�!��@����[��{*V���BX@�;�zc�<3w����
����*|�gtIi�_��2���~�Ȓq�𿒃FBCëRf�̧�/(�{�I�}b��7�<�T�q!*�YQPش3��K5T���Pj @;��{p�'������/�KDw�L�0��ԙ�Ȩ��O�Nh:\���g�|b����Z�@���LHrYo�y����.t�l4q�� ����7b��@Tv�]���E��_=���<���;
��H�N�e�D�_Y�V��v��tޅP��̮��m�N�Jx�I�~^�#�]ǋBx�ݠ��sY��OS�q���/��&��dh5�Ӄ��P��;O��n����� Z��p?�0�i���2u��[�9�|����i"��[���{�Z�`$i��0@Ǔ֒U�\��ZM�b���2�z��o�g���o�ؿōG�n}s��hx�� c k-!՜8��-jpD��)?�?juROa�`�!�'7����~�jo�_%�g�V��3x&h�E�h�\�O����m���F�ע��/?�4M�"� ��5-+�@�b�f_��P^Ď,}6��g��c��%H�:m��X��ʴ��?̆<cC��GC��zx�u��DȄ�Ki<�` �2��̱�Z�Ge�a���v�tC(r��H!t'A.+��^�����v����a`m�	ć��B�ulyXZ�{@��^�����$N�A����kA�z�1�L��(��FŁ,�K�o�Ȅ�)p��DM��t����ωݭ�k�Ѱ����Uic��'�n����Cr���Rv�Hϱ{���� ���J�n��cx�yWM3��ZVfR�(��E	�^5gå�5�ГG���3'��j��`%$��pt��� ��Ģ4k���J{1�A3��v')3*;0Dvȧ���P-���83��l��^8A<A�{$w��(G��������kg�W0�DՉ{k�3��Lm�À����/���d�nF�����^�.�B(|��'���7����?�GS�S+4��sMY����\R�.��J���p6�bjZu��������N�xἠ�(��@L�j8��R!>�����D�l�AxO��Nq�EW�2p�&:�h��@uz&"XBn��ՠ��U��97)2T��2�=t�o��Ô���e_���,�@nA�D����Y;mf3�Ż$K���4�9����dZ�����9h#Ȏ)��f�L���fy�3:���Zb]��H�`:���H�%�kqkL�2F$oV&���M�\V@H�3}�>���J����*����$=�W��!��Ĉ��r�ө�z�y�ּ<9j|n�l k-�C�ӊ����$�IDH{�	�*��*��c�����d#(�a$�_�ĨR$x�ر�G��h\9����{/�_+�G�}x��)/-��Kg�=��ѿ%�e9e|��0 `L�2G!Ni��g���gH�գ��*�ԘV��$i��A�4+��_��-T�?V_�=1�����,���Jo�I��D���C�ͭ)����^�Z(�9�2���ݘk�l��B�������-@����m��4�e�M�(Z��#�z'E���h�솽A73��8�f�&�8�)�I������#|�� Q���ih��R8&6r���FdxM!��7d�n!����8��g��3ΐ�Q��-N��%ҏ �V�H$��᝕.��<�!
�Ʋ�,�h������}���gfm�;p���m��vK�?��Ŭ�[@>�␽fET�2b��T�N~���u�܃DY�]�p�{IN�)����?ү����/�J����cZ���)#��{��Hպ9���uS�>Oj�{�z��L�{��.�DK?#���?��m����r|�5�C�:`_ǃ9�D:U�|#&�*GruVE��R��"�9BZE
��c�S�
L�������G�Q�L��L_�L��s==a��8� oũ�5��o�t~�����$Y�:${b�[�x��,,	�^�]�&*LXgG"
��V�`>�X�O_�C{���s(L���qJ��u�ˎ8�#k��+'��b W*YTr=צv�N�T�E��&g>�Z��t)b����ӆ���/�:������;B�,
I,�I8a�}8�
x�y�v!�!+�M���S��qeiXS��i���%�(W�$��/n�{"pHt�fRr�І�ī����^�9 <�^n�� Yv�(���̎V���X�N	'��uo&��fk�퐗��x����'�Ǭ�̿.�Q-�0e�A��һa�����P�	u�) | Nv�C_��4����J���J8��{�An��U��Ԏ�][;�d���a|�jy�d��g))5��s�c�#	�sQ-����$3���%HvN�e)[���nPG�Z�- �Ǖ�:���Fr/�O{<,ּ�6��v֬����*�����QV��[R�tr�TyxNB{R��\ģx&N�l��u��=Gm"�"��2Oss�b����`0S���6諨[�c؂������)���[~�s�6�vk��0%���\��Μ;������k���͈��ha�q�9ׯ�T���t-�:�Da�!��Euv���H��֙t:8�(w������䓱AV�����G���5�]��:CI�@Q��>�a��Qfc$�7�����Y{���ي3�3��;����m3�F4M�񤝨�k��ᑇR� 8A�0�<p�[�q��Y����bnl��  ;�=@�V-��WFˤ��>��%� �%�OU_���#ׂ�!�����I)$�G���8���at���/����j0�C�xn��?�J�ر� �
�/���u��Z�_�>�5cѿuCM�?$L�,��}nH���R&BJ-���1�ʋAcȽQ�$�����|>��@�)N�R7��&�40ߥG{�P�Mit��-�8}h��Ei�.J�'� .�Wk�F�o�Z*�g�- u}�t�e`h�tI�q���{Y t�W��w�G�a�˷ߝ�Z��7�zb2qrH"��I�e]EQ��G��N3Sp����o�N�oY���M�5�?y2���ŭ���ٸ�E���B�$LOD��x�U����$����_7��M/>��S��xH����x균���'���[�����j3�|��/����+mEs��d�Z 3jy�2�f��2-^dj�	@�nJw��$u��?��X얆�#��U|io�2�uw+��屒����.bO���Ĉn���?��J�+'X,���W���H�v�&xQ�>U�L��I���E�f��0op��	�� �F�7�_
(K����J�ȹX<����LeԨ��v*U�M�v���d;��a2�pT��	j���L��~��i%uz'����PTh�����|���X�{4�U�t�-Ð-�֬���Q