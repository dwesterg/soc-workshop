��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�s��W�;��Hj�������R���9P�޼�ϝ�$q1_��kVu}��b�b�B�b^��%%�%�/��d@	�O��+J�/��f�Y?RO��!
��8H�Ѣ�m+O��4�����5#��̏�����,�i�d��ڶ�@�.}�WJD��.��D�??����WD[.�2�1�QCy������ݵ��8�s<:��%���т.V��Q�8�����7zJg��3<5_�?���@#x`�-�9�!m�����7�fc��E�9���=��.�!4��P>��
���: HVc��Gf����4�D��@gВ:�Q�/~� ϛ$k$R�NIH����)(셻kHX�?i^C��ߴ"�<]��2C�zP�w��9~^7�lf�(al��G+�+�Y�[�jT#Eo��B��I�9s�n8�Qq^�D33�������V�/j���u�(��۠5�Y��A�$��_W4�潕��^(^T<c�lO��K���^$R�X�f���別�vҝ��iP��|���J������*^V�o�Z^N=�Q�I��,b[u���L]?0��o��=!��RE^er��t�� �4JX
pK����s��+�A���j�B�6@�0��������{�y{6VAv��z�xF������ߍ�׍O�ݱ���4��趀�����Վ�S;B|7$~A�cɃ�'�ee���j�ƙB�Og��~�S!�`�Xj�-�4W&��Q��6N�Q��6�OF�^�4�2Q�|�Q�L��g����ތlxL��{G�t8�!�BNM�M��������[�3��R��W�@^��3k�Z氍�m��TU01������+������p��?�]1�O���|sE�~����GV�u�2����V�Pt7q�j-E�w��|���L����]i��ӟX�-�[�Z_�'�:X��;Aؓ|�Mi����Tׄh���Y��g��������P��1�K�gk�*X#7��!uq�}��;�H6Q`�{'�f@H���ׅ-t���:h��^`D���~�D�G�J������Eޏf:�?���TÐ'���D���q��n �a�0�,6ߏ�ά�6���s2���7��y�l}i���*�z!�S�8[�w�������\ASdkl]���J=�`��#��d���f7ʄ�������^J��?�("�[������ !�z,����rr�m[�B��NQs|��(���K�6� Ǯѩ�p�K�<W �ĞčM�2�''��q)�Z��(Xjl>��\������H�" 	]�7���??��ĻC�r�p�%�pv?Z(!����'b�2���P<ZK^�U������u� ���^_*6����5��@*ok��.����W������l#Ր���5�kV5�A@;0��ۅ]݋�S����ą{#���x����:���&H��
N�<c���m�{[��^�e��$ޜ�t�D�K	*Ⱦ'��Y;�K]�x��yV�v�K��Z���0�h1,�_�p��Pw���Z����1T\���	�oCW�ǣ�}��r�A;��#BD;
�|��\�5�(H&�%v��݁sGg��%���e��o�f4B��B?�4����"�3�\6�5��d���Í&HH�w���. 򳁡�Q 6��^�c�Dח~�L��d����Z�V$ڌ�k���N]@BTU7�*�Tv�ߗ���r�?��=n8Jv���|�%�S�̚3+�?��0� ~��si)D�\ݶ�	޲R==�(Y6�Y>_��␍��Y�f��=my�M_��������<�A�6�M���.����nS����#�.���C3�|�a=�ݢ����&9:��5������z�4��y��2�1����7��)��c����ߗ�@��c��٩ ��= �Τ�[)9����L�xo��N���tA�-m�l_{�p��-.5(lDf6RBù��1oU����ao|w�L�Nʻ����=�Y�6s��QS�^C��Q;�oC�Nj���׭��E!�s�4CM�@�4�S�����c�8��ãM���(9}�_)(�F^p���<���gN�b��\���ge�)�]�.�jd�\l����$��L������U���E�8��6�Q�c8�O�J�95�x<5=6�{=����j@"d/�ʚ�^���Wr�Nx�ba=�m#�Z>T��֬d
x�]��A�$����T�L{���:�GP����}�tR��nbkG�И��ҟW��#��>Aغw~,ARͭs�=	�p�oH��{�\�^q �H+v�ׄ5;%Ie��î'Y4�X�O"�bY�y3�Ł@pK�/=5أ�[,4>oD������ի��CTH�S.Y?(�j�1�;�U��jC� X��F��TIՍ3�J��
��Mc���+"����X�7v��<m�>�S:w�WMx�.e�ԋK�t��`X۾h�<C�G���qO8#+k�Z�@ů��O�lj��cj��.�M�R(��0�ʛ�Z~ICJ�o�������=%p���&�]��ؔ+Ċ��ꄰ�|]��~_[�����X��#�Z����+_&T�)�͙v[���q̼���ޜh��NK��ʩb;z��> mJ�4��6ɀ�R���4�9��܌ن|���%Y5���o^��؋��U_�b!<�Q�
f�=�D1�&�����^�7�m��Fp+��X^�[�2��h_�-�U_�r<z �.�O $��������x�S`���E��1���J����ֽץOrW����8�c�^�a'S;{s�o-�2����
y�21�2��'|ۍ\��)�3i'�>�����^������d�H벲-��~�s_���0w9.�]3�L]�Y�f���Mtbi�>����h�������.[�v�V���Flչ�tpyF8���x��K�+hm�]цo�u�GkV����#�������U�V5:0��[y��1��z�$�gԑzm���b�?�+�$��A���4�"���ANIQ|��8�~�p7@I��v�#��he5���T���X����;\
��V���?h�#�[6M;��c����.�$�.�.4544���[?`P�����˕P���eσ9C B�qF�(0(���������o<���Ko��C��}��Գ1k����uf�VN_�ne9�VB	��oZ(0�Wz�(�v�3���G�s��2ux�1�St>6Z����"!30��U$�&�5�������������R���-�C���jz��G6���S����� =|`�kL�������n쵺"�X���^f��i�6��qQ�>�0�pY�o�fZ�����̯1P	'�?�u��h�WQ�m/n%�Ӱ"��V�h�׉W��,�ɗT��:�����5���2ח�����Qد��_s��ZqOC���+EZ ��{R"�cG�����)�ߩ:�V�UC�W/�'�,�L�hM>`x2?�؈Q���� ����<Ll� �k��?�N{}fqW*哋f�9z�|(�E���y�4���`%�����Sg6�~ �%����C�ʅ�1������[;K�R������r�2��X��f|C��I:vx�����挴��J�Y!�Y
���G��4����x�����^ֻ��4:�����A(q_�,1$R�b�O�����kYt�+���C:����+���([+z͈2/�E\������;&�QPu�ɜf���1�$m���]2�'��{�և��9���!��4y[�C� �	'�0%��Ɲ(�!�n��2��u�)l}Ш�����h��b�%R-R<����[��I%OgU�l��p�V��	i��]�n�֗g���$�4�nr{�G� :�4���W�!��7l�G�4D]�P��5�=��?�QL�T���V���⃋B��11�͉`� S�K�XK�򥇟0�0�y��tC��T���r��0�Tg�8RW��8�/RiTIǌ��DI`w��>+_x싰q���.<����6U�N��-�9��ή*�#I�4[ʨ%z�M%[�����0��GW��q<��j$	���u�D�l�M���&R�U0(��_�R��o�
)�ua{�L��A��_ B�"�`���e��~��N�����7��z^-ӻ�����
�EY��@�G������X��m{�O8�Tp8���1���q;���s�(Oa$#X7�9�+Epj�'=�X)��ۚ.��z{lZv7���L�2��5G����.�<�X�-��q;���M�Fn�,���h�ڸ��˖V����/�Y2<�ʹ�ʐ��0f����!L�(Va����MD%��D�|��쀉����(Ȟ^[��Tp�[u.�!���P�����ce�X���ڇ��OGJ���a�]��<g6��4n�5�gq]�<���B��RL���f4�_��bP8s ����ӹ�҆B��r��U`�Fp��ىE�s�q_��� 7�Ν���{u:�N0t���WH/�w���C6`�)�J���uΗO����굂2�}}8�^�yB�����h�^`Rh>���n�g/��ʉnݕ�8�}u��X������:ym�0��}l��#��#��C���Lݓ��D �΋���'�b��6���j�K�c
�HD]�Z&0�����n�:}��!�:[[�Z�P�i�L�%M�r�>0�wY�~'�����O��e����嵣���k�V�lTW�_��ȿ����rBC�)��}�S �U�z�p0�� ���>G2�F4��em���Ψ�0h�]��6.X��#�T_y5͛A��QC t�-����I30Ii錴p�~}��,�d����͍Y��B(�j����z��Ù:�%��c6-��{T�����J�ۍӰ?:�[�$��H0�AT;�,�p��ԓ��F 5+���f�}�1�n�p������9>��$�C)8^4��p_e|�v���"&�N2���rDr��ߘ�[Y,�P9`�>-�y��-�I>���1�|�a�]X����W�cϖ3���şX�+�"�oZ�otɬ%�m]��
�ہ`�� 8�݀# ¿.
��z��8��mk�b�\5�R��W���h��0-�<��D�2���*��Ki��.V_e\�;��t����X�:�[d���M�C�0Ş�E�/����Ň}��L�?/��x�����"%8��,t.�nXߎA�Z۵LM�ŉT�Tg�/!��H��D��qĢ֢���� Ev��)��E�G;9����h-U\������������SH��^�榉�J�'O5l�RA7d��y�n�7i7iU�q���t�2��yG<T��9l�o����2&͐:��n+�$>���8L��zJ���huJ@?�5��:�����i����D���,bnO�h+�x�#��*�Bp���9a��II���r �)����w\N��Z��^2Rko[������m������1>S���SHRj؞��~��$��EB�P3�^�Č���P3����POex�n���8��
����c�Y)����أ�Ds%�;�ז3��k���u�j�2)ƛ�u��������ۊH�	K���7!�p��us��/�y�v���i�����l�t�h���r��hP�P��{ >�U�f��ē�s�A�|��R�#�*h�s���R����w>o�^�yX������?�	��	%�F��F��� b��d�"M��bY.&�F��K���f:W$���Y�tB8R�1٫�ܞ�A�0R �>�������k�&'�v�kA��?�QzV׸�,����S��4|�B�"�uԝFPI]���ņ.琠��e5��}� ���`�w��.�9�t菾h�8��_c)�ηC5�B	�['�D��x�fWA#��{�=i�!��@{�;>c���q��;bXeiY-]!�փs�X��NV�Й9w$�!������	���`"��Js��r�Ӈ�Y�>�l�/W�s�0�"�n��aq��i�:׊4���Bi�G�#�S�f��itB،	"G�jx�`�K"�����5]J'�y��Ҥ���񟙣y���	�b���v,�[l��c�a���+e�$�y��-*�΋��L�D�ʶ����GA��Vz%�3��(���U����P��X$J��s*`��
��'��|��q3Ӣik�޽����\nB�0z"|mK�9F� PO��h�>��<�n���-�G�#�ςM~g��Qk>b@t�m��~������`生��<8��9�D�����]f0ꟛQrJ9$N�����K��P̯%/<��C�ۄ�d\-�S9U��<�2}ش�t��wВ� ��c�F8 T^������=����@N{t��2Rl�4=��(��}<C����>A�����}��*�����[v?��f
�Ռ���U{¡yz�?�xwl7I�sL�,�&��G�{���Ie�ks��u	���H�q.L�\J�O!ϑɶ�� � ���̟���R�a�qV�ݲ�(lN&��ޭ�Fz�}6�gU9�o�0��m>�F|���z��7B�Q�~�X)j����|����<���jO6�&�D�F�ŤcW��|�����l	Ӑ��j��[_Dd��%��8\Bl�q,=�!Pq�ƳdL[���V.����z�K�};�:�^B?����i�o��D�.>J;�� QJ����u���җp8�W}�p��h��򿬪VPؒ����+�7������y�<�A+KtJāƫ�� ��%?Yy�K�~����^ep���a�:��M �Ej��UrP�`8ndZyےk/q�h�����U�:2���Ԁ<V�#?ҫCz�P��FJw��RXn;(��-w	(鹱��5)>+�/ց����'Yyc�^�����^�����|T[���zx����xE��(�\L!��P�f���Ճ7$��qR	�v>΋8x$�7'�fwF"JP��r_��Y�T-��(�(�����mz��1[���\�I-b����)���+�;&��]_�S�����-Z\~���e|�����S�\�܋��������[_W
�^��Y�[i�p5�p�M}���ɒ���7Î0�6!}������f�-�s�b���� ��������N�)? �,��'��r�"B=.?�ꆉL@�,����xB�[�
->4�uZ�'m��ڿ��>onz0"�� B�9٣�̂�q��]��%L�:�Ӛv$��`h%-&��m�-�.����X\��H��