��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t���������P� �N�3��Z�oihQM%?XH&ɜ�S.�Ƚ�֤�x}S��O�c��q���dY��!`�F���ۗWogj���,�Um6�7A�-`Ǥ�de�'�Ӹ������������!��;��vs���L\�9��1Ԫ��V��@I�CD�u���߉9�G��Enݨo��r��=��1G�q������L�_@�=�̞t��{��j���*��dB��z[\�J��F���l�ktt��4�8�eA��,�록���Yi��+.�"��Vۥ� [�Qb��*&���C�H�L��C�z��J�>���r�L�6*�S�{]��١d\['w~��2J���UT��͛]V�@�����)U��]9��(*e�k���L���.�1�����
��x)s���)꽹R)�t���'	
�x���Q/���	�jx��70��tn43��������V�͚���w��>}�?�T'(Xc\�wҳ���[�0/��}
���O���
�Ȭ+��!�O�D��bc��U�4�D&���8u�`)r[5[y�0i��jβp�^��ӄy�jz	ձQv��'���8�� �2�o��1�N��(������R���݇���kƬ��Ųs�tZ�����Y���H'�<}�Y�h*m sN��3�D{sq��<�V��L��e�Vg2�E(s��"�B?���G�3	�S��` ]uS�1��CI�̀6�d���7�h
�̮��e�z���1F����Z�z��O0u����&���A����>߽A��/�D{J wj}O9E�.�8�Xb�g�;�NI�'�ڛt��xW{�XF��c��T{)Y�@�"��T�G�����-K�iA3�6���l`$��;�hILM�#Wm-��!h���X_�/-�%�&�t�Ed~�#��]f �0B�% �T��JhT�0�7�>A���Jq��/�R�g��.�D7oz+����o��B�c��~��4Q���X�e��G�S��U�,��O��=~?�{R,!���T�8��#)�hϽI�[���4m�T�(b�Ԡ�f��(�π4�:�H&�I�L2��d�Z(�+֫�
���[�1t<)�:�{0��l0�Z������ŰF1�֛���aٻc��\�1U}���4S������p�T��W��S=�x�L�.�z���e����H���)ZD�1Qz������O��� 
}�fLem��C9a�A
�Vh9�C�P:�(�k>������`�pu�6y�ْ��w�a��7/��X� ���!nN�a>�;n%�Y��ק}�;����*�'"�����7�*��U��6�����sU0p(�@�W��6t{�"ӎ�Է�i�c'/j��y=���X˚�K<1��&���H��ܩ��8�%Ao�z��/os}�9Ă*N����^�@����$2g�U��S�
*y�h��2|���Y�Y�3!��/[
8Ol{ps֒w�d�Q���&���K �X� �q�Ќ��7�#{a!sc5�e�7kt���p�#�~�=6���N��" !�@Hqk:�2���Wq�	s�O�e��a1l�YQ�}���u�p%�b�i\���<�ե��	��S��-n�H�7N��*���oZ`�{*h_��S?wzz�×$7F���~� �΅�L��`�"֣�+����l�A�GK1����Z^ǯ�nB2��`�I�]P�B��hp�<~H�X��H��V06��5�I�7&���wr�C@L�|>�\� ����(��j�D���o�J ̢��D��sN퇫��D��u�^�ڙ(/�C�MQ�fy��<��An��"VP#�P9�V�N`�	H	@�� �fQ�}����z݆݈2�b�kV��m�O�ZQD��,�R#gΏL�$k��vi(Z��P�u�/g`K;���4w���ߵ��t�V�ӆF�Z+�dUt��FP�ń&M�o�6
٦� � ������qP�-Z9R8���,y��l�}hˀ�I{�L>\@CN�ǒ��ej��Ɍ�(f5�_Z3��8������b�Z��3�d�ә/�Ƿd�;;\��P�Q�Eˮ�+.�jr�>�E|����q���~'��|�_#�g-o�+���K~A.�c$w���!8n� ��Q�cB���-�����&
��`��?�ZpNCܷ6�9Nߋ0E��z���ڛ{�O������b!j���Q$�n��T�K�ҫD�9�:w5*�MT��0^o6�;jp H����D�H��gmk��@Sq1�����D��a�kOQ�a�M��&2:(''���5���G��a��1��@ǘ�1��������A�\����
4HD�k�����#��?0g�uN,Q�ָS�u����d�?\����)m�D{�L�>�ࢰc�r]>�X]OBCg����4X��k���A0!u�<z{�ŗϟ����v�ӥfS��� e�҉V%�jB�n"����9��=z�˳"��CGk��K�K3��J% }���0�JK8��nW�5���1�6v��-hGqì}e��l��c�	����"[|��B�l�	s[IJq'��d���<�iV���@˗۳K�Էٲt��V4�ïK�1Z"*5fo��u���H�g�>&�1Ar�������2_��ￄH�`'�D�E@yebE���M9�IȆn��k�xjP�4����N�0?Tb#�Ǒ}v6��5�2M��@vc�m�/Ck8������{�)�x��]��В�(]���|Gh�����#��	���^�N���8e0y��r�A���]�E� G��V�QTpCJ60d<�&�l�[;�Y4���P���#����B/�!�g���:��:�g����d�уQƧM]��z��_�@� �T()����J��������`-����=+����6��MtK]cO����͏V�9a�������z�}����{�>�Y�,̀j'��"�a�g��(_@<ȣ_��}x���L���ߖ㐀z�]w8�c�H�ReY�xQ��t��J�+��@�q9Dpޔ��,yF=R]o��Q�n�}��4L�@#�y苔X�LY��X3���W�3+�|�kZC���W���f�4$��A�Z*��i��nI3�3o1��\F!�=|�}�q�yP3�҈����\H� E��3"���{"��ob].K{���/Ӂ�#e�HT~�������:.���1誎S��O���6����O19;�����f,^w�� [?�w/4�
�����T�h!~'좰|0�z�#X�3���:L��B�A�4�/I�&�=5dI��R�'H�֚�腣Yŭ�q5v�ȗ���Q'�-�����/���Iv||���A
����YM�a
�#��>J�a	��gIg2Ͷۻ�pG��F������|,P���B��]׬�y�d����.�;�F0b�w�cfմ��ЧDO/G���{��
��f�0�N��ak�D4K�z7zP�Z���B���2)2���q3l���CsG�~��+z�8zm�i��/��8{�R)1k��iu�x�N�k�F ��G�٥Vd(	�E�	&W��
�R��D�ЏRqІ��敭�o#2
�T�0L_�>�ф�Z<��m�iG�E|e�Z9U���Y[�eq�z���t �5��	���u%yo�3ޟ�'��(r��7��$�Fm�힚��dD��L���Vj�%������<M�Q+�d'�م�ُaTNCu����Sw���!�/��������@�<ab)���:A�ǖS�v���gj�/���.K
�9U�S6��$��X�ʹ �d�˂�kD@�F��8��F���x�� 2ǦS���X���4�����K�R��|��N�,�<���{,��	/=��M�ޚi�8����G5���C>����ũ�y��qC��<�!+N���=����/$t̞'�Ҷ�V�D��{l��t����wR/
�C�yU��S�8�j<�-d�s��4��x��LL[s�)s�3��$�J4�wdw\i����HR�j~*���\k�db����tf�"և@��Z�;?�t'�/a�d�t��x
É5� ^b��m�)G	t=b����s5�'V@T�pߺq,���s��	��8��NB�ģ�����4��y���o��c��������(���&�L��`X/N�4���5%���<���WRj�V�� ���Mr5�Y&E�
���!�'�<jv/H؄`b��	Xg��kp;�A�=�<�{��� +�5|���^
�爐NK�:�G�q5"P0�l��,j_�f5j��ˌ~u9,7؊z��d��r�J����P
럍ʿ$p�fŖ��[l�!�ao���xQ�H�ÐPrE����h�gM�������5�>HH�T�)�׎�rFI��0���BxY\�=0�q��8T�0p-W�E)�ϐd�q�7E!۝�Ǡ��3��;��Kː���*pύa�[?�L!�z,W�V�erʈ�b;G>>.��+�IX�Ϻ���+�oy�#AD�I���)?.�=pN���)|�����]2�`�z/�L�%���t��nHjWܙ���/�_�+4v�>(5t�w��y4:��`7�h�I)�e"�;�9����ؽU�aD�I:ś�Z8�a��鿢�3��n���|=�69���)��~�5�xW)��`�/��3��T�*�����j��f���Yك|s�w
i��(���4�K�}�;�{�d����@��Ф�a�k7�c~���G��G�R������������pF��fR��&
|mE�?J-ʩ�KU�1t�	��J��ك|Bb����<Љ�V�]x$�v�g+�9�;��E̎y'
��r�ku�YQQ2P�D���,c�w4l�^�jC�%�5!#��j,������}�5���[dI8�H3TfQyQ�1��zkDfF�VG씧����x�x>�)�s�M����I��>������V�B��U��3GHw.F;�V\�����kH>�Y�CE9;��'
Rnn��>��U�Z_hp�墎�3XO�2�����>V���nm4�f�	�ض*|�@�yP�ButT�ƿN��[�Y��o94�娡�*�y;2�(���E�����Ar���˭�Pi��Y:$1��l1��{�ի'��$�ah>8�O���'ѵ�t��
�����b�D�0�g.�RǪ�]N^����z�)�f˗5�:��Ra��ȞN5��O�Z�7���2����ú�u��~ � ��T�08��/6���
'�n����vpl��x3���p�%�-��zP���%�+�n��P�y�Q\45؆T���c�Kg�)HD�ҽ���k
~D�'�9����V��	ホy�չ��Fr�lƁl�#��f���Ж����S��t�h��W���<��K!��!:� O����:a�V?�߄�(�}R�3���Jql��@K�<���l<6�t�kL\9���)�d&��+�����OiJy���wm��p=��Y���h(a>��cr]�44Y |:W��tM6bfu� ߾T%3���j��v�m�1�����uc�w=��1R�Q�������zJ�|�(�R.Y�0�Ex�w�1���f�`��� �,���a��z�Q�J�e�P���eQ�v�.�P��Y��ݷ�JΤ�0�p�bצ�֔QԟL�>���5�#C�t���r��4j��qFT6J��݁��c�QZ�_<��'��g�,2�&��"��O;e=�^����|G����(����ylN8XU�!�������ӌ0Li����W͌:twUy(!0�x�K��9D���C�_�~��E�e��V�$����>�״����6��%v��6�0�q�>5 �[�0�-��뱾�B�9	�L�قSEx�p��9���O�)@5d�Y�eA��2����ݪژ�p�9F�q;��e�k�b�[Kó=|�j#����#�y8>xVJ��&�p�i�q��z���b3����S�%h�;�2ŗ��ғ���s;(M���5V��݄1&�D������/%V�j��� �ilL�!�ͭ����>:�y��u���a���s��_��"C�J�J6��˯Zx�l~�����i�ħ�c
M,v��jx^Ul3��my�<)d��q����tmS��aB��#�|�Mq�vy���B�iK?j�ɧ��P�T��# D���v?�Cx;������j���%�U >��r �]Z�p���p^�ˊ�9���;���U{�^rۢ!�&8��!}�-�tAI�LM�,��q9�n���Z�(!�S��0_x+�2�u���������z�7鎾B�(�F��5�|�D��[ɚ3��j��!zU�����0G��~1��d��U5H����O�nr�PY��t��}��;�=C.�b�Ȍ��چ[l����sA|\�cs	�ۈU|{{%�ꨟh*U�� X{	����@g�~�&�(ʬkX�'Vb\�F/�৴��Y��r��/(��q&s�4Rg���ܔU�1_8�L��{��W�?�%�iԧU1R$Ya�	3>>��l�)b��S��B��?D݉�f���q�H��/���`�Hg����r/�+M��ϥ`��K�y*�P��F2w /b�t�bA�/��͋Z��e�*?cK?X�M�,g�k��I5k��xѱ��q<�7��܈��X���o�>��o��ށ?��9�-#끄�*��|��)���ƦO8>�)���\����|l��:��2������3�n��Ϡ_�Zؚ�
����϶��8%�˝wz���>SF�WmݞS�S������y���m���o��Pا�U��HjY-8Н1���6A<��m�&0mK��]Xլ�r=Ġ����K�<�3*$�EKm�Q��w��^:� ��,���l����Hޜ�Cvp�/l�4csA��,.Tr<T�����=j�?�0G�=�3��F�3"�[G���t�;�f�ٓyp��vtޯ������ �@�>�������]U����'B)��*m�`]G�u�t�ݜ�S�o(�!���R>�;	��`�3 +A�v�W�7��,N{;�{�̖�{�54Fr\���+�q�'�KI$�ȯ��[f+	ݙ�v����]���ҬS5�0� >k��Msc٣�#�->o�/M��Af6>���c�1�&�y���b+�/V����'g�JwHeڦ�����A�=�P��U})�v���L�����m��W\��mǪ��2�0���9�e�֏��3:��1�ǬIRdd�c�j����T ��80�_:��-�#�u�x��bA��!�NO�X޾�k2Oq��L2Fc��'������J���JG�@�ˁ�lvƄ�J�~�6C�<
:��`��Zb�(�(�J���-��m�R�{����y�O�.qP~ëbٛ�MaC^S	�N��za��,-3XPe�6o��o\����m���<�?��fPc�B�n�����l�VM=�Bވ	�>��n2vc�$��'����iA��Q��D`/W��ݿY��ar4����w@��A���)�`���7���0�䀤v�QifL����xr���|L��R/��yn�9�A��{��j0�US�1dI�Z�������յ��5���̙�ɽ�F$sC-#PWx�w��ԧE�kD�N��X��HH���٪�3�8�oc�o�c�`b�t할/��v�|��u;�Lh-C��H'��\��vІ1o{5���,[������L�s��N�J�K�wL�:�O��Fx1;/0�͒?���I�F�Ì9ĈF���'$��VL1�'c�j�Ʃќ��W�&�NN��u�*���Q���Ju�*�����GN+\��m��̋�ѹ�&����&�Ў	týh �e~`(�k|gA��gy־���c
�kNiLK}�4�p�r�����?b�T��ؑ܀�%O��n�ƻJmGu~����О|�d%��A¹Uh�k[14�,|���:�y�톂Ua��@OK�4j�DBy�5Bۇџ�c�/�lߢKJ%��3�@��j�%)cFu�Ʒ���X�a���I3����������l%��U��2DU�����r� c
���e��e�o/�nPʒM�Ą��cZ)z�ś?
�<`�Y��ZN1���{w�,Ͽ�Ϳ��7t4,�%�G-�p�;;���+�9�����;�`��*��+�'��V_ڸ����d꺨[�Q�9�3Ɠ�.kZ�
y7{�g'F����d�l�Nvf�a}��1������%��!�NEL'H;�M��+�ZgkoG�vm���]bmm��ZWm������a�J2A矂jVM/���� ��y����r����;�W�)L���_��C0bc�-�z��jc�������,i���JZЋ/��'GD��P�ި��/6��ROƐ��sU��-��S�������V!>D��H�}Rϕ��>�<Є��0�'S-��M�<X���]9�L���ѫ�Ҷ�J`���&�QnG���D�F�;����@�Vϲ+�C�i�Z}�l@c<@���t��%V���ļ�]ʿU��Ԯl�WVAl%��T&���{w7 $g[�h~|A��	b�iiFy��|��~ =Iɒwb.�j�G�D�]c��#�E�⁒����Q���:�9$y�#�B#���s� .�~�Z�1�`d�#��M�v��=�\��"���k�����A�@����a&��M �ҩ2���Zm��������rI�v�����K2s����5+{{y���?ڢVԮd�u9�㑦ZW���Gm���I?n��$��@G�˫�p!��Y��\/Uk�G3��ǂ} oYT�w3��Ʊ���WݖHr���_���:�]P��#���^ֵ�$ʝ�2j����t6��:2���^��2�R�Y��]I6�O��A��7b��ʿ��D$
��H[���u���ՙ���;3�?<vx-��|	9��a��|��I5� ��?O^�hE�f�B�jx�q��!��r�*�tZ��Y=t�Z����G̿'׮��7����`�/�|���B&��W��	�+}�Nӭc��5&�CB�Mf��a�2�޽	L~{�2b�L����t���1���0^f ��tO���Z��+PS[�Ò�A�}�̴ZZ�s�E�����1<YU�I�䤗��%��H��op��u%{�y�N�Q��c��ʅ ��ԕ����n>�n��:�Z����R>qY�*JV���oEYq� C,Z��g�D-8�Cϳi�z�e,��Na)�;/�<�J6`+ˌ&W��PFʤ,�+C�]Ɓ,�t_	�貛�K?xYeX�t�=G#���bd�f��c�%��eB�  �7Y��:�O8l'_JhK�;�Q���&K��<�O��Q�l�����ҥ���?�Vl����1��!�cԓ�Ю%�C��g�C0�	�P�C${%lc�)��i�
=3��H���[q����e�+|�-��Nw�-��uh{^v{��D.��F?�����%HK���~���;�](G4B��g#�< ۓDzS�P����D}zڷj��*d����3����>��Sgm��z�"��S�>��t{0Fπ&�cN1*8vr.�z��򈜒��K��5���&��Cʀ��������yEN�:�w٥?'���Ѹ��3��Q�#|��3��7O�K�DLc��J]Y%,��0�!�v-%Yz��_�,�z����U1M�ꗋW�u:�����Q����b2�Nޅ�3��q,��Qa���Yh0��H ���$�Yh�q{<0��ݏw�u�(���*N�o��1MR��4����qQ��R|�
���Pk�e�L�~#���D�5g��aϲ���N�j��E�Q���l��t�Uy��Rc���|�#��!4h����%�W�@����d s5��y,������%��ɂ\j�ֵ9'	�����]=U�!�d��'�u��E���`VR���"x�H��6�?��p'��8!:	���Ĵ�����W�>6XU��
��"�.W��M}."{+��B�.!��	�:�q	��BL�j����ƥxs�u���&��+�NTe�*�5jV:�`T��v��'���4�kZ�2���Q�����[��)b۟ri��:�n�<�W|'�ˀE���T�����Q�cEgg=ڛ�JJ�+`�5�YG!�0�?��k����
�+,��h�BV�C"���&=63G�0;�	�P�K6����^�B] T-ׯK��- t���Q��0-����]r�,!���@и�Z��#���o�g�Z��IN�I6e(r��̹��n�Y�6R�1X7#7���g�xWB~|�{�&��wFԅ�/I�!bu���;��L���anر�G���ѥ7$b��>�_6��3I��^���l^����F��:_}�D�^� W�Y�qa%�Ȱ��.ꡱ�w7|�V�Ŧ4$�}�|�r�����D��A��"{A�)Y{�c0���kIt��!�Y>w�o�A
� F�9ƾ}(��	Ŵ�d��iY vCV��L�`�ُ�(]�v� |��xU�¶�A�����]#{(�j^��M�N�*#g��D�O�x��Eҝ�/^��(S`=3��?k'�?�ُf�Iv�B@��12���R�y�p��%�eD�IoD�W�/�׳:�������۳}�ۂ︦Eܽ	�*�@s-v}�Y�Ws���~cQ�
�C��^��ZH�h:�M-���8e��>���λb<8%}�Ҙ���E����~̡�#��ƛ�9ǌЮ� T�'MG��a����d�7�+Gm*H�E���W���޲��NY����?��EZ���
�����k#Ԏ��*X��#*�z/�⿖�w�z�
��.�<?�s	e,�X�BB�$:�ڜ �sV�Fg!K+a�7ˣ�Xy�V3kP�����	0gi>8m�Y0ssQb�4�c�]�Uf���O�Ω�������E���Н4���M�Â=�vwu$�����(N>���1��ЏǾ�)��]y����ά��=���Eowr��*ܶ���Pf1J�a_y�f=���=���z��n��X��U��@tΚǓ6	�}>e4�L�N�;��Z�S˰^ϣ�2�k�_�w�8����c(@���2��\��g���'�"�=�m��@�&Rf�D��
�a�����}�U��0���0�&\?�5s��u)�\!���L���mk��rݾ�۠�r7�-���W��N�����1=����P��(��,�+dq��	�Rѩ����+yZ`��G,ҬDy��F��"R�U���+_M!���=��M�u���R����9�ဓ�;�M�$#~D��ḥ-���hxS��xnQLT�4�������s�*h��RÇG�B�ff���Ԇ���Ee�t�����o���Ÿ�J��H�Y��A��<{��+D2���1�|��5"0\���װ	I��/��³�S��|�W�;�O�;l)<g�o���B��]�)�C f��\zqU6Ɉ&_���f_W���Ҁx������+*��ܛk����l�ܼ����Pי�T�ۓ�U��ѵ)_+L��-�M�j6UFPm��H,�r�]�0�2�YH�*b7PT�`��@�Σ��{um��B�ĠAy��Mq~��������d���f,�g����GC�������ܛ��G���8Yq\�L�?�X��1�;/Qg��4��1�%,8�
T���v�Q'��s�h�?����.�,g�M@f�A�*7��,:���:�WЫ0oOE����v݇�@����`K�X`K�l�8�#�����5R�Gtw��Ɂ���Ф��QP�QH{?ԣ���Ҷ�U,��.�}f��ˉ���fg�G��Y�z���O5��Z����1Ç_	�Yw���x�*�i�5�\`ې��̢��֑�f
?���_�a ׽���������z�\�Ϭ�W���ߺ-/5��P�.��ʚ�~�3@F�/iH1"�▫�>^���d�-Ɉ��� ��Ѽ�x��ALN��t^=k���0:z���{�t	#t��{�/�/a�aE�����H���G`n�8i������+z
�h@8������<	�{�^��P^[f��ۜ4�"l�4yX�F�b��BhxL�;(�� ������FVX,��k�Vń��o
�Hq�>�H	���t����i�v��ÍY0NMYf]�R]�W�5�&�[�N�x,�����+^��/��i�w�{�}㝎wE��� �j��&�$B,3h>�pp������<>B&X@�Zmw�YIO��{ʊ� ZW���Tŕ���q�Y��
+�;�rԓ�l�������Z&ϊsXQM$��~
���J��BI�6�5Z�)�U�.#���r���X���	At��](�sՊ�����-�?��)�!vՇ*~8��"^��'k�ߘ�x��c�`���(���JR�����O�Ր� ]�WБb���Z��'���v��&�t�h9�Ɂ��|9�k����5����u���Ȁ�}D��ޢ�M��,�$wi��slG�I��<�'B�z(�����,%d�ǔs��C�G�RԹ���?��m�c���ê1٥q�ߨ~T���?7d&Y�"���ec��g�$1y�km��L�I��G�SR���
���� Gw��N��F�A�*���_�Y��%�ߺ��O� �N5�&P'2!��ْ�l���\�8�|�w�*���i*z��fB��+/�-~��lA?d�1D�l�
b#� |&P9���i���H�L�l%��	��)�:f u�˽�8vzH�#�fDv��i�OǤO$�Q�l�_�����e�!�q�A���5~pI�SA_L���2	i��\~Pzp����|`%za�
C��P��3�9�U���`VHE�\���o�NC�8Qv~�6��d��u}��JT<2`�($E�q��cT��űM%��m��A�0q�ϱ��-�$��*���;;�		g"�ѕ�j������.����)t�tL����L2 "��}�����a� �4h,]]������?���}�SoA���FqJ_/	n���&�wEY�Fh��1�7sv�s��7P?�ּ6E���n��?��<	-�D�/�������6��c���v)Nu8C��aG����B�םW�ŋ啄�����	���n2���CE����^l���	}���d&ܾ���bm�ί�XI��-y?���̑�d'd�uD�l����qK:#��O�;���&?�ɶ�v?�D4.󘹟n��iZrJ����AٝR����ަ��pԕ�f���V��o�6z"~ϔ.?�P��SK��"�yuzv+��x�|�WvIY�K%I���|{��e�B$�<Zv)eY4��4�4\OM{��l�?��=a
�Q��kr�|�}����D�wK;����F��7�J E�b0i4����M���ד��R���d��`��S���˥���ݢ-��?�O��P�K�GL�x~�|�6/�sN��#LMe�Y�N4��o��b��;Cc��p�� O�*_ �4 E�M�Nϫe�$�a�Z'�_k�V.���)��G����_B��#��e��HS���Jx�X��{_�g[�@Q��4-�f�Z��w�@E����ҷ����ڿ�*"�z���ɉ�}hML�TS7S��0j�;%:��Fc �{�N���}�H(��?�SFװX$D�͊���:�H?�i;ۛ#�lj�8O��8�ɯ�r�.���|�x��c�b���<<,#/�}�k3]��8����`��ptޓ���)ފ)��֦o�Վ�ڿY>��ԓ{����$-��;��Ne��x< �Ҩ��w����T �N_�Kjs�U��4Fd)���{Of2%�x�e#��!�0��Q�-��t�q�fO���^�,E�U���m���79�Sw����ZY�D����|ގ��R];tk	�[�u�|ޑH��.��$'�cI�����ՙo�4->�j�ȁ��������j�Pw.�1�D�CBN�����=Z�9q#Pr>�_�],)�v��c���5봪{dB"��Hq3���o�ò���JcP=�,�0���ao Kgff(�$)Vɧͫ7��v��:��?J3n�o-�i�^&��6Ie�h��?5k�
�ʣ�+�B~L1={|�QĠ���-�{�I}��B�$�Fע��&��x�#�326Y�jH��K�\���� La�S�$C�QJ4������pS�d�6ٙP��m\P��<��G:}�EG%rL���Ox`<|��?x�*������}��<j�P��Q�>�*�DT����u3,G��>*}���Й"вM~a���Ӄ�^��nj!���:gvĸ�PԴ�����Y�;Je�i_�񴧥k���wq�С�+��O�؜ٶ�����P��Q��nr��B����D��*�,�T>����
�k]�ĳy�,8�����{vG��>��:Ј��:0n�dƄ�����.�v+��Ë�&Z�iN�_��L +DĎ��K��O�d�-�7!q���	�Q��C�#���%��V��e3T�������]sXr�>�2��eߌ%�t0h�yb.0��ʦX����|���aI;���A���^����Dc�mں�^���b�'�z���.��յq�4�O���σc9.��D�����"�'��M�A�P1���!�1g�.#}�.��B&����큜I�������N���k�ω��ׇ�#����!1�w��[�T�%�����%�r[5���7�L'�t�\�D~v�U��Jv�H�D/����
��i� �`<�BJ{6 UQd��ˑj��� �pe��9T�Wq�:����J�W�/"/��c����p=|�����������<�<�6iؖ�2�hIh^�U��+uTJ��
�!��bK'z:$���Hp��M+���e�Tdv/�u<|Vpkٴ�NLK�z���E;;�%�"�����u!��<M� �b�D1�@R�/=��{�Ҝ�.+4U?���Z���Cn��[n�tm4���v�%�"JľuD�d��B��~��폲�Z_x��J�;�㩏L@!�c7o��v����.,Ӛ�(Cf��ӷ[Ӕ!�q9A� �8��ʪ�E���������k���]�`Nm'6F8�����p`Upw��F*C���Glg�e�1�&����ՌQ��2$L�Zi�W��f�[��?W�е �{�W�����O��~�'�hf�p�����(��U�kW�y���: ����5��-E�:e�1?`MNɘ��B�b`/�ܷp�2�D��q�94CQ���Q]t@P�k�Z��o.�e��+�M���@xX�_�h�}��'_|�AhN�M'�U�%ϫ+ъ�'����7�+��N^�7Ƨ�s�C�$���ODg�\�����އ���C�&�v�g�4G3�d�l����x���'�|P;���F���T�'y���Mpq�C���/I�-V�ע1;w5b�-����{4���h\G��oA|(�e���&���� Ϥ�p(��18[��yo|D���I2�Q����,�+�V-:nʞ�Vc`M�H�P�I9��36
x(536M�
��']X�Ť�y�O��F�s�
6����������2)f1���ңhe�µK�TP���X���ci��$��I��c{s�(�9�N4��=_͑~��M��(ŭoR�:JcsU����&���:v���9Y)0q�`W�|��,�ƽ��Z�5jD����8�t�fv��K�6woD��pi�NI��G%�,_M��`����@���q�e�,'ΰ�V�3[ 6u���y��h ��A9�E�7��tu������=�4�"b�f�J���׾ڣP��a�2�)��^B������G�@�Q��I׎�أZ,h�]b�����P'c���_�ת
���%�b�}PI�S���7?��Q�O��dC�ۨTv���-2b�DO�������M'(E�������^��Ӟ}�+H ��3���jjx%cIdH�\*WA��K���DYy ��lG��P��?,���IJ�\N@֪?ؼ>T�_We9j � ��Ld7�tS�رZ�4a��咏�k�i���M�r��8���8LR��z�k2����N��)A�/-�D�ڽ�&��.�e��E.�YA�ITaP#��d��P=�8��צ�!2k����4�#��a;�]bPC���S$�ZG��U�O�t�c��PR+]t+��Q|��f:��Ձ0���%}���p�0>'��Wr�%�i��W���,k���� �g �1����1��xk&�BK�n<�3R��y����-aN�2؎�ˇlة��F��Z"B����a��+�=$�g�����F����#����)��w��e�������m^��ܦ�Z��
�B]�/�ق��Jȃ�8����v-�`���W�����і@�J�t�k^�;ь#���1�IO�D�12��ZP��ޠG�r�U\�Sω������
�dȃ�}��*�ަ�6O*n���-�vh��lk��������$�����e	5�6G4$J� �#�4�H�D��4����}{*��k
=m�{{'�pN�y|�� $���H?j}9��Ş��/��}�F��?��}��'�I2V���r#�G�d��"�[�h�	s�┲�[ϱjQL�zaz��F�1IC���L�a���b�B�5�9�Q��:n���*y�ŵg�1UZ��`֢{;�D/��j���{= h�onUFH�xJb���ŌWk�ߙ�q3�����f�
�-� >_��>R-�&�t�]�6�8�W��¾o�����"ʌ����)�j���ke�4��e�Vuݭ~.���ic*~��l.�rП��31�UoJ!�0�q\��'��{psy\�3�E�ck��9ٞ�-i�o܇�eP�����=��'prr��ܯ�	x�6O���o�~�����c��mO�����e�,�t�Ņ��^��+S�)�;9L$B��C����S���8:�THg۲dyW��罧HFb֨`/�M}�n4J����6�=�{�z@Yv��uP�A"�9~zX�B$�:mY�G\�Oj���ԉ��@�YnB]Ϳ?���B�nd�v��j �ip��h�\K��qڲ���H�D��ur��T{PjHԑ��Rd�rEv��}._X>x��Q�4�O, �*���u=�"szy���#�V���`g�r�u0Yz~~�}����=��B���G8Nŉ���y��ɐ9����qJ��s�/�=+��0�ԩ��R>fcR:M\F��k���P��K���y]ag:ء��j_�-ۻ��n	|�������! �x����6Q�0��fU�O~��%Z��6�wZr/+&���K�A/`�"��g3��a�.=���@��b�W�0.�'A��:i���f����ڨ@��]3�������\��S�e.���צ��n|X)�3bC8��eq�6'�C�=�'�t.$������ŝ}��{s�A�T�������j�:�ȸJhHy�]�Z����-�E�n�^�w/�C�O���I�u���� �������loI�$�:���"�*mu���&�GW/n:��	.)��� , �g��>��B�M��;��,���t�ЁS���
��6�k�2 �M`�b�s�Ϗ+��Y�;2���T��k L@{=���F�l�?J�b�"B�����y(�9�)zT�N�$~�Z�lA�~l�}�v��=M�[�o��n�xC#@q��R!�-��ӷ��X��A�Zs�ʎ�W���y���*�؉��4�}	���� nȫ��l��W=�E�Ip��H�&ю���;�A���L��
�F��w�q�U��R[�t�B㨚j�0��� `�ђoW�B��%L�J޳��~�r �?�ŘI��.[)pʢ`�d"(�ns����"�wpW-Am��Z�(���^?-]l���λ���Pn��������T��Ɇx�����x{|Xy�|��i���������	<0��}&A�9��p�L�A�����	MMG�XX  ��(6dmz�e����-�J�uߌR�����(f{U����_�-{��j��ֱ�~źDd��x}!w�4�2R��NL��N�,X�U,r�Ƌ��J
iT�m��f窱�>� |�Z
~�#�ȋ�
�اV��p��e�`xpy�0�b��u�`�9?	�Rϖ���/L����1)��V��^�\	I$I0+���D�9ᇨG�[�I ^��I�Mv�-�*$<�>ӵ|ͺ� ��������u譜Z@���W����ʀ�_o�I���Z�[�)nUY��O���j��/4�D�����$�1�# �F%5�/��8�!�娞v�P���� �]�*�(LHz�c���:ЛLv�?����e#о*����i�U��eJ5+�hT�_�3�7��ѿ  �D�[����a���B�!��p��*��y���M�8̘�һ@i��<���!����~��޽7h�ƾ��_�E�X�rs�����9�@1�z�rV4��NX^�eB�	�Ot�A�~��|�� �Y��f����7�)FXr�97S��궧eƹ��tT���I�?���1"_�������������W��P�����A��;�(6v�;Ɔ���ؕ�ivDC�@�݈:EƉ�E3�������f(Jh�)H�;�}:J��.%��=	�1�:�$�Q_=�(�%I�a)��d���';=��B1����Gݦ����W��2���^��>�B�L����2lzaє��T����e�\nf /�'FB��j�-����!�!��'Ee<�ޤ�������~����T�a�9�I�U���m]�bʄO%���	J��h.��[a�^>���+�K���9|�;F[e����4�fAK��$[O��
8B[�W�����R2�&?�m$��{~!`�l>��=\��ƠK��H��d>���/8��Ca�ql͇5RD���_S�c�7U�v���ǁKn9;\d�F�Ifs���FB�J���U��a6��'�%�@�"W���5C�*]��E�*� �7.�BG���Bu��҈��J�����
��xFr�M���A�K�@��tjJ�Rh^��\�������\3\�|d��="O�1GxKie¤a(|�'vsh]U���_��0�E�{������Te`eJ?��M��
-�`
1	��2+6 �	�H�F[��v'm�rc�t��<s�7޷o��=ʎ����*����4��l"�E��y�4<�̿�� ��Ǵʉ��=m�������7�̆�͞ԉ�S�n�1917����{?�KA��/�:-򢡆�+����~(��̵�����rb������1�*�5�P�z�"*��b��el���$�M�����4-ᔏ�>����E&��D3?�:���nW��z�`T8R�r��Y�z���5)�Co����+��H�`\d�M��"7Y�K��dz��`�����C\�A'UPa����n��˹�^֢�-Y��u�[�� ��4�}P�-����~���tɏ=�)*���0�`�^�`-C.�5�G��3���)c�!��
�-a���3*r� ,Ʈ:��	��[�)dM�_��C������o���t��@����ٯҼ[$ϑ�3}6X���G/@�^g���79Wֶ�����5X<��鋧���M�u^��M� ���'���mv>_W��(?�R�>^��:Kq	�BT۠�t�|_ K���FH��Q��S�5@���\�����W!���W���(H�Y�^�?��Vm���?��5�]_d U]E���ӝ&�R��f���u]�2r�
�A�s������&{�~�x�S��rn٤����X��N~�1����ge�j��<Y�Nw�T��UR�w�=�2D�k��_:i���gt�]�'sl]���RN��s�+��3^����'Ǘ�m�U�:�!�jJ�J�mIFM7�R��,��v�N��5��`�TO��rN�����{���~�&��-%LP^Ku�(�5q$�!i%b�@f������ZVt.��]��ϒ�櫪���F���4��n���φ㪲B��(Uh�mn�xc���>0���U}h���Q����)�Шz��҄�*�aw��$+��Wx��1���~5��A�Y����������4Y9Q��s��u�Z]W]m����/��֫I���"׺J-Y���K��ߑ⁍~A�%a38>�3��,H�!i��9��� �]���S���9���v��$;~��KJ������-������gE�It��[��U��B��:��\�-�+�+�}�a	q��.n �]g���O�8��9� ��8N�{S���ɴ���K�H=[?�@ß])h�lWM;�\�H����7����zt���ڟ7Q��at&�N�f��+:_��[�c݊h�'�$řd�ץ��'���Kj�
���b�}z�"��c�Q&� ��WM'�HCp��5)���ҍ{��n�
��鮁]��+}�VB��Z7u�C�Ϳ���?�;*��.��h���R�vV9�ޏ�GX?�yX��B��P�W[4���s����P$2?�l`#�L��nh���	58aPAs� �cRg\w~�+o1Y�Q��	�`�ϱ�y0�k��de^T(	Z��ϙ-�fӦ;���o`7�� Ǫ�᳟S(!��jFǈwo��ข��q���BZ�9��55Pf�!��c ���!�G`��-��Zߺ��yb&��8���B��=o{��Z�Ǌ�ZV:�W~��8r�$�[f��*eL8D�T���S��EYa!��$8�hKa��c��,���[��]k���I��4���c���12[Y^ZI�W߇*b���X׋O|��hͅ^׉�u���l)�m�r�B�@\��e���	��1�T��/�ߤfB�ٳn|sȲ ����t��n�K��	���;C8��|�a��仼6�Guk�TJё���\�d$��?&R�P���o�i�����Q�o)���֘��0�a��&u1OlySgHM�B&4NK��(��J99�̈j@�tF��^�y�;����`%��v�B�}@�+�mZ��K!Ke��xk�e��6�q�-2ǀY��)�0[⡵�B����׬�A�]���?75��uL��|Ĺd�u��eH+�#��F@�冉o"�
�z�����cE�yL�u�����%�Ws���w�a���)�(T6	[i�FT��O�lL��6�|��?�Ɠ�F�l�~_�V�vUZ'g�"��8TGl�B勢r��=��υ�g��1�Ѓ������q��?][0Z��{Yq�l�n��O�Ql�{��͎K*�&z�z οMN*+���ə̶�Ky���+c�d7�K0T��Rs�FG��O���>��놂�!�,�2ڄ��l��Q�e��
�1M����D��Ra٢���K��/�)t���r9���1��1y����љ�n�Z�̶�cs���~�u�V�� ��ܶ�ڄ!3�;����5>�f{�|T�K�lѾ{;]	<ryڦ�&�e�}|�
n�KyC��pc���]y���*jz�|�/�WphN���e��ՙ�X��F���L������nl\C��ό�z����Cn?�2+���L�>`�I�@���[RD���íw�����?|q�q�;���'xn;1<�/��M�d����Z*�KGU���E���ޣ�n[֫=N�XOmR2�\��hc�H�=s�́2�"�p+�<���=!da)��`�T�4Aʏ~ �Lz��SΑ�W�D�4����ݷ+';�Q.���V���y}��*���t=V�.�wJ3QQ�H%��Z�~+�2:��|3s���'6��&�ؿ�Bc���ڄ������xP.�S#��?��s;z�$�yIb���<�
@[�<)�s����~[���U4��e�[�JDE�p�� ��@�Pr��v���^����:V���*���^^kr�L6�i���`�gȱ�)��H1��u��w���L�d[l<]���xJ/�؆3��k�AY����:,ް�OTE�K����xCޣ���͍��C+PC+T�#/��dy g)�g�M�c����ͷ���������Gq[�(���8�� ��6�)`4 ;���"B^/j�7����n.����ʸYVS�ћ���-��ƥ���sR��H{��m��$�<��w�k�w%wnZ_L���Й:0�|��5?&Z�W�\Y��>?�T��'��q���jT�߶�����w�̪y�y��c;���Zu��d��:�H�@Uy��������5��c-�?yd�@�x�'�B~�B=�_Q�����1�H=�_�-��=�Ј�Dp����< �����0Y�1���������3l�'V��e4>L��ɛ\�`��e�j'���@4��P�����{��"�n����5!#	7	"T@Lq���nZ����hug�>}��IT��J["k��fZ��:=�G���X:]�� rMH6�{����B�DC-�)��EDBVP8#k��HMi�����K�Y�b"��+���E~]���Hm�s�5�ePj>��@<�O=ǲXy�-"�4fҧ՚E�G�ނ��Ul.�W&ș���|��ڔ��o߉��9��$�	��x���AS0� �HvU�U�2��_@�͉<���dH��w�vQ- �A(ʩ(�<	�����|L����~/�����}��c�������|a>�FK�Cv�N��ݷo�m�\ؙ�p~]l�*Bf����?~A�L
�y�S����g��a�y9j�x����2E��_5L'V�=�X��*"c��3�G�X' �Ob����-�~��jP�3e<ѱ�(R�Z�!?V�d�2��5����@c-��4C
�Qpr{�e��$p��z!� '��,�RW�	��xD\��M<�2���b\�Hˤ���G��Hk��
},|0g?Z�6H6�JE>�r��d����=�h�'�6Lu�$|�����?VW^�r�S�y
m�9)^G_�<o�J
�8��	~�8b`\��t��Q-�}S�g*;(4��H)�BH��$�m7 ʮ�=�u#s����2K���Y�7�S��w��`M�K����@)��KqIx�ha���X�`�D#s~��0e޻��#���2f��ߥ�BN^Bz�v��n6�Acp 뼣�g+���39�IY^���b/�6���&	_͚�S+���@桦����`�*D���3�{����ǒa�r��ſ� �	��\G���L�,�Sn\\�*H)r�訳ҋ��S�$��)��-�Ӿ�j$t2j伮،� ��z���!�Ļ)e>��C���P���&�,W�O��.��N�v�5�k:���=�^�1&���{�»
HH���/[��z
L�Z��� �El��o�+�Q�p�CmO�0��0B_wfK��o�{`};�0inC��[��n�2�U�nV������|e1,�	n����t�������0�ݟ�o�,�h���._B5�]�bP�����oR����E���5p��7@0�3��Mo�@�ݏ��eZ��t�:�F3l��m�+s�2t�K���)�z�x�1Kc�PF*�0������+O9�a{�	���Cך�q�M��Zl�Q�>܆�?�h�:|81� ���s��~�7����"]�od�ԭv�ש�6dUz=��v`��&Ց4��0�s�����\��/E������O����y�Wd���w���l�DӅkF�A���=C}9w�b5�&U�0��jrF�Js
���)T��'�I�;M���xS�Xv�䲴���w���==t%$����ݜ�3H<9�� 91�^��w�M���HE�:3f��jȥ}bd@4��G
�����������1�6Us�M����J"�bϬ	�#�l��ó)����y�cgf�k=�����&,�w�|
��\�)��t�?�7�=���p;�d<s���9��a����E�
�Z��E3K]$�]�$AQD+��:����".d��619�	��weN�8Z_��ב���󝻧Ը�5�0�'e>h�P"��#�@��w�Tk2[�u��2�ԕ�S��3,T�m��P*8�K��?Pb���aӰ��fW�JY\�	q��O��h˞sG�|�~72$-[�p��iQ�0?U��b�C�3+�n��'.X�M��U-�Y]��	N���Vm�`h��Ǽd�gBr��kA�3MxO�*��1����ω�B�[�v}��d�|��T͵���Ʉ����t|�y�����W��a>��h�)�o�)+T߾��'*����Cf��.M0���AJ	�'��Ov���o�K��uK��ji��k�����1#o�뵶���L��'s����K	ro�c�������)��.�r���%$-��q�p����៩${}¾o/S��^��z���>Fn�}�q��{98v�������g�.|S�߅���=-.�3V�yJ� @�f��ZJG�*�[�w��޷92�[[�uּc��0g���[���ݮk���
�rI�}�'"D�]��8�1VK�I�/��s d�e�j����o�i����~.�mU���K�^+!�>9��|+��`[C΂QKp��%x�?O��)�ɘ�#�d� ��=��"O�T�yM:�έ�눮ו6�A+��1��LЂ���/m����A�Q?i�����9�q��|4�e�����ut���>u�)nU�q���"���^z��X��
Ø�!*���~�x����Ӝ]��`���	d�F�:�@}h=�a,����v>h�}��*T��7l�ҵtX��x�}��J�[\0r�6�a�g'DOI�O9}��1��5��j��@ �%̓�o�n�E^��<�Y�2�@W)�ţu��"�Z�x��kk��f�ZE�l
�'�b x�RdrBw�˫f�E��׶q��]h��y3��!"n�ZnO����A�8�)+]-r�G�D%4n�T1eN���?F������m����k��=�e���}������0�YbX ��:�-�ǹZ)��e� �3�/�$o�DN���ri�az���f@����7w�ۅdυ��I��mj]���T�V;kkoG5��B���g��P�@"r �{`A�����g#R���/?�mo���v�WA8t��06L�5 �g���?�P=�m9�XF=R�F&�b�ZHF@B��F�@�췍���~�>����l#��Ҩ.i�4笳77�X��-��~jO�?2 �1`e2���F)���o�sV
n���l�1� 55��$1��%������r�N�T"�.��9=�˧ '�bvtp��c�f�a�_�d�K�d�m�C�i��Zn!\�Lkƙ�L5�;�� %c�Yq �����������ɋJ2|��j���:�1�|��W\�b-�9�j��z�UEOC�5�2��z����?�ި�3$ ̰M�4���r̀:f0��[ON�ҿ�Z�����G�7���Qs�^��A�7E�`���
���~�b^hh��.+?}9�"��'d��|�&��Pb"#��1{>.nk�#�?7��GV�~(�,+z��cm�����dEF�kx.;��ƺ��l���R��ޝ���l�Y,�����\�Eआ:�ۭ�amM�3�����܆���5��~s��T�� ,#�I�}%>F���ܶ�����!r����͵����.ȝMh|d��&u���H?�%ԾC�o%�[ȡ� 3T��z��qi��?�a\F����	�j�$�Ϭ�i�q��o �dz�A/����4������F�_^{�����f������s�TVc��N~���i?��r��K�R]n���W���uW$a���_~�-j��+5u�Y���K C�w��y��}�*���<����-y�� �Ph��������{!ĬՒ�G��xI�6U�8��|�ܶ���PK5%��!i|C��g"�Z|�E�H������;;EŔ��b��8�L��a#�Q<6��0��p5�5j�~L���Ӊ��i'��Z�={؁(�>q��4A���e��7T�gְW�F]��E&�M^�����ŏ���l���H�	ɿr��Z��o��N�����"m�"8��i���pr��.^w���%�{#��4��*����K�u���9�V���"+�������g����Q��K%&+=zށ�����w9N���moJ�6	�N;�GXj�NI�ahx���O �&h�����ts��.]�a��ʟz�&o���ԡ�+'���yr��;8�c��K��q�z��%p:��0:I;(Zg�����N� ��i�&��H��^'�˟E���������+v�9Iȶ��%_)#a D�Ϝ/�^ ���"Y����@"�^�Y�isL[��d�Q���ޝQ:��0^��zcM�$`u�db�ɧW� c��8M`rI�t3	&2�hm.@Uh����@v[��ӕǖ��R�uM��*[��p�Д�$A�ʿ^�>_n��H}�Xs�HNO~O#�on�v�I�W@���Hu�O�����;$��!�Es	Ξ��5+~iѽ�H�B��m�����՜l�WyɢƳ�Q�yI�����6��zHu�D%#�B��3�B�N��!<\��ҷ��l���U�^��[ ��Y��8���L6A�����gu}I��9�Z�;��?�5ΐB�;��1`Ր;�I�{�e�Zc��O�������~��ޥ'��;C�h��������1rxq�/��4r�ٛ_���G�f��@7R�K^=�$"�nH"��C��j=�zf*�L���8��P���v�_�y{z)X��ES=��V��	�	bK���F3|W"ݐ@��)��gU��7A�_]_@��~.�j�`g� �@wT+^_uڊ2 f�o�(��k��p*�m�J�;�v�,~�\:�L���l���8]�c�Uj'����8=��@R���E�:��7lH*�\/,�ؕ*H�kꁏ4��'OS@q¯ѓhǈPu� �[|/��H�=֜�j���;��(?p�/
�6sŃ]�����#,�H�x���(۾ڶ)���s�I���_���r�5]!^��G�f6F���(��^LM7����R�E�ŁK>D�>o�l����܋��2�Oi���/�$�l�c�v�1���K��P�(���Y�z�μ�pa�"�￩����O�T�ƶ�~�OJ���I�K	���_x[B�/ɴ�'���扽TȻ
C~������:{4Υ2k�!ځ�*OȺ��9h5A>�`L�9r�vQj��=#����V���б3����m��Vyֈ^��B8�*�L@�{��xy��E!��{�%H��v�;HS��Ե#�����q���J�� � ��A��?����(�?K���Y2W���5��=(fW!��c8�g�>h
hǯ�Z܂#	J6c��&��U"�t�7c����W*�E���Ok�W6�[:}�Z�x�Жl8=��Ny3��*ak�jn����d���uz>-;K J�]<G���XG�[E�vC/3��ޗ�f���W O?�U�ɐ>��9'�:����0�LX�0@<}�|�(K�>��&Ő�b>H{�R�0��}_kz�5��$�7�u�3U']x �Ɋ "[ׁf�&���2��)�����H�)ۡ)����+P_z����<x-N�̼���r9h���߽!qGN����y����)&i:��M��"&��\��v�
�����)���"�V���x�%��̝�O
�YJYA����'A������.�i�ՋL��ݜ�ͮ�<�",����L�I#��X5F�r��UL��ܩъuł�����W���w��[78B�Yu��@�4��Ub��B��r7�W����<kF$҂�(
�{O�%��6���.6x��a.���g,�&�Qc���YMƚt��T2ε��[ˮxK�:��ٳL����
Q�/:�}�EȜ4��s��#�%��*�9q},#;\��]�Z��<(�t�$z!(r�'H�iګ��1� H�H�Vv�.�{i��i��H��Px��]�dA�h�o����o�@P�	�Y|�W�j:8A���WV)D�){�����6~p�������D��kF�P�&�C�bVt��y;L��h���^"��,%v�/ve:Eӣhf9.u���Z5�7�:b���^��/<�hzF�DP��Q	B'�s'�o����=+F=9�F�b!�P���4��e�q�ș�T�pS�`�*v=��6�H��]T=˖ϋD�6���ވ���T�.౷�f�R�L8�X�q[�=\g��HQ����>�;\�����9�l�;��@�	gJ��������`���'�5��n��B/6I�b,�\0�w�?w�Kf�E���+Dtu;t3E-��9�GY�N�։�T�D!)�*����0z������d�kZU���btw�Ex^P.��{e����>�ea�F9m$5T5"Q�4�ɧ۲��{�/*:��Z���.ޏ�7��NMF���Ы�#�fri��}����g��)�f�r�w�Ӽ��#2��;�%��δDf��~֣׃E��1S��+�c3D��&��{���խ��>��/��c�
<��4v.OHg� f>�m����	T[�����͚Lk����B�RC�c�4ۏ�ihD�-z'��Q%���@����Ù�U���dN	mg/y�����y�/��}����y�2l�2k=��%�6��Ƀ��ɪ?��J[�7B��X=q3��k�ᶿ}$��h�@� q���/ԌE����5%�`��JQ>Ŷ�=�E���نl�N�<�j�C;9?�}}B9�����.�d�}�u:�.%�	(3�z��b��S�oa麒?�|�r����ip�~l�Lpd񌱵![Y�1�E��X�I�l�Ih�
�X<�r���b9��Z�R�%^��Ǔ�'���9��I6�fE�M4;N��p���4��zi��O��Z��$�I��@K7xrR��)�!~*�窡d�u@��4� q;=��2����i8��J����Q�k��uO�&.mb\��2<��Z���ܣ\�nĭs���n�x.޹7D��*��2=y��a;�U�4�(������n���*�J��zx8�V۩�A����F�Ԋ39Y�Y~ ᆌ�G[[+�.�kYr�I��(�85
)̠Y����w���@�C����kv��Y��Y?���0�4��w*�Qr�� �&���
m"�;������c�X�S����as���_�6�mg^�G��;���\ b��jV���n~[����Lk�2��Q������^�z�^�K��W�U0�Pᤧ�K�0!�9����3�(镆��,��1&y���|7�	?�3��J����,�.8y,�?�rG����|I/��a�+_�Q���%ɷ���[�T����":�4��ǁ˛�wo}��ʣ�8�l¶2����1$O�e(�h�.FY"$>W���p޲Ft��V|�}C`���� w�Kr�+{��{��ӠBD{�rQN2]�9�i���E�t!����'���I��$�"�$�x�1�Ɗ����۲�W�������c1�ʐվnK����=��k����+L"��'���t�� � ��v�f�0�Q�M!��� ���X8���҄F�wYB�!:�P^)E���^m��T�Zx���K�i>�7�-d-6v��B�	ͭ��,���D��#����6����H��d��~V��r]L�(W�_
\4.н٩�LL�+�G�M^�?����R�	�T.��$�#��t�^UK���k����6�r���h���Ð4[1��e��\+i3Gl������>z%��&sV4$#�OJ�u$�һ�k[v�N�R�$.��I�?I�ɫ� �-\��㧣�oq���vW2-��q���a� I�Q��Cf���gzal�!V�9<8\����;��kH�I��>PNH���/�˟W�C�*W�"b�b���7�j�f`ٲ.��1 ��ϔ��4	�
=�̬"R[KHk�ꁽ���ЎmzY����]����������b4F&Я��
4��}�.��ONY��Ι��?u����No����u	a�Ksڞv"z�n�<T�b�I����:*�ڳw@o����4�1�A�Ft[�@D�8�c6���$T#17����������T�մ\g�~�>ɶ��Ŭ�t,�� ��k�^��j�X��:Nҫǖ�;�5�Xj��sk�ǁf�T���?|g�������vq��6�?�QoH&���2��0��٫�M�jk�f+�ʂ'�2�l�i���h;F�zf�$��<��VT�V��@z<�j�x=f�2�R�;X�&3�����D.'����w�XoS�g\�U@�Ғƈ�)*I������Z-�7���K�~>{��{ݏ	��#������vB����-&$/�	�x>8�w�+f�=�̝&��زY{ߎ�Q�o��"W�,�Cz�~�n��4�E����J�U!O�	S�7�7��:�e��T��F��`
-t6�Z�'C���b��ߚOj-��m_�U�B��o�B-fK�����!Ԝ�����xI@\�_�vC�3�ƪNb
N��R���д�॰�(��6�Ņ�	D�c
GED��+����ت��B�A*�������1��xp��C��`�e����X� �y�K��
�R	̩ԝ���J=�� It����U�X��x������� ��dE3[�@���=��#(��+��V����􋥅�8HK]�R7��4����2d�M.Ĳ��_�����-cD��>��7RC�l��6�$ ��(F�Z�����*��`���s���0h�e��W�o��O�]�y"ހoz��N'N�+N����qT<Y�i��M�>�+w�[t'�������p(����FL;��u��kƁ�-FR�]��V#�"Eu̲�o����(�5$��SfT�K�YONC����'�c��f�+q�����y�vjG���1/wp�s�%�e���<����P���hA�8<Oq�&�@z��h	��u Q]���PzXɐ��[nWX0��t�����9���$�����>t����<}��9��`W'q�*��Gğ��F�����A��ʳ}<�`u�w�n*�O�jK���y�0�l���9-��������
��X��{X��p����L����O;����4�t����S���e±��M�F�D����g������Xq�t^bM��&d�U��8�����pPZi�����n�ᄻ�����x��K�~����s�9��E9�"��7ƥ���b2΂,�,AV�	(#-�Q���c�����M���'/Ԕ١��d�E����7����c?��yh��Wg��n����m�0Z���ҏ]����rU�� <�8������_$�����k�\h�O`�7z*��놼Yt��^��&AK��������y+�	C��˅'ʞ���DZ�ځ:�{g[���t��F ��W={Hz�#ڞ�S�h��3:o�D�"�Pޭ�)���u�D%�)�1��v�m[ڡ����G�?���
�q=�s졋���mEU?I ��j�I�R�<��c˅�cN�A�x0����/�z�B����	Oy���Q�+�
(������1;s��\x�O���
ۋaF����0�\e�k�䖩'T1�#�m�0[�R�ʊ�� 8�A/�*�J���L�M�(G�?��p�$�����S|g3#���L@��jz=�gx=���\7n@Vjr;$��q�ƒV�8�X� ��WS�`�h�����ԅ}=��r���XK��(:o�� �(R�Ȃ�!U����� I�����'�Z��NmM-�x��Թ���%���,�7�{3Hh��v�njw�2jT,`\rt�^.Lt�t���+�����˰;!���z/��4M��Ho��Vj���8qb}T���ٽ���w��%m�iS,	��//�</��S���Qɩߣz$�,�$.�9-�qr�0��N$�M�a3Pu0������l1ݸ����y���>��e���G�ߧ�ٛ�r�=�jL����ӛ7���DH����t%&9<�Q���4���N�L/�`������$eH��y��6Q�23����"���`Μ�@_�4u�0�7������$W@}[8��\9�q�-�N�H#������G*���]鹖AH+E'@�����}]��&I����#��K�6S=FH�(�T�8⦒H���2�jn<;�rroE-r��!����N=q�H,�u�kV�I��O���.�w���Ș�uu}��rM�ڎ�̷�J:�����/�-�M[]�]�N{5fR�nK%��8�wٞ�Б�W��?�M1��5 @� x�A-0=�t�������ŧp����-=�=1e����6O�y�t����@��������c�d�J:�y�bB�Ar��D�q<��0@�`�`����$�7���<��HT�~�����g�duMfZ�^������l��C�J7BX�
�*��:�7~�����T�}�z�8��;f~6__��`n�h�}�j�h��P>#T���(���>��WP���T�!�1�����A�
-�O{�Ti�&�8��G;}J u�+3R�����M�<���������-�,u(�*ؓ #�ˌ�A� ;%���ojo
�pL��Y:X��\c$�.���I/�����[As�цȷ+��@��j�
����$�Ηe�;�f�ZqI��ۈ�g"l\QP��i?��P��+{=����7Si�q�˞��e��M Z��@�چ(��I6� n�; �N���:�X�b4�9T΃i-���bB=���b���'d��.�'��]���L)xh;1$��F�	��o�x
-��uSV:ٔ�krM��[lHɤ���f �	΍��ǣ�q,�w�c��+)��g*�|-�fWF�o�W����~��q-$���L�u{59��%"��o�od�Ͼ�����	hA��!�y�m��������r���`:Nb_�/v�~A�
m	�y
N�p����M@R9���ݘ��w=�� �2�@�x�"�a3�H$��*!�.��2⤚����Of�b�ĆÝ.��o����1 C�5#1t9�/
�z��wX�'Q��*({�?H��{�ṶF@��ⵯ���X���
�1��>��5ve�� �)7�k�3��Z��+��Lڍ�-r�&"+�¡�.��B,є���.g���;��ʪ���W��r�Ƿ�K��G1���<1K<�,~�5�pO ӳ{�nJ�H*~n�׸�i�4�q,8!Yy%yv6D�9�ufZ����V��=�����1T�o�憄:F�f^}ꚩ6źɕ ��%auϫ}gܸ����X��!��`����A�t���(n!�\{��ت�؄��SصT��y͡.�+;к�j�l�����QᲝ`u#��HY�a�~�Qkܙ�L�����	�TL��q}^``Ý�+&
� �����.��:��
��RbUB4�{E�@����#�9��}\�T�V����Q��<1G"���9�(�����^��rqXO,Ҝ�������m�/PN�.@T��~<B8���I|�7�\5�W0^=bHr��$��.�W�&WD�C���iӾ��Q�Z���pvc��-���_̕7�������pe���]��~%.�,���l�o(��v�4ݰ���Y��cr7��,8�%0���Wq�UM4*U�rF��۸U͟�d3��YH�<�T��S����ou�2�:����Z�
�9%za���_�C<�I%��������Ž��̼P"��6�9 p k�Jx/n���:I��DԵ����G�F�����3͟
�=}���|K44omQ9Ј��<��:�� O)�A8�5v��`n�-���%�L���M���5z��+s��[?/�_$t�˖�@�Y���N���;�	w ��x(���?����>�X_�(-�k!{�׽~�e� =4A?pݧ��`*(��y"
nh�S�w���+���1g3*M��MI��j<�k2�����C_����ʥx�P	c�ߤ����3�$� ��gs ��A������Z�-A�3=�/"WP(���J�p�1���s��0=���.�P�q�܄����B6фq�T�Е��gxF*+X!�%����yW�Jx^�b�o��:P:'�f�rN8�}���}ָ�l� W�M���l/u<9!/
S������ �Ԣ����3'��J'��A��Jw��R���L;�y�s4�W��]�L�+�+�{�DT��t�;��f5R��|�� wI��L���b�����g;����Jz�un�
�27GҾd�|=fdM��C��$���z�����eaQ]����3���(�^!'�h���7Lh��0�=��*ި}_0��lj�1�r0"}�D�M���OS��]54���~�Md+nf:m5��?R����㍫L�%R-*ߏ��ߒw;�8�.)���*O�t@�����7;{�)�'�|Nإ�������h�L3�)x-w� ���X�	��n��nS�����Z�-�t	6,8��P�
X����aU�$!�yW�pCuwy�3RS���9NiC��w�eY^3������߁!�È=�U�`�0K�y�:eT^���z[����o�#��տ�3ss��ѕ�.�㌻T�U��b�iP���Ias��@l�"m@謘F��tE���{2<<�� �?�j&��c�N�u�?f�K��h��y/����~蕓U�'�?ag�/Mǿe�
�*=�?��0�Yt*����x���m0��/�C����_�H��jLGI�=�����7 ��}z._�
EWіw׌s��1W�I�?{
`4��o�<5�9CA�8%9ҽ�l��Z�Z�E��[��*xw!�fĮ#������]��P~
�ۅ��/͙� �c3M��Oϩ�(�O�[?�H1�^B�]`�u�'��Ъ���h�t<yKp�;�i�\2��ά�6fQ��'���v�O�6M�B�Ǔ�W��N���.($���C���9����X��O�YH+�8E�\��R;���@uv���)/L�����s���Y|�ع�"�5s�k��@�Ƌ@&����-�[�,�/���T��niBo�0,�qC��?�\i���a�n�t��\׋���f��s��](,�ħ/u���IM�z�����1����I9Fn���k�x�()��s�E�\���h���r�D�[����/��S�/Z�8H�>��\�{?��p��g�܋�&��b��&�'-=C��dq���rY/��%�g�ȼbc�I�6����v@�&�ky��6<��xs6��tQ�}]K�>��د�nҶy|��I�փD��=.�;Fen��3m�+ S��]Tj�+�3�0��.nMM�0���F8��a4qQ���G�r�����,�g���V��H�~&t~j���aR�a^��/��zihV��?C*3��M)��~��P0xߺ�åY�=.�Ԑ��2��wb[�ޖ3��g�r���D�����K��Q_hXd�l���\^����~����DhW�&&��+Yh�z�����f�����wu7�b#�:�ɜ��T��U��R�LZ��-�;�8y}K�������u3H��m��[䯪�H�FKR��S�����[�tQj��bq�j!�����M����*�\����5�(�Ţ��A%�/<=P�c����F��2a�u�غ/��@��d���T6�f� F�_,0_^"�s��u�H\�Z�P�`����_�&\߯�Q�]��0�����
��M�+W��9Z��{tm��G����I�4.v�̎�{��"w���0��p��i=���qȘ�*���	i�"y�w��[`���!�P�ة\�M�toY��X��[}�q�����2��gWbͫ�:�R/�J{�LAP1�\��`M���8%B&�M���Ѓ�Xvz�P�|:�E� �+)�&B8�T�"#���?�s�_ʙ�*e��Cˉ��E.%���ߩHn�/w;�M]�i�6ϟ��=�q+P��=6� �o��o�;3/$*B!a�h���&�����0�&�Ią��I\M�e��PB������뾢�(��:O	�_����Vh+m��d<8���~H�^Tk�q�� ee�����h���NW�\VՖ쁺�0e�G���P�$PG@4'p�9�dK�&�������?+�I��n����R1Q������>�FiT<��-�#�SB/�0��
D�6e0&RG�0��W�2���-*ѥ�������kq5y����p�����pe��!B��_��d?����Ϗ蘬��5���c���_���f���B,�֮J�?ϝ��7Vy�M�=>&�����?�K(����~1 Q�ST�}xat� �
�N���띻�Ӱ�;�|��mws�Q����Z	? � &��M�GX�����[[�ɉ�H��<~��S36��N�M���A����ޯ�2Ф;A>�b-�QR:,��F�*�c�P�ihM���_$�c��b�lɿ�&������ݢv�����jMK�~瓜�ՠ9�E!��B`y��+u�o���h� _��[���#oӯ�p�mx��ܥ[�e�@���0:''*Zp��D:D=5�ȧGR��S�I).��9�cfjuܩ�	��z�Dj�^��ZiٽMC�5&/�`Y@ih��l�E��M!3��.��ʞ��q��_��_�G����t[�PG:*(Wt�h�O#21�v�#1V,�5߫���2�h�:SZ�?��' ��bp�g*��l@��i�E4���m71{���C`yO�3�@���'�ތ��ꏣ�Έ����yWo�B�ƍ1BK��	��<��QuD��=���K���v���Ƀ���ǈ>�a�7�H���m�ϧ�a��fv�Q�lIR{ӡ��k��⃔��u�&�r��h��2��_������'U���b�����N!Ďm�8mJ:b�T'���5��K2˧��oOiA�7_�{|������������S\"�����v��+��,nP�R��4̥���k�P���q��듴n`�{%���	�IL��qTƊSKl�Զ����n��2��%����]s�����4¹��N�|�����:��{by�#��?�m>��&f��jq�������0Z�Q�9Wk��p-����\�P��f�<�6��'��0t�mT�J�G{��\�6z�6�GI�Ѕ�e�@tM���z�꘯�a�0o���I�;��٫1Bq����A7����X�Y3|_����`������9ϊ��ڡ��Mp2p�����7l�������(!/���E~��e���3�w܃̈́�(Ҩ����N�%�a��x��Y_\DGH���*0wQ����#ﲕ7�����/�S%P�`&�VN۱Qg��Jc�g�)ܺ�,)!;E���\���N\yþڦx6Nf�MIH�����(~j7B9����$j��\��{��[�Uc�y�e�;���cd�����9���CCC�s%k�w:.��f�a3�S^���	�FHR�g��1��T�22���V�n� ����\�S��H}��{m�g�����r)_� �E|��s�]�#N\CJ�(s^��{����R)�^-V�H�>��+��F^�<�Oߐ
�T��
�@�[�;�X���C�  v��0��Y�d��Fz�G_l�6"�y'�tmw=�s-��q/����Ѐ����h+�2����R�"<>�e���t1)֕X�\쑻]sHK~;��L�'+~�=7�8v�} u��4'��[������8���<�B6Y��E9�"�[�����P@oJ��4&]A�l��[1��B��>/I��#���>�!$��#rw�A��:�u����4i��0���l*��R���NwC�yI����g���xg(U��+�'���E=�8T��x� !������;^�����_W*�ԩW4��|y�G݋`�9m"��N܏s�]�TՁ���(|�<y�"�0P(y�xсVH�vX�mt[@��W������Q���<��b�otO��L#���ѣ�����60{�%pR�\�2�&l�>� T��2}�H�4�7�4D��7BXhqF�A���P�NT��ݮ*�R�@�3~�A\�9:�x��)����gf�l�ߎ+���N�V	�������������b.��ݢ� KX����$`�(���j�xp0bI����`��@sm�B���;e![IR�����D	��.��OVl�o
-
�;�lФ$�P�i�6@{C2����@C_8�<�R�[�U��v����Z|^���f�=�n�
�7���ˢ�f-s��� q�C����}%�{V�Ѹ|��MD��������f��������q��kI�-bOp%eZK|�6,�n�|Y��Hgͳ��z`Ǿ�GZ��+H�T�!��'�i�ί�����݀X� fg����]s�t�"�w�^_���"49�&��=[�jy�X�<Ev&�Ư�ί��J��l�S����IF3�^��sm{z5�Z+������n�0m�2]�Lm�ì�,<�e�`�����h/�0N({���4;���m�4~�y�P8,�t��V �Ћ7����$�(�P�H>R���$h�A�b�Ҿ3���%����F�K���F�͓^����G�b�y⑴?-7f�z|`e�
����>"X%�9^r�RCJ����-T�?@&�# ~��=i�h��ǋ�[~�"�!�0�Q��'��o@�Yqi�/VH����־��Ye�/���e��R,�K<�g�S�q|��2H��5���,9�&����O��%@��6�X��T}�f0ѱN�N��l����5��4�Tb�s�_#����G��*��%��3�V$���G�"����E@J�Ȅ	��jk$e}> �^�O�r0��Ɨ`���,[�h�̏��L��(��B
Cj��!�A�ɽ���L(��T���A Ҡ���ͼ�e^#���`w�n2�e��Ks�|`�|�C��;�fi�h$��	�[]�&Vڟ�Ɨ�E���=���X�qA�#t���-|�)�V��i�˯��$�hfF���s'՛�iZ��#X�Z�_Q܌@+1��$xl�fu	�F<ǽ#t$L;xz��Ӟ�ۀԀ]�EЈAz�K���c`v��?fM_�[��ni��ݹ3��ӫ ~cQ
�`-t��ʚ� {2��d��J�DNS;dŎk�D�%^�rآ�Wp������ɽ�Y��4!)�-��T��7�0�OA:��;�;sCĦ��Om.�u�ɮn\��E���qp�kh{��N���j]y.�����rkS��Hgzb^V�Aۼ��n^I2�������BO�g�@�5�R"W�������!���F�n�o�V��7��B�.��u �0,��)k���hǎy;��M��~�����~�>���=�_��� kpĹu�YB�^�3�[�%DW��Ի�+B�Bڶ�k��G��6*Iø��\\KQ]�,����^pG���"=�W�Hwc?m���R�Y��9�:�"�#�Q��f���N�"_�轫I�*�ԧF�3�!����g�e����+Qy����4��h��H�ͷ8�Q�"ew<d��*���a��� ����ϥҝ�{�jELSuR�r
����K�n����y�'O,7O���r�����2v��z%�s�$)ޛ����&{gaL;�#V���>B5c������;@rU���릸Lb>�p��#���X>����Qn�5�r^�-A�NQ�nd��T��8���45U���yC���c�xi���S�ؐ |�}lW&����O~Z�4�NM��>ni���X���x��$za��$0��~�{)�w�}A]��q��o&:@��[.ǫ' ��H |�YNBif"��I
���k3o�Xb\b�kG��6���u%ـ��X��G�C�P�W�"�Ɛ0�f� K�ƭ���>$1��yK�S�8�A7j��veEy�&�AQI�,�0xy�L�\�t'���&H��d�:��}���36%�X��W�.�Y��!e
BV��`��c��f4$핷
�UXl%�<5-�l�a���'��W��b�`�a̀��.`F0(�u���TxL��Aһ�kw0l�`X���8�T9��75 �"�FXFk�9�]���ɇ��b"�w2���g��#H�Z��U	3o�S���ߨ[�jN�kVaeYmW�Jn���х�7+|�9������ݺ�]G�>{�u �/��%P�J9y�t�(�������j����c�N5)S+u|c*.����s$<aUpG��^���Ȓ��s��p�@3Rd��Cl�9����\�^������=��5�rs��%�9��v- ��V�PD��A�vY˝f�@n�(x4�B�oޱ�*(<n��y�=�2�l� kw;�kuΐ'�� ��X���(�c���y����^U��J|�)p��W_R�#��3g,��p� ��W�(�Ikv���W�Z�{��3!�mN�9��+���E`��sq�kFӣ�\�>��*7T�:�\T���?�Cyٷ��#�Y6ӟ�=�ΨHc9�`?�&�gA"X��q�b*�h!�^�җ������ )�E.�OT��Y�� �E��:c�m5�$�_����:�l�F驂H嵻� W$_�0�p�7et��Q`��3�9d��6?��?	tl�����/OH�#���O]�d)�kW���UG{R�O�|�a����n/��>��+<�u�-/���L����1�SE
e���޵��=g�Op:.=q&	����p5󙜶.W�m�
��y`�Nf�ǳE|�FQK���T��*נ��v V�@N��~�Db`m~Y���s��4�{*D�pL����I!Z�}��p֏�U<4�()��TDF����� 8�=u���5����K�'D(�S?Q��#�����meU�'���7����Jn����]�����}.W�`hW���sx�X����L�˴�D��|mĦ��'(�"4w��f�;���6�����sp$�c�6��p��	y�o��br�M�H�٣�q	Q�]8�#�g�C��q��ʵ]$�O�:��jflʈcCG�H=�����a��^������;i���/�'.v�:M� ��rzq��r�Ƒїq�*��Ąӹ�������'�Ԓ�,�"�Gb�zZ��9�gE}Ņ�d\������ف�àH�&�;�b�TM�Ŀ�<2b���H�C$��բ�UN�����b��
��, t�%<�e-r��Fp��
�;�1~r��2E� iE]?[jN��PA��D��h�S��PN������L9�B�#D�)3~��$
��,�0���ݨp:��.��R��'5r�k���S8�t��2���k!�^�PǛ%�bI�`|	h Ɛ$l�ۚ�:'My�K/(��P�Т~��n>�P��3~ъ�h wU.uL[%nE7�l504[�O�@)&l%���P4���B��(E�&AH�LepfL9��mxED:�&�}���	�I�2��9 %x�1������,��, V��BӃ�6�<,�8��~\��e6���Cɟ��]�(Ijft�1�P�m��+��k��k������QР_ۯc�B
�lN�|'<�>���ȟ��/�f�&kB��(߇Ն�K�Lh�$����U�=���s	�S�p۶%��jG#n�f��)���AW��X}N��F�Ӕ��S�ޮx-�lP��|]xq�A�[�\
�[����F�����\L�=���c�TIk�s�6���v�u��8�J��*7BĔ�� *�ܝ4�o�j��?���f�Yn�����A0��y�[�����/�~R����\���LA/�_��gW��f_q2�����l�K�"�}���a>k֗���,>4�E�A-���j��#m�qή�Ǽ��Cb�}����;OM��,�mI^��钶�%��?����s7�Q��z�N�e2��q�-�h�y@��,�']�G�f��>iu�G�h��p�<&�4]�����p�f�O�]Qиƻ�V���;�_���U2�j;���)a3&E�-3�fש��.?ܺ�f����yg(�U��^��-�0DѮ��u��j���Y���r�JD�=��Pn.���a+-e��In����)l����b)����j�L�BA�uM�UO����C�[��y��q_R��Z�.������l&U?�[xˮU:�k��2j�I�.?�N�i�J��w{���CP��]=?ܴ2�����Z�ਜ਼���Z8y}�*�0�dҠEꂹ�� ��Wk0I��ۊ+����,���*�G�bj�BB9�b�=��N��od�S�M�\�i������O,���Wk�L�l�9�Dn�=,�6�dN^l6̊Mm����*�ϳ�5��!Yj�;�5���iǇ��4��\U��ϧk��Xh Y1��z�_Hb�g�-�!oS
�JYU3J�±��n��?�Ĺ��'�	���I�<��ٮ/�dO��1�l���v���Y>�i�ʚtW��6\E���u�H��zy7݊�"@��f�	���bi�&�"�,��މ��X]���&���۶��l9i�ڮ����K�-F�o[���Җj�J�����<}��~U*���;��:�^f���	)�f����~ls�1��E~/--��ye��,��	�p	(�(K Y��lO�Ei�����
��H�QԦ�3c������O:�z?��	";b`
d:-�Gw��lg7��Y7�P�@pZ[�S��Ǥ�=�'Kp��X�uy��{zz=��H��7�������+ϸ��I��\�R��J�+��ז����=�.��<������8�&�����NG݀�J�ڝ7��� �3��R����-�2��)�N���NH���#��cN���l b��-uj4+�t�GNz�l��O�,`sE����P��+Wt2�2��8"_�T��O�~g���*��'��K�<�AY�{[w��?�l7���:����ǴT��%%��v�uRfE�ǃT�=at�;Ki�Y�3p�],��]X��:i�]켕����~m� +�Y�E�S����vl_�{ya�ݶ�ßyD.C��9�虷ւ���w�:��v8}��F^��Zx֭�6��@�B����'k�~���͑r��E�իCѝ�86J0�a���A��:�d'��ߪQ�<�C;d+�x��:��˯sը� ۚ��xY�&�~(�
�@�Y�COw��mڣ���z�i����W����Uo��>B�)�����4RI9�y��e6�
<��s���'��0z(ͽ�t͸�՞�)E�d��@�,�=f��!�T2����h��
�O�{DH�Ƅ<[g�6`9�@���F�Z�&jaR"�J9�#h"��j� ��Q`<˥?]���7�C��$$���B��-Ud���XP����$�,��Sxǰ ��B0��M.�e_+p��CD���،J�?�����V��hje��1x��ܴ ��l[]5-���n�G��l�ݖ=W[�|$�2�  �}c�4~bo|�0'�m��m�9�_ʳG��,�l���c�~�=���pg�Ҥ�L�?�A��U�:=�����T��P]������=}�T�3h1q(O�X�}�6��.|�:9��՜���fh5P��M���e��H�����G����Sr���>4�Xȥn���7^4E���]��G.� V���������[Q�
�3��O�^�\��2d��^��,P-BW�S��u�;�v=�^[�cye��3Ńԥ�r���W�������c��a��8H.t��(��]CH:���4B)��DdOk ��=��Vy�^"�Q	����"ȕ-�Lsn�<��fF��k�#	I@p��:j(�ӏ��B1�B�p Z��� �d0h�E��Ϣ���m;놡��6ѱSܢ�>�Z^�9z͓��
�nw�o��+O�>�|3�6?�K���sl��ȸGR��	��2~�У��+��b;�u>�|�l��5z�������O�ŀY�]�+L]>ң���Zܧ��]��n�{gປ %a�ɼ#�DB�6!	ʫ_�3]`���e���wf��>m��{�S4�z������s`WhNvQ�\/�v�5.�FV�
�������W��~zL��dC��䓱}�"X�`Y|��j�߁@f�I��T�o�bg�D�w��NmG�̾S��|��{?o���z�Q�i��%?����!(+x��:����f�.�S/܊û(�h�|�o����s/���
-�����r hHN?1�NhdE"3���YOl!����L��F�p˛a>��q�d��p��$���rI��5OiiD@�dy����.���8X~W'_3�|�Jހ��Jl�lxM) H!K̏�T�W��0äj��Vo���l;�x( _ra�I�p�a������	��]f!yL�2Wf����A�V�P������|=� ���l�嘂�4�7�	 �	�;�Wr�I����(�u9W`���]�C�����}�9!y�m;o����>� C �>_������啦�j�>\?���GܞɻO�%}��/V����xc�=���E�Q��#�v����'�`����]�����c�d�0�W^��+��d�ec��Z�^Fb��,�(�[g�yG�4���.�ڲ,�J7x���A����!��8���ٌІ���s�%6P��T�
���u7����b�8/$��;.�dU@���KhdH%�h��d������!o��%h�b�AvXԌi#��8��p&c�	[
�W����M�G	H�s{d����X�PA�ѵ	���b�[�R䭯)���`,t�3�9I�V	���.������w�1"H?����^�Q��ȍ�v��>�Ov&��qPds�v��(Z�`���٬�g�ί�tv���g٠��%��F��{�_\�zix,�v�͢^�<���A�n�Ӣ_��9���o�����iż�V�Ox^�"��;�4�> ������$Ϝ�o��'�s�K�xӲ����F|�/�N�1N�B|-1���(F������_R�2u��H���A��sZ�`���o���L�ޖ3���`c��<���u�;�g%繸�0>%�ј29A��u�e��S<�9���PSy��^�
誜�üc��)��V����xֺ�,e���ga��Ly��-�O��3��f�=%C��Z2]��٭��:]��`F)\��r��ڿퟬ�r��Zנ�4�1��N��a`��=�h��x�+va���P����唾{�ؒ��[O�#���ͫ�[���H:[��1?"�s����<�3�+���vF��+�P��CG>�xٙ�=��mU�&��	�,�q�t��#}�ubbi���P�/�R�+5Y��ܻ���Y=*��+�k��	�����A����c�f����`��	8������l6J�Ӿ*���46�qy�.�� �h���.�4��Y��S>yίj0:S?c�:�۱𸞚'�N�1�׮���Ll��]�~�W�BЩ^�/�Q�T�/.;�_��j�rl�� J�e����Ⴜ!�����-�q�TO|�>������2y>p���53�u��%�yB�*�YE�c��-2�� sL�îI��$�g��@�;f0��ȹⵜY�ހ��i��\erF#�XM�wu������|'0�Ӗb��L�d%r��1Cu�;��\ӄE�F �O��n�k�#$w�d�}¬:!_a�	��j��&s�J�[l�R�A��ږ�dֶb	����nhhk����Bkm�}S���ÐI�����E�\\�wBs6�,ȏ�8>��꙼�b��e����q��������<�<��3Ӯǃ�H6=PB��O����c�	S�,�Bʱx�T_k+�;�Jx�`=fi�EE*�<_�Rfڰ���q	��ը���mbߋ+\h�	5�����ׇ��A��w��V���[y��74�����ï{�@`�$����X�A/�$����T���n�Z`�ЇY%���3��!�@�0n��J��J�~���p�H�����N���s�Μ��5Zm| ���H\��\ ���Oq�`ٶ=D���$��N0�Q�ɪU��mt�ֲ��Õ��_�^��N�v�F��NaT]ĉ� �~��io!��x)��+2�=�4a�F��R��]��L�2�ٻ���g�q��r��pv���ص�C�7��7J��+��������k�k!�p���3w�� �LR��w�,g�Qqt�|��Q��k�0��Tb@�Ȭ�+\���^���h�f4�rQ 3zoX��t��k����n Ka*CW{�n��>�������a�#�:/�ENi���������
-̍IOU�����nIFf~5�P� ��-���$��;�5ω�.R}��l�>(�C����h����F�kg�l�����UY�%B�~P�b�m�3��k�}��w"���4ޡ��_�ڃk5�w���	R"�J^IGk������ǯ�a}tU������É�D�|�O=�Иx8:q�����;r� ��c�r���ڢm[;Ri��ٯ�M����2��*�uɅ�+cz�3��)We��s����m��b
*��CO��n���_���en��=�H���v�Ǯ��
~,6A3'y#� ��G �n���H�NB�ɣ���g�0���%A�:���)�+,$�����e��A�#_au�1Ph��f�������B�q��	Ōo�I2��ڷ�_��+U.Y0j��'�����/���2��L�Q^�z�6�?. ��Y��K��
��R���0����?>O�r�7ŋ�w�O��D؍%��6ǂ�n������/�8�K�[��,��H܈�����#6�K �_������
l;�:��z�3�����G;w�3��`�����)\��ES�ȡcwJ�b~M=:3�qR�FU��q�;�/���	�b�?����I��[�G��+�dlYP|�C$C�9E���)=r	��:$�\���ذ���cZ��ɔ���>����[�Ox*1v0�!�J_Lm�iC�[���U[�l�=�w��߇�Q���H�m��
w�5��hו���	A�P#����L�M��w┿�څ���xwꇖH�R;��T�߀�hyg�E�3"�,t���pS�lYOD&�ޝc\U��-��B��Q~�9��@���!��|�_��]$E��Cs��<�U�4�Fn=b"���Xճ�M�Ma[�BRi�M��7�W��D��
Q�Sd�����|İ;��uY�y:�Sp��HL�b�˟	����c�B����-���(O{d�6B@3jғ^O�N �TV���8y�Y��Qf��/z��!ڭ3a��4 �*Q˩�60�_vfu�Ύ�n/"@;�%qI�U<\=掉Xr��>SQ�����{G����K� nQ��߳�%��:���vV�V��e���M)�AGX`��J
B�}&�����B�ʫ��-K�d4�Y�����y�Y�� ��#���K����H�0��u�_q.�q�笆F���{K�"��r̺9���WdI��z�(��)�u�xy��{���f��^5��XUp�`gx�[��~�U+R1ky/.Frd��^y�&��)�hk�N��:���W�=cL�`g�>Q�k�F���E�b�eUz�֊�y-�����N5��%ʨ{b�a!�P��#ގ�cz����W���%¤�sm-I��<z�-�n��B�~<��kd�)JI��V��{Y���3K� �'�`�2�Um|���PE���1!:������/�l��EM���
��E�U0$k����v4Q,X���}3qf��{�=�`Q^v��5Q
�#��`4Y=EAJ'x��yRK�&b*��'ѕ��N�/�W���z7�ZҮ.�$�B<7���k�S�62���1����o�u�l�؅�םU�k�֐��E�X튜����U�-�`�u\W/܈��55x�P�$�A��K8����ٍ�o|��E�b��{�)��� ml>G�k��b;t�%e]�ⴑ՗�����-oq��E�X$~h�C�2�h�\��8��E���Ĥ����[��V:J�c�Z��J��zW���6���տ���![I�Y�|1�l��h�� M�M��fs�r�#[�:���B��s����V��ptd+�ƮY�F�"K. �A�xє�];�%R6b�w���ʫ?s�(~��;����ׄ23Ta�n���8$9Y.��V�%w�rF��W�z�g�&��u��^��$eGvC�hZ$�7��8E��T
���V|I��q���M��h�c�^�	-&c%�\�$�@���+��k��b.ᡸ�|b���}�P�U2���Қ�~e������3p����M��}�9t.�>�)
���v��
�j�
_J����ڧ1�v�qt���/�H���`��0�3az��[��	NN�L�( �D
�.#g�B��4<u����EO4��.<�Vy�ĭ6|Q�ODH�p,V�+6�l�l���{�{��+N��
�y�&f�nj�V��ݰ���y�����~T�[���L|�֖�����g+�����|�|]y�K���zV�Nr����)g�J�J�5)�z\"��i��Q�8��?������9̻(�Ox�)���ۥ��{	���n!�c9��a4�"��р���h ��U�*`���g�Oh���6�D�/a��W=��r0�8t�� S�x��>JZyY-�_�z���e����|��R�'�'ᰔq�lV��z�rjf�Ȁ�{�ڀe��z��5_Q]��Us�i}mmS��D?I�,��0I+�I�%E��������tc<�����Wj����~~0Y"��Ԉ��|U�rgiyY���L��e�4���r�	�5s&�p!�PSۿ�ǲ즽ڡg&���w�<Fa�M��mEW�s
���T��H�s4��q;��I����aFg�v��r���P�q�T�_lC���/��췋H��<?h���6m��㼈�k{�ql��M�4<��߬d�����R\�e0K(2~+�1���Y� �h��� p
���Q�rq�_g�:��Rmo�d͠�v{���"��D=�d;u��qJ��o$�ө9��6f��٦1~,�w�?MgG�8��NqB�u���.c�Q�%�t���|�qq��L���JCU�#��m�����2��h�Q�%fU�����#��7��i�lEs��Y;� L5;#�;m2�ˇ�/���~u�H
k�nSz��o���z�zP3"�Yy�<�3P�!E��&��#]���;YĪ���;'m��0*���D�{�I=9F�X̩M�K�E���L�6�
@��0r+?e��R��	7d?�D�.EAf0C�19�l�������MΉ��PUi���Dگ	����f��tm�d7��^BU�&?��ِk�{dGd��E	�VYU��K���@|�Bx���E �����v���l��~7�i�Z\�ze4�#�$��5N%-����H?.R��Y�9&:l�Й��8����Dl��Lt��a,PU,�.� ]����M�7:�i��l�C����h�]Q��89�-!�����d��>�[U��,��R�����Z&N���N�	_�X���z֨8���(�����K��mï�/���EXg||X��t�Zv\�!w��r�;�.e8RF|4����e%���X0j�	7����	�^���d"iA0S��a� ��a&�����Ӱ����1�����}6���D��{2tP�|��j�{N������0x>�a�'u|�\�������ۃ�>�S;���#�>��#�6&������Lo���{g���5�c�UAN�tv�b������u�7��i�w��"�[[��/?�ʞ�/Hx~W�ę�w$w-R�q�)f�Ψ���5MN�a��j�/K:�#!7�M��܏�c��	z�0.��|�F�	�;f�N33���>W�AQ��΁X���37�����M�4sW�:j��׸�MVl�^XvB��rU�y
�,,�{�{v��T�#�y�$S�sE#�>��hw���9/@�8	��bCx�@ՖCu7��~�>�+~|y�(T=~�:�Ü�N:�V���)r�Y�]|�L���V�S͋:O4w���^.h�>�wo��ڑꊬ\�d�۱��M�����9�c~[��j|]
��aH��>S�~��y���@���+��(r�K�2(�f���N$�!V��u]�Mᬅ�cj�X�ijo�p��U�Z�g1`�%kTdo�"��R"��3�p|Xm~"��z�Mp��X,�G�5�����b�s��^g�Ԗ������U� x��Es� '�b�F��Y���~x�t��ֈ��%�2JA�^��<��n��%���}�r����׼r�J�i��Ǵ�����)dM��艶J������BS�=}l�\s.ƺ����T6���_���~.�^ݸ@7T&�~]�1�^6,�R}�B�wm
�s^	gH�
�ջ��_��iղ���AJ�`7�{`"<6���ڠ2BKIj9�Q�lx��P�G��s�0�/q���f!X� �#����Z����}6+�!,�R�`�ՋG�zʃ��i<t�����<�W�l3.`�u;�5a����Cg�C����?��[%3�}mZ*�����[O1�ݟ����\"�J*�88�k��t��:�+\	<!ba���w��袹BSk��±��I�뵢��X��o"�)�,xv�����n&I��#p�/�|9/�">��}&�)q%���^�N�o��Sh�!���%7��ӫ¡P�9W��4k��A�8}3��(ժ�]9��E��`/��-�"Y�\G��*��3�����%����Jb�A�Md�è�%Z.�M�$	������O�8�R�����5\7���qp(��YT��7��l5��N��)x�#­ԧ���V=b��{�ti9X��\���}��@�8@>W�X����|�~���+jEH�	���FU��:ې땓϶9q��s�9��~vi��"[.�Lz�KQSC�?H#������a{���as�N�"N1 Ǽ�5X�0	�Ȧ:�C0?��MX�ťd�-�`"��NAڃ
��V��<(�@��\[I�C����μ���%a�E�� �cB�)Z!R��lG	���wcdhP4pN��N*��0fIq1}f���o�♧��z=�O�W!�<����6�%ϖSw,bK�>�-�!=��D��w������� ������{⽄���DL������Y�Zv��=h�,���4�Z;�&6* �\;F�X=��B��%�e�)e����3�ۃ�bO-�y��LuW��g�#��L�H�]8�C-݅8�!ˤ�_2(�V+�XJ�T�
�
t�ͬJ�C�jgN�+�\r?���+
���� R�˱ӷ��ȬK�aMI�h6���
�3���*2��H���S�1W�2��U��יL~S�<�(x	!�K�M�.�;(kp����]���<�l��[�F_�1�PH�ʬ�>x��`
1ȭo�e�R9".���do#��n�&�s�"����&CB0�B
N��<�Y�W�)ʕ8
��������o�tр&���_�,��j��jp�x���W�t�Ƈ�$q@j37Ż�/˟����iR�B�5�{
qk�2g.���U��G���;7�5<����g�/'��p�k&�ħpQxӆv����ܼ#���b�6���\��[3�:��r�@�#��kg�e��l�]Ø�����~<�2����6��zU�'Ըe����������,�e��S�1�9N�Ɋn��9���&\�� gV��K\���jn����J�M�z�NS7^��-�)/x%;%,$�,�s�1���M�TG�����.�zY���*�@��l'��P����O�v��$�9{h�+I�u�-txFg��B�(�8�O��*W����vդ���G���R��W����7��[�Q��#��4ێ5��V��2�����R�R����/I$��ro��VDO���0����+kֈ��f3"~R�N6�p�f��;������P�rs���y��|]��?�O�oD����|�4!��q����d�3O���+�Y�Gi�w��Y�_�fu��8�g9�@d�s��Sm��Z���O�e�
,�q�^-O���sl�"#��*��dmV~��,�\ç����P�~����0.��<�Z�����]���.�C5�8n�R���F��Mg6,-�y8HY�`���;!Ȇy��aɋ-�hYD�q��y~�ʓRV��z�_*�(���??��C��*|b�`��2�Wr��iuG���a��#d購��]p����g$�"�&������YgsTO8>a��N��J�3=
9�����bL'�T��!�ǠB��<�L-o�H�\�M���"<�	G?C!�D�nx7PV��[�\�9 �u#��а�=�ef�9{��"XLT�P��:Q�����d���OYg�M�����9w��5�x\�;���$y��
��Q6��b�N��ۈ滪KIpa貋ŗ�-V�B�..��HbaMI]���yݐ]��Aۖҫ��|�J�L��zv�e e@�� n�S>��l3�I�<g��3s���dL�l�$��\���ryL�g�Ʃ/�!%�m�^k�)��܎�?�x�iهW��M�~@�-
��BG�*���M.�U���x��~�0��D�J��`AO�Ϯ{o7f���l��@`56�G�kD^�f��*�f����>F�|�Ӿ��Ō)LHc/w{��CGqV����+�q���KN�Qz�Z����_�t!�DE��4>�(byA �/;�'U��P� p]��)>��fO�߿�{Ύ4�[�<����0\�����K�Cݾ��y`d�n��,i�j��p��y
��n@�=���:�����A���v�����t{1e2��Rs�Y\��cҝ�O�y9��t*�����*F�|�8�9)�~Чl�1����2��W*����
��#�m�`��ƞ�z28ܠ�<-_�Y�9x�e���<�˓�v$k��ۅZ��_���yaa{S�Z(���@���$q���I��_/�G��Tu9'�T4�k�3�fM�ՑA๳X�F
'-�Q�o_a����ht���}�A�Q;؎*U����w�n���Ԇa�����	���Ɩw��1e�a
BX �/$�:]�W�m�I|���:'�R����qC��x�Y�%��K"�u鯢Μ ����N�y��� �4�ʸ�~'�?��l}8�r�ّ)��d���W-��	i�9^��� ƺ���t�JQ���)Hbd�.Z�" �Tf�z�O8���]���*�Q�VIe�z���&3��fֿ��%_()<��� ~��~���<c�?�rS���q��Ɏ�f8�NbN=-�i,(�ӎ�h2��*������V����k�e������ГS�9� ��BY�C��C�娪vn��&����8�a���ao�ol��X�y����D�d6,�a�R2���3o�S¥$`*@�?K!�i�%	,+isl($��e@FXG�O�+���u�~��YF�O�I>fsS�:���[a��]�����k�`2"�d��}7S��P����j悋���Z�G&WC���m�����lk�hF���N%7�!d<3H������{�%&�e�3�MgV"�^4?	��K*�������XP=�H��˂��M���(xIb9�Z쨺�(���8K=���Z��i�h��ha��E\(�&�)�3TR͖����p*&%����ad:�9W��u4�� ��j���?�]�-����m4��;�@��+H�_by���)�{�Z��.��5ܲ�fa�7�,�c�Sd�|S �<y�B6��c�����A�%n����Y�4
�x��H��^pZN�����h��H=� C��1J�Ϭ?e��Zz��_�';+�;j� u4��U���ȕr"	Y98
��4���."FC��/�G����/��r���4�i(�=�N筘Y^�kQ�R�ȡJ�㬰Է�(P��3}8��g��5!�����"�^�tu��0�5�ˡ�M������z�;0��X%T��4�4��&5|`�\'Y�Z#36�����p]���]��։$�4+�b���^>�v�o��Y���g��
>�͸B������O��!�t����5��Z���u3F���������v����c�.�L_���='�'*r9�1CC�zʣ�7���i3�ـ��#L�m�_��݈Ы��-�.oq/�\�2��(�p���L��uL�2���(��'wB�'N:5�vq!_����f�=��ɶ���;\s��!W;�>#�8�`K�ǖ S&�ϑ�?����scW7���/o��#�ց͎nF:@�&�!5y'G
��U�~�pF�#�� �rY	4���<�uW4��FFr�G��_$�y!M����bց|S�r�5�kA��@�Dʎ�cX�B�
�Z�Y�!j�hzL�+�75�'.$lۿ1&�c�GN�/f����2��_iTMŔ��xɪg)o4�
;�l��)��qDl�o�����mc�FV[�$<A@XpU��:3h<����e��l�C}mpcF�'�D1LV���/���p�5e�:)!����R��:R��Z�J�X81ѮWZ@����U	��	�s��9�i3�eZ���G����!��%�g�׍	~s�h���^��꿠�C	"��K%�q;2�C�`�``�%VmspP����u ��`˰�|�`k��Z�U3r��bj�~��Gi": ��$��t���}���x������G�1�f�t�E�Z��Mb�5��d?��rn &*�� �6@,;�cN����:~@|���Z�;?MJ�,ۋC:�Oh��	���!�������		�d�����Ok���E�R�9����@�Ӳę��e��Ϊ��hl������,����UH�F$E�0�,N6�ePG����w�x;��}�`���C�&�ՄȔh���9g��`�j� Șߚ�w�&i
��Nuc��T�񧋿1m�8��l#,���~'�re�Ey�c?�e-0_�|Hݸ��d���r�ş
*=���~��q�Jikg+�!C�k�%��3� �Svא^���B��K�.--���}����,�zJ	��2��L�~�B�\a�$�@JJr��v�$d�����^��*��-�0�P�_e ��FQ����qɤ�ԏ_{0�"�ۚ�i�����/@7��}ð{��BEj����W$ K\m(?Sz�q�Xy��;���/T��} �Sh^��0O2�����슫!<���>����jl��#��jVڬ��������p�y̙*�@ '7o [#-�*��v�%�_G���N��n�|��J7i2ؓ���=fAKx� C&��/����U4��Op���}�Հr�6�,����]3\�_E�ٲ�ڇ%�l�k�C����;ڮ�B�뿢&n�t�}A�,u�,��7�Y�w��>�����1B�{�����������X��`Ǣ[u�!��jr�]�,j����?���N�L�Q����`t��*�"��=�<�-�]�v������/_r�`z[�znKj�M��^e]��qWG�=+"�'�y����>1ԧ��k�#p�e�<_��u1��cX~uId�]J�1���nY�$HT̫�U�E�e'����� Ȫ��%�$�m@ا;�4a8�-���(SS��I�SY�N0mq-��2���������
�َ���j@��)�<^{`����PG.������Q �~T�p:,�U�g�l���j����\ml����uPR�J�`ҙc^�~���6+���-e5Ȉ�H�z"�,��f�VhN�jT�sG� �8ݤQ�-��a�X�x6���XOrv��ڥ����������U��+ ���L��a�6�����0W�M�Ἁ�I[�T��r=��	[�14g�͐���B����	���&�\�n�VWn؃�M҃XhJQJ�;j��߳�=a E��I��s��?���'A�o��,�N/��)�S@zjW�͏�2`]�גLjvd�u�AH���N@Ko� ��I����Z��Ƙ���9�5X+f�Ч���h�#�m|��;?���z���Վr���d!�s%�+�b_rP��?��7����Jr�(~�}������K�lN1#��b��;~��q䗲	b��:��(3�q��YR<�j��gQf�����w�qU|!],a1�h�{�wW8x��E�0�_��PԏK��&/&n��l���N�{�=O��U��I�i�����칍��ln���i�^��s����˞�p��-_ܪd`}"j��O���v�}��r"6�8�÷n�X	z������K� ��q��i�d����Ӗ�^eFUhi���\	�b aY
��r��&N&~P�GP�N"��@4܈���`�'E/��b~��ŀ��g%���m)��Ͱp���_.w���u
C��3
�"	���[����2�o4)��A3��_)N�k$�%vpj��T�bW��X������g������=뷍�wn�ﭯ�{VpN�LN/1����SV烫z|f�Z��B�G��s|`٪k������O����?zM+WV�(]Ek!킭o6� !�ִ��ZVi�[�$�9��~^�ȋ;��{��8 a�ɐ>T���lT��e�T^������p��2��9k�d}�`	���K��,��x��8��������i�:�PԚL�T�~Z�.!�zfIp��~|-��q���;���q�&/�d2��&�#��ư �H~��w�z1?)����0�cǕ'���$)������` /���ZO�5�Y�\ǁ4������C�[;�[G��/(�_�3	}j�3�@��u����fNp��GZ#�|fTk��ל�>�rv'׃9�X����m�/J��}P�3r���5}o=jِ��h�=�í�B8�_�\J��8ŠK�D��j���W�@�^y����Fd�۝R������J��$��;�Q~����x&��X��|��n��cG�&p3lץ�_d�����j}{�w��
��Cr����?a[���Pr��L%;/���hu���?NU}�>���lą�t.8RB�/�/���P=����B�9.�2Z�J],DR��ѯx�� �����~_IO}ά��̓8Ao|��e睢�p�Ki0�a^�}Y@ �z��歚�!}%�P�����f����E��7q$�G2Q򱏡�nQ��Z��h��1'NpNy���<�`h_�_�T���5ݖF�>�?)����8
�3��L��*0k?e%x�߆l���_Ѷ��@0K�~�	���&G�ɓ�zҬ�ܨ;��Q8�5~��5p,U,�q�&�/����C]˫�n�Q�YT]�XѵWM@Z?�v�otfIw0F�|}�%�u�Nqp��������]{��l#o9���Y1�ʱ�n�����6U�����Y��S�:U��I��&|�l/��2�E0t�=�n�u?�>���od���>>�C�Z�������N2�;:(�HYlc�z\�2jU�T��%sQSL���e���/@EMY���!�'G�l��;�6�*��(�4���_ٙ{�ڳT���'�Gר1��D9Y�Q��,�څb++׆2�>��9[M�3�&N�l��M��@-�� ���)b_�Sx(�#3CR�H��4=�| �ū�Ա���F���T�N��$n,�g�Mq������k�0�mYIR�����	P��N��΂iR�,XR��[EjyT��T+��N�u�1�Ibuq��T�Y\���΂��îRU���B�+��{�)%SV�K$ċv��I]��i�ͻ�ar$#�`�#޸2;mE%ځ���C�Ҙ�� ��t[?ˋ�	\�\�k�ࡋX�ZIp�����u�	޵�r[
C6�J+��N���9kI�m�V��*+(>6#90��.k���� v+��6��^r�>a:<ސ��E�GR��.z}� _�~	�L���ky��?�9�=�4��"�XT�5��1E��΂�E^���̏���>!j��7�#��Q3#�N񲺄�rs͖�e%'^�K��Y��V����$�z��s���0JӋ�["�|.���`�΃�J�&�`'���£ɻ�x��o���_ְ;;Q���c��,��a�_������lZC(~K�6��6�h�9;ڍ��3�+aH2�m�s5!\ ����_�t�%f����<K��tʫƇ{����L�6�n�d����UP��&����X�L@�w�}yb�/v3C=�1�9#�,��u*��+>|�.cD(
�~�Q�!�p��>Q'S����H{p�toHk+ E`��/	�mַ�Dl�eF�Rd�f��.k���з1s�#-v����x0���z$�;
@�䟎��`V�9S�K����.�'�ql����w!�"�+R\p��?���l��1�#�V?�=��F���8���_[m�����mn^ք+U����P��}������R��dĘ�L�$��,xx[v=�Q��L;E5��riHe�����"2wz'����!s�N��t�ɽK�meE����Q�u|u�p�G�@�TW�2��ju۲|���^�h�E���� 
(H�M���������c���Xƍ�GQ=��V�
�~�W��zz[@zvV��L�܎D0�hx���2��7छEa<`Y����#�]��wؾN��9	�H�Z	u%��k	W�h�8X8Y)�A�R)yv0��a��~ٓx�+T�����M����>L�뜤��|�p� KH��c�f$n�H/�!���/�/�n�2>ڸpG��/Ꜳ-p*F�y�{�ClI��-��� �x��\�rS�F���.������?���W�<g�g�TA�?xI��)Xq��6FKdѫ�i���];��p?���NR�ӖTd!"LY���(�[��j��� �r���,F)s�}�)��b�i�	������ 6�n_tk��{?v��{�����~�+�#26E�Hy��H��gO({�ٲ�#�[
�����&�u�Y�k�t��І�U^^����1���l(�A;sa�<r�]�j��(�}��/�6<�k�Y�{sm^66<ԝ�XC���>����Y���� VP�	��oO����)W�YIjU����{5���� ���
&��:o�v]4���pd1��.�{`��n^��~I��/�ZX,��ȿ:2 E+5���K��n鎅�L1���D�g{͢�3E�`H�Bvi���d�qj:�k�萈�s�l1��	��o����f^��r��.�Ղ�Y�Aشr�jh����RJ�Q��$���[��ɘ����>sҿxN����3Q~�2gt���E��	�'��j�L�懬��t�UO�KM���f7���%��|�~���K��x^��D��z,�m|�=$v��	|Â��1�q��_�k��JF��?��YW|��txp�2~�%Ы�J�y����O����=�̯V%��DU��}��dG��@����s�$�)��tJ`�R�C�����)z�Ʃ�����,:�� ��,L�h��
iי�UB�<���A ��aK�X�r��	��ď��iU,��}�H8-S�짏�䯉ٚڄ��Cd9�fJ%�����e�*4Z�*�����81y�)tb�:����7Ah_V��+��iIZt+/u^���?�Q�k0#ssZ�)(��U����H�j���ı�.B#u��,�M���_��_�_vO�ů���{����C�q�j��>,��,�
�v�(���!��^�B)hV�u�!��i�
IQp�}��eT�T-��x��-1|a>�?�D�4r���b���4-�)䓜����nF�����9�������I�*r�c�(��diD��3
��9���ѽ��3Rl&Z�jz��Ƒx�*i�_�5,6��ʽ\��1��=�-XـH��t�A�xw��\RM�0���)g�'VG��^�uȩ�:g֐9������엺�#�A�'P�J�e��K9��f��z
ݘ��Q딏j�(S��u��b:̾�ik��&ö�S�[�e2�>��ӗ�t��]�^���i}L|J)
	2UT����7��p�^��K��m�4]P~&�8
������I�Xeoݝ��/�,��*d�A0��_Hm	�Nk�!b�]�|�.���;����L[��Bz��Ry��I���a�Awv-W�S	cƆC�<���.�i9,���5��PA���黌{$?2���Ƣ�Ƅ���T
	X�rH�.R�ܭ4sQ�7;KFs:Q�Z~,�U��P�f������*�.���j��>�@H<��}{����O�mei��F�nQ�_�'l�햐�_n��������!@���4-�}��^�*5"���N8�@nQ��$��g�E[>�M�92bqष5��T���l��z�%�w�1�<MvJJ~����;�ɶ��.1:j����t�qF.?��K����V{E��;�ys�^����HU)� �e��q�jK�IY��$�ਬ�����t�~�#�>=m��|ӏ==J��b��K�8�o�R�}�Z�L@� t��d�]h!|�Ih��O��C��>~gzr��K��ч_j׋�=״����:XkL����f�^K }��}��K����[�|Ķ-�,�����؋c5o��4Z�� -�s�Z-��;V�:�i2�5��W�ͽ"n�ϣ��=��0�V�
(9N�� |0p3�c����qZ�'g�� �b��`S�c�9��έ��eU@�%��J��wM \?�5t����O�-�Q����Ni�3�8�O>�:�S�W0Dݺ�<=���.��j�y/�U4�мR��iI��(���я���X3�;~2�kS���8~�gZaYH8� �m2��gJ\��ƕ�%�E$���]<M'd�}�f��)��,I�B�l��K��q�'>�J��:Ǝﯯh���c�e� u���ڸ����w����<���i���	Y��@��C$Lc�'3����aFB��|�4�+�%��&O�XF;�,���<^V!w,�6H�NC��}����㷘���%a�҇!סz;�cRd�Hl��p-^ y��v�~k��vu��3˽"/��Ws�R\��C��?j2J�r��w�����M�κ�f4r���Q�+��D �\��LAi9�
��|�������̂��f��rb��~[��I�^�F���4R���1�c��/HR����Ii�Ho44JM=*�DX�9�$�X�3�(�x���>��i��[��r=8�T�I���Ϭ�v��C[㻽pﮕG�w�2�e1��":yW�k�:D>�i��@s(K�z-��oa��1z�ؙ�&H�����R\�0�3��:����xPj��W���i������A#��B����h�$��-`�Y!@�w��7�Jbb���o�T��=�0���WUg��p�HD%f���@�1�4d�i"@J$^>b����\��i��W��g�8�QX�Y���kK�k��w��MC�s�\�u�������=�L��Jп�0P���E,���u����J��ȇ�x�ߡY���v��	$�4`� ��������#��я���q�G)�ߙ���S VR��i�F�$��<l�U��<��k���TY�W��/I�	��$m��s�Q�2ן����j�=h�D2K^��a��m���Ѥ���-���K���&�>[�<��ؑ���q릚�}%tI�q��VXHy6���k*�}��\�އ��uK�v��@M)�-�V���\U�X���2׈�w�Ql��2�%)��0�b=y�WN��t�?-�o̲���HiG�Sծq�:��Md��(�uya�)ǠS���>Qj�I����!��Q�<���g�N�Q��9%O�𣭵��ܦ�a~\>��1�6n�H�L�/=5K,��,���ȳ�}J�}�X�5�ޫ�/_\? ��ϴQ��߆P0;�J?9wq�D��W�������Ӭ������P�����AOq��]j�9%ZfJcpg#z��:��֜��Ri,�"f���Ig<�+�:��hM�cׂ�7�-H?y�d��C�/P�+�X��aR�����D�`1T¯򓄹݋�Ġ+.�8��F��.�I�84|$`��ǝI�\�pf�xG��k�;c�^��LP<��u|�{��ヾ@��z���Q� �����!F���}�]�x�h,��v���w�`�î��n9,މkC��2A�P���]�$���\���7 �����u^|(���P�Kv�r��u �`�J�gTYo�'V0��q3o���p(*�� ���*9{����cjr矏	a��9�W|G���,��<�b��j�� z�P�,:�c��r��f)[����B������`��3j����r~6.�S�Dn�؟�R� �k�v��]�l0��DC��Z��8Xp��{�;d�|B-���iimt?������U-ļ�g�Ż?��M�k��5J����ZM�TN��d�1���xDC��8��scs`��Srq)^���n��@����O\����T�|�2�~��ia�q��j����֘�0�)a@70 �Il��co��ܝ���\d]�Ѯ�Ql�.��皳��O���M��%fo�\����c^�(�]^�������|ᠢ�U/&U8���� ����z$bBv�*��W_�2�(���P�dh�b�yJ�5"Ҍ(&5�Ҹ��1���:��x�*��b�կ]�SѦ�d}�!_�g4��OK��+C��xFa�m����7ܴ�=K�^4y��"T�t��m�N��NY9Hc1@F�"��q��M蜋f]����(�W��$�&Q��ޅBצ,���Spvkp��Ѡ�Bf	�σ
R�)q���EDb��C�� ���y�'���Y�D�SG!U��g�b��+;s5�q�>Ȑ���F(��IlG��u^���%�'&¯�Z�eIv�a��+I���-��@�I�܀A�]�`}�ʓ���.(Y��E��� `
r�^Y��?���+�v�b�����P�<���]� ��ן�=� ��`�x&�"d^�!R���v�����{�>x��5=59�J���5�R�	ZO\Z��'1LPQ�n��r���;^�K�Q�ii��C����r"[�kgB>k�r��U�v���1��z�+�rrĈ�$)LT�r�8eJ,�n�w>���(��M���J��%��+�_0x�����-��T k�<{��N���W����	��n&n��Ɐ��q��b�J��w�j\���˺4DW�W�
g4��R�|��QN��Vy<:o���,���8S���(�`ÐK�3�`�r���\*k�VDqǀ��T_]oJ��!Nd���~�ǵ?�5���G��Mﲋ��p̩ͯ\cZt���*2V��H�d%��'���_�,�a	32�n'��J�fU}L�U6���{��T(���Z�b3]�5҈?F�j1ҥ4���e<���|�Lr�5f��ŀ{Dc_p2�h�v��ޠ���*>��[���1o��:8�z(<A��^�*�2�U<�(l�	 ���~O�ه��R�L��İ��,3e���[�-���2�GՈ����K�Ұqƫ�*�WE�y���Z�:\�epw�m���m`�),�I����yt%�W�L�mX]Qq{q��*-6�cǗ�V����G%<K�cm�q�3��;(�ӥ/���U��_5ak�1��_����-p�����Z(EnfDw\���+W��<6�p3"�OA�"4G�e�76VB(�)�>ǰ��8���% �0�
g�6C��n��D)�$,��c�{m�.��9�h
�'�B	�]�ǰ�G��l��Y�����  3~`�zp�ҟ#_�0dBe�������ay|c����L��W�(ky��(�E?�!�L�e�����u|����a-��jd"��ȡY0�t_����`P�E��X>�(f�#��Ώi�\�ח=R�z�s�}?*�\� ���P��o3�;w}T?v�����\+r�x-��d�u��2�#U}���j�">)�ɨVh��4�B_���NU���ڹ댜�ߑ-����d'8Ȣ���M�9��(�R�(�3���Yb�ǚ孓0C���"�@)��8uQV�5]��5��S�kxb��#a���7If��U�x��Ǚ�O
�6[ҸA���,p8�rF��]�_�����]�~;E��������y�%q�~�໢ˏ&��
�+�.�;	�E��e��9��ݵNW�B�!�a�<L����s���|�-��J��4 ]Hd�q9j*��={���i��e�>7\>�����o�CDk��t z҂>���vk��;�iH��W`,��NX
:�B�B�Ӆ���l#��ɤ�F�q}$	�5��v�eft�t��/{"�}y��N��Ð]�	j�	����;�\[|42 ����7����ۦ>�:�4���(#�TҦr�ų�2�����tY&�;��(���.�r�9�x61�h���������ʃ�)�xA����5v ��A\�W�B��`��Y�kVA���`�{����a ��p����	▼R�Č��H	� �C�Pi.AB�!A�4)��`�FyJ~�1] p?�h���i�!�m��݊�-�θ�돠��;�pjtP���}��fAZ�K=�,ӆ���_v�}���r��n��&��g�Ja=���XP���ز�=�(��-����5�Jbx3F�Z^$L�3^2�1��{��s��@����@�U�	�Z�d��73U�{��>.B��,����䥖P|���DUŶ~=>��5���`{����U�(Yj����W���
�����{�L*ľdxyɪX�46&�WjD�� �v�n��NS'L�js�B 5� ,8:�t��O-���`;j����[_̦L�X{k.���=�@ř�1�B
�uk��͚=z4��-AH"�!:���C|z��#�2z�H�~���P��K	B�ͨ�������hE~�ڛ�[wgB�؁�8�y���4f7�]֫�ۍ�Ұ�V�2a@��P�ꇣ�)щQ3�^#��;3\�������_���w���i�M׭���X�N�l?>���p�%��.�yB���6E8�r��?أ��8�wx�T�5�k;��oG�vf��϶�`#�\�p�8b0l�G�����1��xwĕ�YRs�9{�j����W'�+r(�*�b5ua�I�Oi�M�K.)�C5�
pqY3��ؼ,��]��s���0x��aI�W� �H�E�DMn)�X$�s�z���������ᜢ}��88�5���{sD�¡��0$�#jG��y���y����Nȷ]�d�!*�b0���,f���*q�l㓣���t����(����O�JΡ1�4(g��7	�b���;4_�Z��/���̈́���V|:T��G �/���dG��lIE�g��Ɓ��d0�<�J��Q��P�d�vڻ��i�Sfں �^���p���e�!����ɹ=�w��E�� v�T_�)�h냑o��c������,�H�
$�ߜt�!1ޫ����0)ݷ�a8# �h�ٻT�%]Ԩ�:�#��Oq�H�n�&� \��`���Dbr9���5���M�0�vm_J�-e�����JQ����!���a�:����v�[���[Jip$��ef�,R,Q��s�:"�k)4
��'u����IA
�B��J�N(���և^Č����.����59wB�T�IW��P S�|ͪG[V�sm���u��Ym�Hѓ�>3$�>��+d�E�zV��q8�(�"�U=#"X��Ys�]|⫹���~b)����4�'r�EE]�+Wf�~ԅ�a0��C�\��[���>k�T��'V��w�㹯�~eg�GBD�(@8�S�;��*_�u�S��0�ih�V���m��|j���u�:�PA�� '4g��:ms��;���]���J��p�b���(�tr闒�T���r�����h$��ܭ��C^x,��j	02]����\0�
��g%��p<m��F�����V�����b�a�/��N�Ӹ|{�Sd�	i�e�{-�h���ۢ���Tִ�{>u��i5gڱ>��(��g$&8"*D��G�*�� \���n�j����朔�6���b�[�������Kd0߄3c�����43�ۏ�ԇs�.R���ޤ��*��LA��&��#��?��D�&�Ls��.pVk7�y��4��3�)�W���lkR�:��6n��[K>2)�u1�A4�{6Vݶ��"�!�zD9��tJ�.�����I�S���}��� g�K��U�M�7�$���I���2ɘ�b�<|��56��}V7��|�g�v�L�եg�������O	35d��a�Hj9$��1�=B}L|�\W;�
�`G�P11��Ɛ����/��~�yh��A�ώ�IݙpXK4���&�����Vn� �3�5~ ��;�Aը�_/Ѐy%���]�]ˉ%�JU�:��X���u�KOа���FZ�FF�<l�2�׌��>Pz�N�W���δR�-=�FIϿ썤y~d��^_���g7۳�W��0���ͷ����^�u�~���j�s9g�
Z�v8Ly'����Y�k����_�K����7�7M+�젅5B��R*o����M�!*��i�ß.��_�tB�L˸Y��oxؼʳ��d���(����W�@8ur�!LJ�y���.A'�\�����0]��"x�炚�#'H�W9o�+(Ԃ�*���s������tr��� ����⇀�*��X��Y��R�����b8�.�B -���IH�&����	��#	��gj�$����a�ǟύ� ����6r���@���Hh�B�}���d,����������|k�P�޹�ڦ膃iZ��޶�t��Ǣ��:� {Oj%6��1�,�W�q*�`�H��Z�f[Fn�pI�{�T���ޟ��R�l�oބ�a?f��K�{bP	U�cIu�c���]T|6���+���?��83e��;G��i=��!����
<_� '�VKwS�,6t@p%�+���ά�``P��_��Fl�����w��!�M��0���֞�4ta<����?�am	���Í�i�uWy���(/#QT�^B� ] �Y��צ^���m�܁���uG��3�(�.��<��Hxi�*I���-D8\lpu�L��Δ���v�!"s���T7�좄�l^W��sJ�H��5f5���j1[��`J� ��Y-��L�e�Q�1�r�ĕ�*���ه�)�@Fՙ/�%R顼t����-�o���7�� �ƛ񌣫޶V�	�pRYߠ��x��&ϓ~{�O`W����YtR��Ԑ.�@��k�(�a�ˮ�~�ж���I��w�}�l �Q(��У1�7KC���d4�6da2�`�X+y�T�N\�i0���&���)�ʮ+<s�_�o�O���j�c�K@��G��=| ���u��3u߰����C?��B}�=� �H?bж㌌Q�?8Y8$6N�U�-~�QV��{e}�U���m7����:�u�M�=x��ͯ�j�U�a�/�>POF1K2&-?����J�x��|���������?'��C��٬�s�{!{
6C-1O�v��p��K�D�;����H��ޥ#���B]q[Z�����T���ݥ%$<F�����j��<x�E�V���3ce)\g��(8yu��f���$.ޭ��N�m܎�o�g�Y�~�h�(֤���I\5vQǇ�D����I.�׺�^��۞T%��ݗ�<�ȇ��B>��i��m "ƣ|�X5O��r?f����J�g��FNG�jްw	e� �Ձu�/m� �`4W$�B��d�M���.�ZC� ��;^��C��Fu�4�ZC?���u���<I��G�WY}Q�~��
�|�G~9r�D�1p��$�[�������+RK}�D�ƧP`�3��l�-��se��1s(J��*�:��c�24�sW��I+����0�rI�9�p���޼��P�j}͛�ûJƉ� -*]�>aD*�q��������'�&�E�+���@��v&m��1���C�޽j[^��~���n�2t��#]�り����&i�e:�˥IC�꾨�����L��đ[����2?�x�e����v�3�M� >D�$��xJ�8��1���wH��*nI`%��a��ա�P8ڈ�� ��ӣ9�9���
�]��c���fUp�H~
�r�����̿�����[{�X<��
�ZԽ8����%`�-���h��y9@�G!����u�1��JS����mnHi<��Y�+�-(ִH�A�&�V54$�`�@t�����Í=�[�=�,�ΐ�i�9:-�ڜ���b���S`i�ET(�=��"~lb�e]Gt��g��`��J˕%�z�W����Ѹy��x�$�="����5��x;��V~2���dG'���0�2"~%`(�gm���K[Ks���@v0e�Py!3�gt3���`�a-��'����d�f�X�ت^m!��i�g@@=�̒��%N��x�d�X;e7���&3�� �������R�\Cz�G����]�Swz�M�Ӥ�P�7���(�\�j'1Ӄ�Io��\1yO��Ľ��>'�	���CKB�7�r�켚�L'X�+6�M!�1��9iu>��U)6��mt0�vT�ԣvBāg���������):ه�B�z�}8�fA%�'�	���Q�A�D�pJ��U�2�ڿ%��`�0��$��c"�5�P�O_O� ��u�:�gueҞ�?�45���
�?9�,�M-�����d��Ժ����>�&��is�Mn\�$>E$�=Rv~��D�Q�y����~w�.���Q�+U�錆���aZ���u�$��0=��U�Xl�g����,<�m1�dj�K�9E��K�� ���.NA�
��_�{�}����`��sl�3��9��y
Me�Q&L?��n��=\B����{��C�=?*���ޝ�J����h����(��0�Y�LH��\�(Q���=�J�MѸ�����ז"F;�IAxS��x,��w��?����^6l!?IS� �C�*T΂fZ�]��HQ�m��\�b�P����#�=�j2��\N �����O�p�4Yu퀭����5Z��$�:�����(Azu�����˷��Y&�
��L{@l�fy��9a�:P!��Ӏ��$;���H��@��b��Qؖi�+��BtԌ�vͬ�;@�i
�@7��0��\>"�s�.��x�o�
��K� l?�}�N���$�$���e�ȹ�J�6).����z����6vo㢞41롆Ae�!J�hY����,5' 7��������i���guz�����~��j!�.�?�9�0�K�r�����
���0D$�j��S����?޺���
k�^TNp|4\��֓�����s��e U|���������Ux���-"eg�<tq�
�/��֦�)L�F�=���ͩ��2ش�����0��̕�|	ػ�¸l=B�v�b��\p�\�R,�tj����P�CK(c�K�ҿU��ڦ��cH��w��@���f��7;��дћZ��jz"��T}�gO/�䕓�FvKyMB�+��[غ˸��ݖ+�����\*�j����Q2���tԫ���qE�β$見�jǉL��8��sR�!�Ƹh� l���7��t��_��K{̱����xAV6S�)�� 
��cF��SОB�>K(ٙ����;����~�;蛰-$0��[���I��v�g->f@�[��g�Pp��Ht���'�SL-��LSUhlÑĻ>�/",��8�G�ѴN.F=F��X����*���+z�8�g5�R^�	r�-�����$�|�QT�1��NmTkY�K�x�r$�K��4YE�ؙ�R����#��a�,���Kb/ΨD���pP?��s2�����&� �Ϝ�y��Xb"f��(�~Hr��P�/�z�m�ݦZx�x���&��s�(|�Z�x���C)[ǯ`Z8�vS�ҧ�|�@~k�F;@:ׯ:îJ/$�J�F�Z��PSP��ʛ�]��&�,Qr��:T�,r�� �f�s'�6��tZ^�sp�:l�Y�/��>v �(:Y����m45:������a�|t�B/q�W~�����s�O���Zv�o�[�:W����>l�d˅��[.x��~/�"?��}X?�޵l�j��L�Y!K����2�����
H����@'ڒ�g��!�Z�CӜ�J��h��Z{�t*Z���S��ֽHa�Y��3g�#�ٍ	J��gJ��M=�Cpts�
P��䟞ٛ���n�$5P��9T��=k0p2p�f��P��U�p���;S��{���o��('[̔���ܞbx�������T���4S�{p���K�d�k�Z1���/��/Sg��Y�=�Ձ3���>��+�ާ�d��#_c��}���eH%y)��D�"F\1��/=M�pR�˱.
d)�&l��o�5R��uhZ�7�	2�%�N1�l>�m )ޘ�.�b����e���2�U��Y���X�d�}�4P*�W`֘��FwF�S9���*y�EM�-����9B0�L��?�������K[u��-�����H����V�~����j�"K�;�HFa��;�'Kt��P�����5��8�C��'t��Z��KI���Gt�J|�������ٖ�0S��ƨ��Z��Wj�?-#q:5a�T@`u6iVp�l�}a]�PFz���J�Κz �����z��:�P�H
,�6˚.����n	z�'{S��B�MI�A7@i�+�g?�{�5��˂ͧ���I6�Fu��xŷ�'�
Э��]ھ�Hh���J,H�T�J�5�&�|���]��<q�0J[BEC��1	�z���`ydm�~ߔ�:}�p�*uO	��v���iMջ���2��s��L,#ҕ�)sb�B��,#c�Ș��m���?Ni��Qtp;p;����s�-�._� ��s'������9�����M���rш���@��tfO��*1��z����%t��o���o��M^'��Ζu����z�k����1�V�x�9�lP���8 I+�t�����GPu�h���mu�9�W������s��ۣ��v4��,���u�k�Q:��FM�U��<㳽��4�a:��ӭ/� ����,�.���LOa��?���*�3 e4ݹ����<>�Pu�0l�y�)w������A_Պ�.W����;,P�d�XB�n�s���<A#Z���&�)�49��Uӛ����k���7ֹ���	f�Dg�� [y�8�v�wvT��7�4N|�tT@�f�<}��/�Uu�/3��{G�\�E��t^�/����+d/л�>W����H���C��1`tj�������]�An�$:�	��� l�eP���}�P(���i�l~�鋿����Lp};>@�!�����A�j�����E%�sA���L�NE��KywL<)�Q�����.��5j�y��Dz|�)�Ƿ�C�ʹ�{� Y����&�O���s;��,��g� ���y7�V�W�.�G��L��4��z���#i,�}�,z-�zW5es����Q/�:����d1�u��E����{{I����<`����r����2��"B �_��D=�I����d�+�"�RN�%��ơ-�[��}�ƣՏ;����&%9�@�3��O��2ҍ�%ZmM����>�9���Y���|C�I��X�P���(o��yG�x\O�"Q����K�a��TM��5Q����R�brS��!8�v#��?���<�éXm��h&��6{ 0h�"Kr���6���4=�)D?�2�z��hي���^d��{+�(��� �)\�뜡� �X2��6ȗ�KΏ�'��q�k���Y���ўS~01�4�_��5���HWό��3�������5o�^3�3p�a�a��ty�(%Z�R�d��I�/G`�J"ȳ�9*@������B1���TM�:A��DtIX�vMJSkIGbiltwL� �mP����Y(�i_`�`�3K��-����^\K�j��j����:��؉�죘�_&O�Ģq��;�2�L�����h=�Y�2���d���0��3��ܲ�%1��9Q>kS�E�A��Ô��x t��R���˼vt�Od�����}b�y�3x�	��@6z�qH`H���߈b���${��k9��,��O��V�\�}��G�_{�/�~���ː�j�==Z�B&�H�AAe���s�e!�fk���l�^	����Qɂشʛ�?P������~�N�$� P������Kt�(��U��j� ����=����zR�L�����>��+�U�:5?��ݲ���vC�7�p��N���'�hJb���P��(��)���������B��S� U�[>9	���q����zn�2$S�����i*�"��eH� ���aLQ�"	��ae�}�/�s�6����ƺ���<��m[v�IlP
���Z=l�8�w����]UF����78Vdql~W����+�2�-NZn#�mn&���M��j;ík�H�)9*�5�����I�d�_%�n{,$���4�h��z_y<R�=u� �S[9��P,�y�I�с��;�7~�;*���:v�������L��WY��`6v`ƫ��O�Hf��;�{`�����w�CLD��U���W�B�׷��q#�g%����&j�x2��}��L.x�;0+��D4^�2"V�׵S�>��Z�A
�e�,��_�q�E���}Ky9`��
$5��8�� HT�tй(��5$�q�^� H��KU*O�+O-�~��p�Q�TAx]�W��[�h��Z�-"��Mo[J�F��t⍳�[�܊�8tô!y'���H�`�QZ�g���tH�����3��e�s
s"�5�X�P�f;.������u��� .�����Q�U�ܥ�R8k�g����(�v�fd��^1���7k��KqW��4!�q�و��4�midT,��!aU8ד<�Kݧ 4�ᐜ<�Vk�xS6�_��}�P�
$��v#o���j��癑�`��˾#�ޛq�ì��j�`�ZY�Z7(>�z���֍�5DuÚ�J'�%K�1���<�꣒Y��-��)��'��W��i-X��f/[��}����G����@C�����Z$E����Gz㱉�L%%
.�!4,Czw{ n�ȝ����}R)�,���ԇ$"���W�w��5^�>���.�}��9��j4,��0٢;Y�Beƭ����m �����A�KmޗQ(�\�;,�P���a���tW����>^�"�3�-��x�:������<b���.�\���C� !ZIx�S���W#iBp�Hvc5�F؜�}׉�q	��;6?�Eഠ27�S�k)��~��$qj��������Pt'2�)*���"���NZ��qd� ��\?�*�s�bZZ�T#1���!����cm]?�t��9~��A~�ާ%��Y��~�F2�b�a����ĺ*������}��E{da���$(���9�f��Q�eG��:\�V>E)avU����WbP�k�p��VK�-��ϰ���V	<�O��<%����8���YE�^?���ËC�?��eo��c�8w'���uW��⏎�*]6o��	��Ӭ*��×XW4���Nӿ���xGLO��H��hA��BC�T�6A��%��h
[�#�4Jg"-�4AAC�[RzNWì�N ��j��z3���9���Tr1�#������z֒�k*��7>��^6���V�j=�9[��Tu�L��*A2:)�
��a�K��rm���[@9a�U��D�,:Y�5�R�l���͇�;�S9�4�|<ӕ'0���}:�;s�G��U��+2���`vn�@va;�b	vD!��<��7T�*^�U,�#���M!�v�Fʅ�M������Ѥ�f!j{pp�U$��A �Q�"-W��w��b��Av�'��{(�Pr������O��]� �W}��2�����R��V��E�>�	@<�
 ��|�蔱{!=���IO.��a�<�!_�"�����IR���������^���X�U�V�*�d(h:���2�f�"K�Цu7~��B�lQ]�h�y�"��+������f�N�|��,��x����6P��[ꪌ9�%�$�r֟h�#�9B�|�	��,?��6���E�ijLk ���x�y7�BēJ:=��7��|=P�OA#�6����\�hr�/Xy 6Y1s�6����V׃�TD�`(0�NMB���?Tn�f`=�w�ϰ��%T
�Q�qO��в"����7@#f>DedL^�^���r̟�C�up��S�u,c���`EL�'���X@21f����CR4��=�Y��AƵ��"1��րm��pH�>4�=����4-�h������*�}O�	�0|�r�~?��,��b�V��p�z����Y��ȆK0���7�8Lֈ�x� a�  �G&0	�7V�fѩA�E��2�44���b6�X!SarG�a�?[���d�^��nf<��66?�^{�Տ�6w00��~&HC1�c�-1L���3Q��Ш��!|1y݅5���w2�,ec���BC��?�K��c΍�=���2����b5�7��j��%�M�d��X�P��KǢh���uñ���e�٨��J*AG$�bkX��|~��Ӊ�B)�2�Ws�7<j���[�Ir.�>��/
;�:����#�2֥d�F�@��p��L���W��k߫�>wik�+�KI/�GZ�3o���9��7���@/�1b9Nq��TV7��u��re�6�':b~��Q�+��x��)|+����9'n�l=�����v�/��6u�iB��[)no-P��҉�\�8Xēn���V�<���{��� ��:J6o"�KYQ�)i�Pt'�A��R馛)b��/zQ�S�kP�7l��|S��tY:}ɇN���l"���Px"�O��8�nO��|r<з��S\T)}�0� 0O��Rz`�XtU�����I@�cx�N�-���������������`oh�^.�Y�6��@b�X�3xuV7��y$��]�����l4��?C��A]�Z�R�mZJ>݀��Fj=B�cv�z���/�����*�bk�����&�UFd��Mt.<�y'����2 ����ҟ7fmLM],�/v��'�0;�Z�-+9}�k��έ{�1���8 ����2o�W!��v�n��>��C�Ė�u3� S�H�����(�����������Ϛ\_m�S�gA�=��

WVPR�-Dq$�n
x�HZ��PM�9�A0��,�f��nK�=cU׮���	���8�l�t�
h'X762}�K��z�M*�
`)����J� ����m3��)Y��Ê�Y�͊�N�ȁ��b:���к!E/P/A�X;,o��/
�J�6�w���j�c��7�l?�Ś��Ў���6�}�-y?�����[۟��e�71_�"� �b��v�D�Z���\�[�Q���K�	�r}z�ڴ3�|UM�?m�i���62�Fn�>���q/o,�w�t�yth���q��&�d�Q��PmJ'��QC�>�F8����_�~a��v��!
�e�|�`m��o�K��V )������9%��[✯S�Ȼ�I��F �x��-�HJVNH��#!�7%C�{�u��d�tۜe���=8ڲ�Q��v|5����M��ăw�=�_�x�!�\R��gB!���cT<C��#��%�4�4�p�e�8�]����Wm���w+����%Z
�U�5�i�ղoJ�� �s�G.���u��r�,�c�-W���x$���c�G&c�[��ݭ�G�	�h>��I j�O�Hy�i	�\g6����{�m��.��4�i���J�&�E�GOu�T�f���~~s��*�I���p�T/�|��ȣ=�{j�y�����$���d�H��rͪIsִ$~��x�r+��Iuh�^����� %��L��1}�e��-�/���>nߞXa�6(A��d���4��*Z��� ;˗�/T�ǖ��oYU���o~�s�+<
�|�:jX���?)��zy�$����<û� $c�zodc�)��~Q���P�?�Xs��wעG<g�]�&��u����S�����<�bl�"�ps4��j���e��$�}8sf �l��4zp޷�[2ny5���{�/+/�h�6֖!�9h3C0��x�;��ЧBb��vO �í��I�~�A�Au�y$$0�h�
�#t�W����ζ�{����p���R�n��ɷP�L����*�H�=8��q��4�^��ÇC�u�e6d���]+�⮜
V#��聆�5�-�}lYm�uC|#{p|(�G /JF����k]�בI�Uxꊈ#��� ޒ�?Gru����yPo��`[�%�IY)c�	6�$��F�Q(�@��yˤrz.>3�F޷3��ڇ'#l�m
��H�R6��쨭U�P?%�<��c���`W+��q�_��=׸|a��XFݢi3������̉ϛ̔%��y 9��K�҇+���rj��	͎*u�zT\�]���>HL�<Y���;�j[�-�9����\�)\6N} S�^Z�xK������j)8�������=<���0��\܃ÃqZ�G���N��K��``�%�~ѓ�rk��7�����}=�����PY�����Ύ���d�lb���h�<�`�����D�۲�-9,���JNG�8q�V68��_MR�\Q�[�1 �4� `n���4��8�ԱxJO�X]Ru�wR.���/�b�d1�+D�E�8����c��@�rW����o|^#D��.g���&c���o����參���g*���ɑ��R?gqv�-l�(ю�w��۲Nb�-�!ʹ<�6�I\)a�y �O%�U	�b�����+q �k�l�!��d�P~{�KZ���+O����'3_����V�ks�I$�g������`���0��z��}�Jn��mœ�^��Fpm��]"n��l$Ծ�L�N���6X�'R�'�\��[A�;5㱲I��FK��m�E�7o�{��L��R� #�1���O������؛#P�����O����l�ɂ��uݒ�O��<zE���t�z�bm�/!	��"�%�����E�m�-������x����e� p�=?hI�����B�*�]�ᙹ�'W�.
�͋̈r��W
S��m�ϰ���ѽ
��dL$�N�d7'��UN�A�w�e�i�Ok�ݺE<6�ep��a3��Q �8�X ��k��h;}�3 �qre;_���{���D��D~Z���
�@��7<��x�%®qY�i��ʤ�jX�pN`$��3Hv<�:�4��nXȢ�r��r'��\��mޣ0����S�O���"�Ldl;z�[�f�Y���\)M�8�-��Tbֹ�p(�_��w��-}��m��"X-�pn�[�a^R9�
�4���î�ٵ��c���v�Fda���z�����2�6=18���X��q��zf��<���B�f�� �ZN���+[b[��Ä�<t	4R�D8�Y`���v�q��%�$��r"�� �p@t�x짟` +!˼�jWҠ��d�&q��viKh�ພ��+
XX4D���f9�����o
��h�wJ�o��D��\ֺ��T��"WPJ�,�T��E�. �g@�8��]+a_?�4���uR��r7M�ḍ�1�uo5�N���c���Y�p"��t"-�_�����$꼐E�@h���B�B>�H�'Cy�����<-�O�����(Д �`�M��{-�z�	��H]E�D�E	J�_yť7���F�Gɋc�&Ժ&�1���W���蒋���g+������#�R�Fmj������zY��į����"��}h����l�~HҰ> 1�լ}h���Q7�3Q�" ���<Q�M �,�3���d58. e2鍅�ٳ�U�1������`��0)�o���竪"?jdؓ�����J�>�e,�jS9��S�����]���Lu5� mj���ն%Mr��T7)p��'k-��K�w�#��gO��+6Dy�r��L�kN� ������[��*��A �����pA��΍��<�bb�a����7Y%��d���º`S]<H-9E�cD÷���N��R�'�\������W�����v�$�*	�� �������tF���<�sQ���ɕk��� ɘ6ײNw��j��B�6�%?�o�,^%��30l����GzG�e+��7U��ſt�}3�����|�U8��yS��9����d.&5�S���%6�yduQ%�gY�������cq"�?��z)�'�C��}'���4�P���o��7��	��9���
x��sО�]�o�kܥ�vX��B5�]��	uC,47`&�q��18Wh+fo��'g�������:�(����x0rS���x�q[V?�i��n���R�7�{�x�U��]��	'\��>#�+���Y�� �T�������+ 뷽��!
�i���rb�����L�Y3�t�^���|`�x����"�����*�}pե�g�̌.|d>H�X(��U�]#p�xi$�ڙj�Lb��33�n��ZqE�ց~=qϏ^���U��{�C���G�p������m(ƽS��#�L��3�V�S��X	e"A˃�@N��\+�շ�L:(���9z��QЌR!�A�>�_~ok0e�i@��7~e�En�����!QU�D}q���+1��*S �s�0Iuٙ�Z)ܾ��T�qA���+2v��R��'���7}�EUb�{2:jO�D�>gŊ0ɧm��B�Y��J=rj?h� �����DW	��(���s~b�"��Y�Hp)�9Y�S�?g��&=�]���w�3��Qp�q@M�|E�ݾQ#�̱Ϩ����6���p�]=�r"��bs�[����n"6�F���s���$18\�q�J�Ne���ƥ��omyV��\ĳۨ��N��r�dhG4��P��v$j���WSAϜ��2�6W<���̱i����O�j�+Zyղ�/�9<Bܖxm�����@EBI�o���s�~�8e_�r��`�D:̐X;��/�R�gBI����vsy�����:-�l	J�&��LO7�;P#]��fږNR"\7n�`��an��x�{�
ԚL����f�� �5��{F}��MR��sh��l���3��?Z��P�6����⃒��V����}�=㡍��.�`��C�\�8s�p����f+�<^��2E� �%+0���3�kO6�%_��sG���q��|L�3���� �� J*�rj$�w��m�=!�Y�}�<@-q�mk�ӳ�&��d��B1�G��Nϟ��w�I$
��B�x����7�]��C�Qp.ZL3���CC*�l�<?�t˿^��e�V��.�������Z"ŲG�Vc�:��j�<8/I�%6ߔ�=_��!ٰ��N������BS4A��v�����d��<f�3^'2�XOt⟤�r�;�+�L��bc�e�"0���F	�[:�ӽ�]%�G�� �U�(��/�㚾ڷuFM2_��[_z�H��-�*A�#m���6Y+�p��|e������Je���`���=��Z�E�\	��Şc�tt����m���ⵚ�8��[VϰpIt�nn/g�GZyjZ�.z���ЮɄB/�pa ���������y���3�"��e��Y�t�4����`_�ʰ�pr��Řlc�s:�n�/��3o��̩�"�QHN�"<wB�8���p���3�w���c_����r�9z4I������$(��1�=�b�׏�uZ�ڼ>�\jX��=�&?[O����fD�D����-D�����r
	��Ts-؊���~�UN�[Q�F4�n��s�D�@�{�CQ���/������TU@�)!�ӝ�^X��s�Ы��\�I�0f�5�-�7����9�Lk�b�����
�;:�+�����J������p��n q�\r,���15�}���r�ʳ����z�d��*5�J\:O��DbѠ/�^i�MA�ż��=~4J�D�0:f�+�F�a�~8U:�F���XLFw��9��}��:G��zy�k�oƁ29��{ƴa��I>9��Cuc�G���:{�}�gE�(������'9<n=�t��^�������걔J�Է���_CZ�%�M�R�W��;z_x(�������uJ<殻ϼ�7���c���7=|:�o��x}z�Uò������H��:���Ho��0��������kpBm����Rg�%J噑����'�y���ejkJu�����{�	U Ӂ1
SlW�y���q��oy��Y�W/�j��g�Aڋ~琽!/n�	��x�aZ#�0�p��=�]�IV�E��ǀ}hW�z�#�pjN�=4�Nĩ��W�8鐐�f�C~��B�C�G�3�=������\C��޵��u���n/��݈7`V���+�vޠNO�W�vŎ$R`���^��7l��e-]�^�%��v�����>TT*�O*����BL�U�_'�)ݔ|9��F#B J߹�n� ]γ����P�u1������efd�<'ے���7�1XΝ8?j��b#��ߙG9|��]�S�,��t�#��2uy~3N���IԠ,X���ŌiGk)�͋z��Ld)�r[Q�ntWd'ql��zbl��L�0��sѶ���d83W��!����=����:�2w_���K�\�]�P��ꁞ����jpS���samƟ�$�����Z�A����j������S0~)�tz�	@Q�J�Ց[
��.ܱ�<�D�ip\��(�Qi�m���)��ٺ廜ƈ2���9╠����`�B�	(H��E�&F�W8]^�������D�{�MN�������elO-��f�ѦJu�Y���!
�%Űf!p����w�S�����;w� P���9�����p���������-~�K��n���DT���������(�S�E�RN��*�P�YPw�x.'t��l�̉��˒ �&���W���h7d�#O����j[�-��ۥƚMbT�ч��/�K ���Ԙ�X��%v=k�OS(m�{�Ƕ��?������^����o8����\�hL:�2j*�N�(�̥r}�Zzb>�8��*1;��O5Wb5����Ç	O�	��WSݭL�8U�ɛâ����+f#��\LT�"��"�dԤ�)X�'4�kyf�&����c��w��J�̥�Ҭ�z���>a�G�H����3��}ѓr8��T3��BT�GC?��)],ˆ�jnF��k�+�W�d���5P�p��?Os��w۵F�H�%x��a�}q,� �A�=��G�%����C.���!�A�h_3+)O�u/�u.���f9��m_վ��AnU�%mAsW�B�M�C׉��}��yu_�B
�(bk�Ux���D>�֦�@�[U��-�� �1�xSa5���Vh�F������u��u���#5����e|��M����3�T�*�6[��C#��=T��W�G�ш5�M���t��Oy�䖥`�xZ17�f���=���R����}@Tc2��Ъ}�%��,�+jk&_���k��I3��&,W ���)�����ęuS�ߤ�`/�ޕ��n��]�ݯ�@ҥ+%�_�vw&��1R����>*��+]U<�=�Ax�����C�����f�.�����9��4�sQN���/�Lx C��JouI��[�	o�#��e�D�[On��v�E����O�f�^Hy_��$�����d.��\Rʝ�{�Ta�zdN0���@��p} @�h'��1��l%֖��L:�������>t�;X�	'�N���.��u[i;�6��X�4%F�Kۮ�R�0�"��q�~��Δ(��	�ph�Dc<���A���m��d'K��h{A����<��'�I���K>^�t>��qeED>�R��-@�W���7�p��?|������c�#V�j�������5�֩�)�����C��=[�/��4z%��2F���Z���� {��D�-L�Vn|�a-���P�_���oP���'��&�7-Y5=��#@��&[�x˦ϕ����w�vp[����<2�:t�7G`y0O]�׻��}�Wh�8&AD]wy��vP�*��/(,E��3x�j��ߘ$lrM��T	J<<B�x����m�dr܌� 
�YS/�����r0�y��~ᵲ�.�$Bk��ai0m�(A*�=��C�&Qȃ.k��k���d�%�p#]zK$��bhG�2���I_U����x�[cJ�5�L� OF��_�_�GaʾQ_�V7[aּ�B�w%����׭��AIo��I/D
�o���.ŷ@	Ŵ���?�}�S�=�OD�!˗�y�/ �64�Y^p�9&���B�s��Ɓ�Z-~jy�t��,|l=XD�q-C���}�=�ڤ�F}>*��W��|�T�K���d�1��*��X<f�L/tw�yiT���b�k�C�4�FP�G0�����Li��ͅBam�̤��:r�r�+6�?,|��Ma>��*����n@쀣\����$��U 9���"/K���.�b~z�*���
\cV���zQ�4�Y�B�	+ �r�����ю���5���B7�t�3NTȈ��ܖꂜ�a'�-�����C8�Fa#OOF��=�X�� b7TuL×�nd����U� ��4\�o�R|�ZlS�3�Uq濘sAx�4��1���rW�ڎhHvp���+3�К!�ˠ���rN��'~��?v9�N�w���C��:�zXp+�e�� 8���u�6��̫(����SA������4=��E�W�����@emXH&�����G�?�n�9�y��>y�q����+|a��~Ɂfv��e a3-eG�jX"cIЙ�j.^�8fL��*U�Ԏ�]m�����Hg8sR$��š
�O��@4�P�a��D.V�^4.�^ܻ��H�^��/55N�W���ahGo��Ƙ� $��h���``j���me����QK�jhM>�z�bJ������
�����&��o��m���]!��֨��j��;0� tOk'�5u�6��4��DZ��}$C�7�5-z�E/v�\�n��u;�]G���Bx�a	0�0k"�*��WUk%>�r�Zª2�sH;7�R��;��V�<���� �8����!p�'��!�M�
���~e1h�GuP��*5�C��Y��'r�q;�k�]�Ś��b�{�ﾵ�.�(�R@r��-� Kڡ^ms�a��yp�/���r�8��1wlwB��>�ڈ�C*E~誧�:���-e�y5q��k;�� Ϣ7��/�&A߇������n��a�E���R���D���@Ό̻�o]�,G�?mͺ8a��yN1�H1DI�^����&��0�Hu�x��2��&�� ����`6hU������d��s76�7�(P�O�ŗ\<n��~�� *�Ɋ�T
�x`���Յ�-w�1��lf=���l%>��[�V�[5�'Wٚ�0�r�6�����aպM���N�Tý�c0V���mH�#�I�cM�{Ow���Vu�kSʹ��l�Y��VRr2B򺖡�ӗ��6�V^͕�I�q�[�]������1>�����M ��_v�;�������@ڒ�>-'�<-|g���|���BM������|^�4DD �B|R	�^�����K���@b#},s����:���X�m[����I���I�t�) (�z��f|�氊�M�#@4��#�3Ol�ێedf��C+b"�Z*�íJ��p��� ��qF� ��^FԻ%Ů{�K��
vBTԚ�-6���"�;/���(b��䏃�@qiNޥ�������D�C;@I�$��De}܏����K�rS0�����X!���"�آM1�JR^u�6���&�0��xLr��6����V()�X������%���$	�W����Q�"�~��L��E��U�L�G�$Qwv��^��xj%�Ώ:�0��$������w�����+9�,!���1���-0�c�iفU9�bjtp�>ר��3Y)c�X>���O�ipat��e��F�O΄}��EɝN��Ղ�y�d�H��49N�%Ht�p�#��W�}mk�0yg_ݽ�/uZV�a�����p�����@B:���PB�d[7�-��w�Э��r���T�A�z���)L���y�������24|��ާ��1��ER�d�'�Ŕ�U���o�5�$�l���&x��!w�a��f�U~���8�.n�)������5���G;�9�ә/�o@�N�N�żR��
y�i@'i�~,�L:j/�k�D���DWZ� 3�d�<�=~1ðe�t��@��H�BЪ�B��\f`K�7���ݨ�g��D����>t�����*G�-*�PR'~�,����]�#<OQ�j�����t-N��c6��S,E��9K����e���u���d���,1Z5n���U����Bl�6k�NE�֡�L�kl�e��t�S>π]�F�]�?�U.�Ъ��n�yz�V�c�[g�i��Sx��v(���^�ƧźҒIM���':@�Y�1�lIj���.b�xn�q�gل;�m�$'�g���AQ�c�w�fߨ@3�gn.�G��z10�iaz<��5Yp�a/]��`��b߻O���+P!��N2C<$
�e�Xs�U/!#��b�>�CNat��շ�'�v���j=bS)����̓M�M�:�ԧ&(R(�*��k�c�D?���Z� 煕�SI�E�7�h���m��/��`n��$�����NJ$8���ځ9AN���y���[U�pҬ�|'�E Ni<����qr2�6��F��2��L�ӈX�����
�i� eq�\�r�p��1Yh_%����0��2�1xi����#iE�/�J��R���-��u}`�d�����N��G!Z�iE�a�T�,�?I�>��b��v��4���=����6T�'�>�F�����U�=hN��H��RP:���'i��e|�?���K��#����W�3������FDl��vvmL!��n���S�<f̷�0�n"�$?U�������W�K�K���
ͯM��˦op< 
���$VOS�T����?���y�[� Ok!S�6j�����@o,G���8nd.TE��'���*9��vq�Z_�����$����>��H��P�����A���j��W��/��2���q�Պk��r���ź���� ���8�;��K8���2��T�T���{7�-f)��u�c�Ày ��X��<jC2E8Í��k��Z��]��b�z� a�u�ݥ-�=7a�d~�6��S*+݇YuPL�W���-�i�{�F	���������ɿ��+b��0�G(lt(�ɗ�YA��[$᪑�k:9]�"==��w��`ig�?�7,�Η�qoc�A� ���	![���<��=��y�����{e�V�q�-}�5.�j�g�~Q��;$���{*�/k�64➾�i�����0����D�5�i1�T��'�o��zZh�J*����t��S�.%*�Ҏ^#�Z美ѳ��K6�Lfw
q?����R����f�U͇m�Y�|���
^�s���<��eH6��h86�ЈD5ev��q!#��خu�_��q�>�b�p�P{;#T-����h�ɀ�W���!5.|�:�!�U��A�	�o|4�w�����5C��D9�YR���D= +L9�������E����ݿW̫��Z�9�,�ݬ��/�[�aފ���0�[Lak�nV�`)�h^O��'{����v�!����Ӳˑ���lk����g/�����*�7��(
I�@�ilatO�U����&@��h�a��r�#�4BD�7�#g�#���q�T�� d4���8���ܑ5B��k����e}��Ţ�����wB2����fEݓ\/f���,L�����A��a��*V ��w�{�u�N��N��a�����I.х�q�5�'&-�SXP�]�H��k�x����p}os`rmo�*�+vQ�G@�Na���6�+�)�o����/ԍ�-'�jz��t�a=d�}�m� ����0lԧ�,���n�Ca��}cK��V�	�RQ��5!]#�-)!,���ת���ҽ��	�\@��~��I��t���������Y��IE�.2 _ I^�TA��msj2I��E�L�}5�8s{�8U)��g@�j�;��{$��W!|W�D f{׋i�ڞg۸������P�m�%\~p@jJ3�����]Q�h������0^?�=x�]Gf6i���0�TI��	�E��e6���<�Φ���7�&��|��V&��b9[\��	��;j�fO|)��i/+�8��igd��5��E��};�*1P-��&*%5�.*�!J���_O�r�d2�Ku2��� �o�����lԀu��pUF��u㖧�����!���#�V��v[v� ����>"�. ���3�!�Q�nWn?�E����t.��T��G�,�l�C�d^�8Na� ���Lo�f|�謊�LEb@�\ם�p/�����;,t��}��E�AG��[�$�y��� %FU�*L�<[-���d^�Nhg]9>w3�a_��s��������5ݲf�4���+$b�����E�.A#�%!��� �q����	T��%���(z��mE|�L���G��ʅQAV�gw��&��L/&UD}�N��g�[lM!I�[����V�|)k��&�9���>꾕�{�w�7
�pܻ��;`��M��v�Ȼ�YȫEj$Y1"��i*��dP���=q�	�XH��'��땓��W�@*n�E�P���۶�ξǞZ�%X�{ܞ�9��{�Lh�5�҄�ku�	S�u�Aw�C?�����i��gV7�ݻ1����ەTZ'a'B_���+ j��:[���=���0���&rV�ёP��R�`p���|��n���ɢ��j��A#� ud�>X�s|&��6D��\�-}�\�u\�����}"1jp����C�}R�����5�