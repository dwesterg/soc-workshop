��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQ�k��s�#��ݎ�4Jh�}������!2����s���kW�YCu��ߥ� q��j3��:��ʥ�C0�S�m�lf@q������p�Q�A����}�X{�z�_�o�Bۆ���rجv��3 �;׽'2��&��yhQ�吮{t�RiF�J�}/n��'/�1���>�e�a�E�:N�c��!�>��n�D���TꡦDkn�(ni@ΝΆ'�J ��0�}uH��[*���q�j5ɪ6�u1�����n���SUO����)����زl�q�f_��r?x9��T_e�F��MՌP���t�n��QO�����v��d�|�RO���@И.:���!�D��d(<��<�Ewɓ���;���(k��wB������1��;s�ĂA��,qhi�d�a�M��>fԾ(͆��/-���G�����}��˖��((����\G��/���:]���H��m�>��������9~_Xaǝ����|�MeDd���>K,�J�=�H?���GYxc��%<yi������Q5	�P�>�h���h)��^�³��:�[_��HR[-�/L���U5�[G~;��=�����ZΧ~l���`5 ����;�>��ε�Cx����X��@��N�Q1�[]`���b���
��4���I.���9���hw��1$�ö��,����3�q�{uׯ��WԽ����x�e�B�<O��Q�Z0d&�|���/�Ȗ?6��°�I��~���4�ZK���=��6����ߵL������DN�ȹ����H��kQ7.
�h)1s�.W�.�ʟ8*SFGJ]��7�����nm��XX)�4&��F\�������|(�Mo��eA��}���A3��S��.ZŴ�5�$0j����OL��GRH�6$>�j �!Bs<�n����f�����)'�$8h$�H��a섂Ł�3����ߋ�Q�57+���B����P�_���V��M�q6R����!�O���(\(��#��|~���������A������~}U�:�F�R,��]�(@�1�0���Ͼ�1������į��07�8/'��jT�|^�)T��b�C�4j<&��A�����Y���]��d؛U��j&��e���ϥK\BH'дgR���%�r�c��a�3���R�i`�� mC` ��;(���%��O+�>�g�v�r�'�m"�lN����αj^j;��CZ:�S��g�dB�	cɳ���ׯM�^��ք���j&'�W#�8�IAe��J�<'��Ҡ/�!�����P��n:�;b �_3%	x�+���{=���4��6�o9\����Q�otEp��U�p����-u�q7i��OU������Ht����B�F-��@&}������6�x�B6��8hr+��M��Gz�l��Q`�g����6/q����a��q�} �qe�ǧӂ��]��$�̓���2�E'�_J�z���C��Y��f[�<5I�s̵MEM-ʻ3J�2�iVB�N\7.���������Y2��=���R0��8H6�]��htj����Q�q~�p}5�%g�'gJ{�n��u��3���T�d6�<�AZG��r�����]K���f	$��1}��p��������DƖ��߷O5h_k�CͲ�v^}�	�=�_�[�]|� h�W���/tEv�s�q_7�LnMp���(�o���.�q)����gT��������f�b�I��.�C��;��*�t$�-�L��0{�m��q��ϒ�٬T$�+�� "$��X���]O�N"w����Kx�4��z-���Z��`.�]TՅf%M�v<d�@aGk�~w�e�sN�g����j�V��^��Kj� O�u�����׻��9K�
,}�����+F�ٮ@=��Qto�����m�Im�H�3_������/V�{�'�U�h/hk��y���}F� �i�u�O�IkǤlVf�:��7N��W�~�N�<K��i�0�0�nP�MU+���G��k����(���V�Y�!.�D|�%�<��tR���i�<BR֘���y��ny���8��]�9���c�I.�- ��6���NN����Ѡ�.�W�9�����+�H�lr�gb$��e0�Z�T�5 /[�ow����X�_]A�Ͳ�U��n�O/�F���ˡ5P���_Է?�_]�)��R�8�K��@��HےL�����8{\�'�ױY9�o<TϦ�S_�oqz�z�f�J@��&���2p�b�3��Ȑ��G��w�qp��J�x�[���CN�<�c����o��l��)�V�B�~���-s�d�[,V�����������!}0Ƥ4�x�J�b"�����L<f�ۆ�-��>[����8�=���[�8逬�6f�s����:��7�5�p����5��pSUۼu(K�����4��3��*Kib ��]SQM7	{uf�,���r�����O�N]K1�����<S�5ql\�m��T@�5[�K̤��-�{l\ �;'��I>sÅ��]�b�2�Ȉ������FD��v�������K�a�Gb��O� x�.�j���+䯸Efcl?�1]�H�j@^�<,Y�!C/Gti�wȚ�Y���=1)j�c�sY�
[�f
~n�2W=11d<��_�>�Vk<��[�ҬN�NG�k���m�M.V�������Z�[�H6K�Y����LKB��w��$�}�ZOJ����E��y��x�O�q;��!���aP��"�[6?F��fS�Bd�m���ǀ,\/*�D���b ��c~v�P�c
�)F6���7S{Sn0+��{c�رA�ON�,��N�79FzH�D�|4�Dֈ�8k�{�ǉ�t�Y?~7G����V��Ǌ��U/��o�V�۠A��U�D����Y���Ubg�
�łi�|�	�K}��vH븩�1+]�OӰm���$�z�V�);Au��#>,O�na���(��7^}�,|���2�e=7ѓ"�;����i��3�q�=e�!S8�4�����Z��N���T�+uzJ���nG���@͂��`Ke
�ַ6Y�r��>�_��06�	�V⿢�����)�������ẇ�Q:��s��#i.�`���W4��R��zA�E�L�k��Afk(ح�m�/椚��!/-[A��eu��E��	��b
��iF��9��Q���"]�U|�B�8R=&N��al��R��ʋ=�m�~�^��#�������{]9፰[���֑��&�ៅ>W��U<4��]�`n��r�!n*�j^���[M�Y�*��k-����(,����:U	�ö��)�?v9^�y�n�"u����`M �Y�F�hO��.��Ė��!&}'��t�LR�Eb��$M�aT��/`d��F��˥���/��N��[�=Q2�����y��J�"_�B3�g�x]W�)���ľ4�C��BVg�!�^cx�)�{�w@ǽ�r����G]&�,�y.j��^�{_R�!iηL*:� ���i�D�+��`B6>i1z"�gM]����oS����]M��PJ������q����P�-���X��|� >(����{��n�A� %�0$|��M�7���$V�ڥ*�X�?�;��rԁ ��ז��T,��D�A�sHV��0P_���y����hj��n0�]뀰����
��Fy��a�Η�
#���j'��dG��7����1�/33�)Ad�ZoP�m���kGو� u�^�cmQmGj}#��������a����K�i�6т���;ۧ�8�L�I$3��!���N�7�g:�����nV�%�L��������.<#^i�Mi=�b�m8�4[��}"�u���]�(E���?���kv���\�X�жB��:�4�@��s���������m�^X�l�
J�������KL��Ä�q����-�,�MŀI�E���,܏.�lx�s_�0˰c~n�/�u��YY'E.+x뙦����s�Dg�g���DZXl�=���[�c^s�ZT(J-6x0Rǘͼ�UQ����������5-BI��=�,���#f�%*V�m�7����|F�d%H̭��<*�jB�v����S7��f�aO�����Go Mku���ƥ5W��.>�gCC�G�u�S00�)q�oB�_7킱���<��s����33�����T��RM�1si��w<��A���A&���
g�.P����ע@���R��&qS�nY��F������f^niS@:sh!�B�U��z��� *L֫�'���pR�%�)�Թ�܄;�Ȟ����E5�}9�����BAWN�֑l�ꩺ�=���y���Z�;y���Sڟ�Mp�<�J��{v�0�0`�Dַ)c�d$A��p-R�Ū&�x'� ��K��DYNw�rQr�ֽ���yc0�9����i�'��Gl+Li[V����:�E��b�� ��<����J��秞ܰ�e���A��?�֯�#��q.�R	[�I@~y`#V�-{JGf$b�=���Ⅽ,_��K{η��wkWƯP�4���!͵IÏ ��yAs�Kɂ�ߏ�R��[p�V�d�`' ��E޸�kU5�Ծ��lxFjdwNfY���3��裖�Z�h��rx��XuK��@f#
���-�9���>0M����:L���_�K8̂Q0�_T����������PW����É���@ZR�H�
t4d
�`�ā�'��@NIȑ��icL<^x�V-��.��S�f2�T	�n4�����XBs9E3X���J��D��N��Ϻ���Ч_�+z��4@�;���[��d�^	7|W��VpA�����$<�l�0�ฤ�v:p.�..U=�P.]t���h�����.�vx������Q���=	H�X�HV�~�Ř�Ѽ\+C�;?�F�Mb�<E4c�B/eXؠ�Ĵy�7[a�<XKI �v[|�u:�.��a/O���h�C���6/%ѽ₢��KS<�i �AIB��jT�T�J[�ZZ�h�B�I�q{d��a_��hm�������	�)�1��VL�⽞Z���2��v��_|�Q-��+�v��aΙNw.�ZC`.�B��Q�� `��E�E�In�~��]Y`H�g8�ƘGe�U�Ue�����87�W��n���hl�7a�О��_F�A��Sd�M����r�R%�7��.��� i�7��z����3:5��k�����h=�Y��35��=�&N~32�jP��?
���a_|v�wp)P}�a���:��@�*�8
�$��olw�+Zr�u�@��N8�-����V,g��^V���d��h;#��\_������b�ق�u����*ufz��G-��I�D
�A��n�����CD���_���=�G���,�KmC�!��{������j5�eMx�e
;N�Q{���j��5<*|��2��i��k��s�(�����P��V����2��f�b~҄d�N�
WqF��"�H��U���wuLT��'��~gւ�ܩ�B�!��3�c,L1������� 8�C��E@�%����xn��J�p�O�|����o����y�O=m�˴�A<�d�f���WkR�Vw��#F_�DC���G��AC:�Q�d�݅��~UL,���G�.S��(�/(�%�ë �.�7V:�w5����[�'.�]�J��`������8"�k��Q�<���r��W�]��-k��:ǹ���v#	��[3~{Ӄ�CR��5Xs1#Cx�D/Npl˦�O'y�;����M��έ���X��I�L`��X-w������)�񐙏5�q5ea&�Hȱe_���(�֡��A�@�@��`.�M�w�y�"<�����D�a��Ӗn�H
A���dÑ[kn%*AF��`o�J��o�O�����z�I&�).췭�Ʒ t	��$Tu��c/qGZ�:H� ��`�4������3|����Ő��ŲW��D|���KR%Ux��ƙI~D��)^��d��=�t�}���Z����%�o.h�R{�q:��8a6K�Ǡ_�捊��xhd����;��~E��6�����?�T�[eȪ�gHi��Rp���%�x��HL/�������H/ڇl���Ş����;-/ɵ����/���~j�$#��*���<��RԬh7I0O��51(Y!���
�2��Zf'iu"���ԃ������`%��ߝg��W����z��&�A��{��R�V����R`�3]M�9l�D��<P*p�>�N�K���[ZoWdI��1O����W��&�&���_�2.},�9G����f�?x�Y�,6�n��/Þ���5�Rb������5%=�z����&��҈oX#���a\����1�?���#��{�n�n�^ZU��&�l�'������v}�10[1�`�������#�Aj)r%l�'[��ykJb���ǅdH� +(SUG8A7RR��y�G�S�X��	���ZP'���W�o�!F6�������-m.� \�:��[���R*hx��э!���_�8Y
�`N�h��{bq�N,[�1<���!��cG�j*����C:����)�����ߺT��w?�m�18��]�E����	���F[��pm?*�"�K�!���r�� ���io�t��"��Ow(m�I%1�>¬+$]@��ʸ��L+t,z|�����F�?{�z�-?%c��Px9T�x��Wo������+��jrlx����FT;:�i�o\G4�:�Nr�F��6�ux�+��%�g=:n09�ľ�BW��?�7�9P�V���B��o*{� [Z}X�ߔ��}�
d�Ƌ|�ͦ%���1F�����'�x
�icLL���J�w ��KNf{�|@��9��R�G4��̯{h`f���_盬.&�<t���U�w�N��g/��i��m�f��c�x�	ILц�)W~L '�:s!.��tB��\k>��;�U�G8y{Zb+�9eٜ�b �Cj�p��Ɏ#�B��vJ�K�2�_#H~�+�C��A�4���`���'��Q��qs,�Wj2Zgd�o� ��X����=D�(WF!���D�aB#v�:d��:�\�$���z
��Dƺ�sb������{��~�������P#��߹?���>�#��낤�W�������/d������f�ʡ���r��d���y�^������c-7��xѣB��0� ������ޏ�����2��D&����eն��� H�_�{8Ť�_�8/�h'4y�hz�<Fk���⿲Q����?����A 󐗆<�9��NC6f��3�y�y��X���&��CݏQ2�t�ȟק)�����U���C��vDO�I����g��tI����1�,�{�RnX�5�v�oW%��T_O��~��U?��fl���5�&��6�:w��?�yjo$Ӓw���^J���|=��>u����k�Bs7��܌W8��Q���Y�2��	(,@�f?���	�����4+�;�?�f�)~y�����;��6��f��N�ү[c<S�����3�
�����(i�ԍ#f��(Ù�lR�w�<قCM�,r��><O��lH��F"�xo��0�@����O�XDz4��N�B��.u� ��P]�[n>x����V�3�B2�	��H=z����q�ʏ��W�f�X85��91�s���"j��K*�Ϣ�?*��65�Z�����F�VD�D,)e4���L�=0�&Ί���2k����t8�)<�֓D��w�,S�F1�c�yF�����`@"�{�nXw�?ͧt7OS�03%��ܱL���.2M��J[V6=�S�!�l�<O�e�4Ԓ��~3�w����h	xM���Rg�sj��{��o�� eE�u���DV�#�Fa��in�b��-�Y JZ��tJ���im������rgƛ�%^�vI+K��ɛ�ݏ̃�� �n��%kcz&��.��熜[@{��b5�b'le�
��e*K�� �o�y6�Րnۛ7�붟��ߔ�֙m����z��ާ�igi��)K��d�� ^�-��Y����� ��*�f��et6o߭�҆�rH�ް�����r��A+<��������g��IDX���4��S6�mX�.�ّ-��»�S<�7��F=�$t�v��JϞ܃�������Z���S+[=?�Uu�\��$��.������Qn�N��)u�o����KK�a�iGX*�#���8��b�n����/!���y��Z�R�ta>�ʱ����
d�A��qE���r�����7d�x�/)��P�?���U)O0i��3� ��@R��(�o�N�P˺�A��*=!�7a�HN�
 ��h�m�D�t����^�7�i��=)iE��ױ�]�1�"���]0Ң�?�1���{ܚ&�j}�l�9�M~B�}�A�+�(��HJ�$�op@��Iu�2�dL�0���NH�������ؘ���I�@�Jp˨�Z�Q�s��{G(�C]��5K�Q�kSA�?�s�6��"P�M�̺u�K�<`���2��a��j���y�lB��#�M��$��w��E��}�����q��k��J_�>J3�͓����0��F�L��R�E1�ƻ�S7#��|���� �OY�8�1Sl�Jy�g��Gt׽�Q�Q�M���_J2|�� ��/�j���	���ظ�H��z�kE	J�����E�As�ub�g.� �g@l[�����}>����.��N�
W�x{+'��E�a*��z�o�AA�|��������`ѫ�C29A�(2W̾�̴u�&e���P9S#�m6(�"ğ��O};�FJi��3�o��ڈ�,�5Q��[���ߚkYu�j�P�n���9��r$4'�LWI����P��\i�!�ۊFJ)������4�*l��L!��L��������I6kF�1�?A�w4��3��%�������&�ru���iE9��(;����~6|�M4?��T�~�R,Dt4���F}k�\�֘vn��r�7đ\_�7�xhI�--�f��]l{tZ��b����h��uߟ�1�V�n.�obǮ�0=x�"��
�3�yU����A/W7�<�Bl ���ڋc���
˧�����̋%�^��ׁ��R�"�jX5��39��l��.�V e���ˁ*�u&���O��J�L���b-7G1���A��ў��	YCt�m�?2
sZq=V�B�������	6 �'���4�q��wݞ,js.G���+Y3�3��m�����MPc[d}L���/`��;�r�1��3s���L���S;�,��*��~����K���c\YC?�Trp��t���vf��qTD`=iD��'��kA�@�NJ,B����p�����z�7<ْ�f�h�҅��|/��Ts�����xt����n����?�eW���sl�Q���1����o|�'�+� ��� �����%A�Ͳ�Y�����kVW��i�q�:�0�s�)�#�����>���vl'r�����C����F��sJ��zk�O�G�aBtr\
����c���_�Lٓz;���l�^K��}�\�c4���v���mfc�C>��|:
�6.]�)}�Ë�s�z
����yxˎ7ޮ�%(\Z�<��^��4v�m��'���`4cX�^� ??PyT�!Z=��ܪ��U�$���������	����.�N��QӵJ�(��됦��ǫ���`Kg�� �&酇�@8��d�b3���O��;�����[?�Kr?ʯ�����@3�A�%"�>Xcd�9����t09tSS�n|�E�����`z����EW�=�f�<U�:���i� ��2�a޹x��������:�p�Az�6k���,p� 79��R��O�����>���pm}��k3�;�"G��vY�|�����*��)̊�����t
�ZM\�j�:T> ��)�!�Ns�T�#�SJM~����Ҁ��ŏQ٩�4�G�y�v�C��&J���K��l'׹oK�+B�������S�����t��O��Y!� ��/i�o"��E�L�R���e�m�<6��8�C�xEGs�� �34u�-��n��`��-��� �����U.*S����d�������� �a0>�#w��3I6��*~��0,*?w�_��I��V�ߕ�����x6���Xp���ڗ��z	�9���4'f��˰H�@���ɞ6ʏ��߸X�
']4�.<N~�=,��2���cR�-Q�HB9Wh����3�#ly�k}�-�'��ᣵ�%?�v�-4����+�Vzȝ��AU�%��Õ����S�;}���{�d�*>awrg�����9�l����P���p��e�%��\�n�p�D���ۏE�$�ca��ق+ꐴ:&n;���TW]�x/v���~�����0�E�a�ݘ9ԍ����v7����U��z���Pϓ�
a��a�9�R�!�@�G�;�y.�
��6�(&�.���>9 �Ϋ����DS��.�@"��˴�u�b��RW²(��)�����&me��|��k*���U�HM*�A�(�xaei77	в���9Z/�q�^u�A�u}�[�}:!5NF�Q㵹7�g�
�̱Va�o<����q�XŦI_ m����{�Rs .��9��!��a�z8Ӂ6Ɍr
�����gRp��W{�S?Bf�t���7���2s�rmv>G���T��.S�������r ��7�pv�-����z��i�]'uq�s@U�otm����J�+9��6�(��Z=E��?���"o9��Dt���P����"���l����^m.�Dv� aK�	�4�C��$#��=:zD[ӭ�_Y҄{���;o�}_tܸ�>:Y*�:I���1øʴxSK�Q'%�d^tF��TY��\�d�!4��� �N�A� �j�jU�ld�h�?��x�LPR�T��k�3����45-$���� ��;<�M�dFH�?B��l{��!?����S�t1��
��=DO;�qM��W�#�@�b1	���		�f:�� 0/%��D�-��[�����]���$U���)�e��T2��������Ѹ��� �q\zӁ|���d�����>��W+(XwZ
�[�z�ͅ��͏Qv�:��G���öa�&���JT�$W��k�emX�)��Cŧ��B)�P�{l,,�L����*غ��rH^tYm�G|�-x�n^� �1��O��X��fL�U2:��P����d���e\i�O��{��ų���G|�ki<3 Y���Vה1zQ��8�4��=�e���w�$��?L��F�f��ȝ7�D�"�	���%�!���Rv�������2�k��H<Nj�ʯ%�+a|o��G2�qҝ9�Qfb��@���1h��ZﾖFY�aq�1�
� (��r˯�qH�pN��`�˭3�\Mm&r����{�������JO�Ⱦp��K��L��m���n �Σ�c��*,v-��鶴|Cj��@.Z���**Nh͒�$�bs� �w乛[�d��>���-�jۢp�U����Z�7's�"B�<_�VP,yl�K�p��$�\�g1V"Lf�[���gҀ%<qT�o��.B�M,�x��1�HE21�෉�K��o�(V#4npР��T3~�4�_���tHa�Ui.�nQ҃'�'JϾ������)�0�n#�-mK~HlО���2{`5���X"7.��pN�B��/mN�Mz/rc�� ������	k���4�k�т���|��s��q�ϛ��1�Qo�@��<n�g����=��0��;�?�1�~f�/puњS^kH=�S���p����P�%��:�6o|M��7�q�:GW��ay�N4Q:S�8PW�^)���i2(|u��m7�2Lsc��e�~��Jz��!)v�!�n1�*�ٚ�MH/j��?j?�CYa4�c�P&��������T��d�Ro�Z	��%vwo�?��=���0���aMv�H�<7����`��>����f���vu��(%������H���1l���S���J�5�y��,?.��UM���zkac���X�v���cJ5�=xbQ�)e��:�~��a��Ԡ�*|=�:�o���`RHƙ����K��(����l�h$�h�"���UF�>Vw|�-]\�5�ZA{LIX��2�_X��1�xENT�2ɯ�U͌�|p���<���~h^����g�����G�W�JO���iߌH�g���`�=�b ���,0�6=[��#Z¿A��� ��k�o�q���i�=�+/�\���z���?x<����
$��U��y�~T����%GL퍳h�^�^'��w\�����6�BꂥW�l��44&����V�wp�ow���:��K-�EL�3���l�[G=��4Z�.�g��g?��t�x��Wn`{�vb"�Z�A_ ��K���Ź�<�Z_�0��;��[J���*}��=0kx��4���!Lhz���8��*��� ��}�Y�f��pYM�<����V�dJ������+:g��v�S�M�\�;�1��dt�,��׭z5���B%�� o|ɘ�n�<�o#�_A\�WPdG�{���J�$�h��m�C2�1A�M鈓�uql���`���'�]� kQx)ր[�Py"�wI-�9&S�a��L̚P(bC���Gpb�c�Q+b�]��K_,|M�ӻ��ƞh���Ⱥ�~�_R�^$��as[g~�#'{䏐���� ����P�R�(�Kղ�%4�`�S.P�1D$"�������6�{�G�/�N�:�ٌ���nIPD�@,�a�D��)�I/��pӆ{�1[v�.��df�F]h��Sn��o^�Dy�.���z��Y��h���_s 3��ɯ���a>�!��`n��,l3��� >*Ҁ.ݟJ��|�>��V�6�@�7����_��;2[=F�Hp�Q%ǻ���$�5ߝ8���쑜#й�\�5\���L�
$�c1~��+�A��m.Ӝ�E>����y���mHgj���{'�Y~P�D!�����eڇt.��/bhc�K`)Sq����Y�ܡb�����	i��^�]����K�+��?9@x-�A�"l�R��PY�7
@O�5������"hi�\�d����u���?8^�`�'bY\ۙ�e��x��=�\�b��̈#:7���y�)>�Ɩ/��l�QP'���tg�o/gcP\r:���ܚ�k8��B ��n	@��	����1I"﻾�R��폰4B����J-��9����\�h(/&���S��k)���j�wX���i7��H���E�G4�0��}���/	�������(��݌1�p%������V���<���
&�૗�g�l���V�����F&�#��ƒYa-~��dS@�5�NK�e>y�R�1~�QZ!�T�����Tv�2_�?����<E��xR?�I���&R)�CF uc���6d�u8�}(��US/<�������LY�w�O�R��� ��d
����W���>@_�0��kV���#�At���9x��e�,8U���{g���1_�.IΨsZ��UyMA�B�Ȥ}���+� U1���0�!�氹�N԰% O��S�d�?�3��M���L!cbZ�vO5�3>O�0U�����<��Y�l��ξ���KӸ�qo���4�C�����W6Xm�0�������GF�o#k�`���})<��1y���3x��<8(��Z�-�~sT )�����\�J�J��gLD������.��feJ'S?O1"R��@ur>�	��ր5����)TC��c��TuPIQ��I�qQ	������5	i�˖�z����p�ѷ�p���6�ZY9�o��Q�)�F,�/پ(�amDE��P�ś��c�t��4��u���;}o�9k)e�IU��ٹ�����qE���
cM�&��ŵ6p��hܑ���ہ'�����xo�V�$���}W_�#9�zD} �y����h.���0k稀�/q��[�t"{��
�_��@<��àg�|ڌ�t�U{hk~F�W��l@����z}��+�����1�D�����kfo���N0/#l&�[
MVؽ���c�xcGp�k��xNPjЬk%�y�\��LZm ��i��f�iuCs�7P%H̋����n}�	&�u���g����vy;*4�*;�YYy�L���{��}�uv��.>҇PT/���ۋ媏Q�o���86��_����Ȱ~!@eI)o$�����R��d��)�G��9�q����歾X6���R,޽c��k�9q��@��+���<�1��O�q��t*�⅞{��A=��-0h�ӷHo���XM�Ƶ�{�y퍼�7�D�u{��9yv������<�j��=�S�������р)}u��h1�d�2d�@/�2<;-E���;N�N�]�w�� Ru����.�����L��/�]+�{6'U/%�~�iO�Q��Dj��<����J��.����]F��/�//M�ТW���̪��]K"�;I.�\��Y9�!/�Q�M2g���gR<����z=b���.Ms�A���Q��O��� �r��� "H�dܽ��3�HZ�:�s��?����S�n��/��Y��H���z������<�ȡ9H�,d��j��]1<���Uȑ�? `��5��y���e�f�Vc*��IVb.c'�:�$ $��DHY6B�⦚��j��n'�;��65�+��dub�*�MƧ۳2w��9���	�a�K0W�M�\���&�;�"��D{-�k��P:r����q���`H&��&��a ������-{�Et�����cP:������B?��2�&*x(�>P���ɽ� -�����4�Q'�Y���4��΀��#֡�x !�2����q��=�d�*�۲$��Qq:' 7T�$��v�ͧ��NY$��V�ŭa��?D�qݑ%��ίn9�/wz� ��E�'������)�L'�g5Eu��'��sM��U�M���u�t��k?�k�G���1�<5F������L�K�z�Ά��o�횽�xM�	�� �A�C��͗���p�9չ�z����N��ss����R�/�� ��Չ��T8O������{8�����v��o|\<�2k���䥪q�fb/d���ӳ̪�����&�շέr
�(*Pc�������n�v�
�������ȇۋ�~������w^a�i�o����x5�Òn��V5튻��8�ͳ휝�OV(�*z-�W|�.[zNM�-^��ފV�S�δ,mҦ7�~�W�����2NLM`0ĥ;�d.ۈ
\s��5��=����|���RETsp�W�.��G����>y��[�Xj�ߥ�xM��v�ߺ����3���1^�l^^-(j"p�BP�;�_�OP@�#/@�����������ܒ�ҝ�/�:� ��p��H�Ɉ�D���nh)9���3������Y�D�Ẏ�C?�V�՜؍ل�_���a��ݞ����_W|b�Ǵa�����m���%oX���.�eE���<�w�LF�hq���JZ)Pq�]ڴ����U�[M!3�l��V7�+�J%�����9-⤭zI��(�|�@5[Uƪ*������/}j��~�PP8yM�r���v�LUTo��>x��]��/����`.~-NQ��1�&Gs*,4��y�䚈NB&�G8|���n.�s�P��l`���a.���S<�=ܡ��[�Ƅ������hZ��&sʳ0嵳��hA�x�l� ���dT�4y����S�Uw��+��u���|[��|.�3�B�|v��cc���.c�h�ek��q�,h��(�\��$h�ڞ�X�yk�KC�v;�󃊓�9wß��oI�(;^.9E�e�[�p?�^H�cM�"d 70h�ey�}�]�3�L���^�R�$o�3du�i[��)]���,_ͱc5sUK*�1������d~��-`Ȇ�i2v�lH�C"Ђ7ok���a#)�C��QB�7����>�)������s	��|��e��]�#���oM�3,Dy�ѿ �8��8��n�hxiӧ�ˀm�ռ�3��Z��|t�}3 ���E�LŚh�h���ݾ�p�49� �90{��6���D+v�I��u}1 B�������v!���Y�^!ֿ�����{�qBE7�;s�?�?�/��m%pMi�^:�f���C=�;H�H�c]t�Jv�fQ��n�߹�c��S��e}��F�4&���`xSk44��������J�9ڴp���ͻ4�t���p�6O?������0�H�^_�s���;'�bc���G��N�C�
_�j9H�����+�-?�V���[3R�𑗲��R����>�y7"���T;�5����s_�˕�T��w���(%�6���1�#���Â���ݿ����ڎ{
_���j�;I��������T+!�j=�B�!�H�Ax��Fͻd8pt�T4��3���I�u9�×��x�Bd �!����a~^&�T�5��t�P�as��*>P`&�ސ����������J�@ˤ�o�T�6�T��r*��B�����;�b�X��g.�j�;>9�ݽ�/W���"�% �oer����M���Q�eꄆ��}���|���������p�o (�R� �?Cu�TB�����66I��1"O��1��p)ȫ��m@��*���}:�4�MP�7�=�?���Z�;��{�Ol�ï��r �4���O�_��~�^��̑J�VIV���̵��u�AH����K��[��`X��D����e�6"�>WpHɢ�@�Q���ю�'A�6���r�y�N�I�QS�:�@^y�|�_g#���ejP�;oA��c�w'&:>9*�}P��tm���R�#@�Ȭ�p� ���aun��ʿ��|0�j���~c'�i����~B�l�%�Z���RS���t E���|AZ����'6�A�}�R����(͛� �$����J���m~���vx�)��wg��AXV�����O
܂AO�~ٕ�)���A`R�������	���g��־3��Şgu�x�����=��?�
XGR}\��j�X�L{Y+L�)�]��˲^���^5]�\~aj��t]�L�vnJ����Lt�t5)/��s1���8�𪥫��)���F�� ��g�ί�!�+���8����r�5�3����к�eo�U��p�C�_����iL�X�����wD��L�8�"У�q�bwp��*N-ʬY�g��@5_R9��,11k
�s������I�{��f�g7�b�z܉R-��xU�r�I?�$O�5<N����/�����7�=��a�ٛ�y��h�����H�P9-�g�4�N��;F:[�U��7����8��z���@���:��ҁ��N�~� KU{;�|*���up�[�8���e��c\�S=�^��٤��B��s&r�p��2t�[���Y��ʁ%�v�N�D�Zݡb��Sd#M�Ga�<(��إ`��>��Y5��{��`�*-hϼ9�5��������ɑb�4R�$�F�ѡ��]�b�&T�$:��Z�����N�i"&��c�Q� �dz�)f���6�N K��u���X97Y	�wL5���Dk�b�*�ʃT#݄	�Xxd@i3z����Xb��$�I#ո�QR?F#B�"J������P/����Z��d׌�)+M��9{{�oj�c(P{��en�ͦ�#v#Yd�5���x,�Q�XF��QS��dJ;9����t�պ�ey1�J��أ�4͂Tc�&�	���/x��э��<sN���q_N���̷:lc%RH��e�(�j�jɏV��������l-|�_���
M
�OO4�UlE^;��$@阗�Q�68�k#�����[�N�陊���\�~����Y�z�m���!d��#�����x��H��2��
]��4�n�'xQv�T�������E������ pq��c���l��0�IJ�!�Jz|����_�P�A�^��7Nb�Ȯ�w�V�&D�@Ɋ����k9���DK� �|P�L4u6���5���8�c>�
�f�n?�v�q�r�).��@p?:�fW�Q��6@�Sz�2F��9EN��L��o�=��R������^K���D>s��+�H�dt�S	P�Q�|�.L�JY���Qo�c�Hc�*�Gs��0�.��@)�>R.��]&�@�x���~�O��[n��Պ8 FU1�_�լ�_�i�6�Pɳ�z�i���O_=�WA�u�i���-�8�����bԘ�jD��S���i����f�.�s��v�huz��m��#	����?$���� yՊ�����6^o��vTsi����*��A<-b��b����kꊂs�B�f�E�Lu���:*
:�+�2�0}���%qŽ�[H�ڑ�#���h�&�"�w���л�]�5�		}�!��;Hq�Y+C� �N��g�^�
�EF�����W�'��V���56$6H~�� �~�2�����Q�z��E�T�r��"�Ro�����QM$r�9l/��N�e�Mr�P+WD�"*lߐ�)G��5�-n�6؈!�y�y��i���{�g�j/]Uni��La�V�Ĕ��N/�P��ҧ(��/�Cm�DΌ_�[B�-��S6u�.�_;��0s`��i@���f�a6׃=�u�K6mL3���Z�q锸 �����̡��,�����c����<y�[x��N����c]��M��^h�t� �`߷��fK�)m�=%�n���6��������pH��l���֕fk!6����ZQ>���%�Db%�A����{�i���<��n�#GHS:�!���	�;ܪ[��x��O�:�}���3� �-�E�I8�Z�n�<���;����Ȯ)�7F-��?�uW���w����K�ޔ�D���ǫ�.�8Fi5��Kҕ3�C=���������Q9��}o����-�!o�ICFBY�}�gK~LUX�*�i��u�mR:���Z���#�/�xHAs��8�2��e6+�V?�\ �)l9_4b\��4��(�G\�X���S�$�\�Ia����Bu��x�q�nb�GK%�I 0vӃx.���Az���<����s����_u+�[w�w��i{�b�e�$R�u{[T���;�y�e��A]%�9��*�f
�:<�[�昰!�p�1�HO�Q��tȴ��խѵ�e�
���nN7,;����{T��Pk�& E��Vg��� t�5���JN���O	�1�x�/cjX�,%�2K��o�|���V�^�Ԋ��AA_8zV��.�ި'D7�B�6��}w�9���� I�8֦d�$��m!%�o	�CY��Ŧ&!>����}7���.������B\ǃ��b����v�͊�c�Q��Kh4�c���/T��v;���-/���/uS���|dhn�A��t�_�hM�θÎ�ͣ���P��'fA
���.�4�����a�O�J(G�/2T�6�E$�_T��(1��/,�"�<�
o��Y1	D<�¯��N��	�X�%�r��__�{��6V#�څ���e�|����	���;�0B�i��o7k���m�WiH�D.�/��jz ��l�c�f� �<��࢔�pڱ� �bl�����4�åk�&(��zι-Q���
5���-K#.�V���܌�=f7���4,c���o��4��=����޲ĉ|@�!��.$gHk��[@� u/w+�[t�BaW2(�8
�ΉP��_ţ*�x S�C�n(XBɇ�9�~���c�t��:FBe�NY���t8A�^�y"�~�_$�Ȫm�S���4�b,RZ ɾ�h������-��(��-���B��u֚����%T� (�>]���>>R�[D;y������mA.o=	v�����U�G ˗a�]������ɣ}�+�JzB_e�'��q�Ut��ׅ:=l?��߈#���>�1}*��gi�g�kO�D�$r!W�^�{��0*6�3�ҚO�9����Ƽ�M�<ݸ��0Ef��;^>���'���`t���kʟ���g�L�A���l0�f���.��7T�i�(��$�Z�4���ı�6�"�,aj�"�"��)^a��c�{iA2��GvەL�B��]���@+z6�T���ޚ�R�~��� lz��zӁy\�� �Q�W.9S"�����vi�����El�ԋm؁��]���M��6˟!�_��aC3�$Y^�&��Ž,�h�J}�z���C�B=QUY��8#=v�+*�R�h���3H�k����pU�e�����ʰ�H�vGL`��v9�HE~��O�U�Ke�֘���H���<���T^0����[����es�EE�%�;��S�kbƵ�s�%KW�Z>D��eC	{����� 2��P��^(w��T��Vd��A�(0|ϱ������b@BTf0q.��c����>���i���}3�J����t�&@~�tp�Խ�=z�|�O��ȐaJ�t�e53�b���\�5'�pA��$�����{F��ʨ"S�b5����6g:���B���&N�3�{z�S���\�?���F	���]qj�/A;��^�U�o�$�g\�_Sj���r�p�O���9�+�F�+|��{_ȑB��m��s�F���3�F��E$�Ǹ��7�F�1W	��<�(�Ye���c��M�k��jm��q���ĩ��Ś5Ť�Ώ��I�׌H��$���oDY���g&�ʙ����;�[+�YG�4����5m����M�8(묢���4JQ���]u�,��E���M��~?��L�9"���X)?��֌�͘o�Ǎ?�͇�ju�'�!3M%���!V6�<5b �S�IT,�иQӲ�*��:�ǆ�C!�=�+����&�@�3�оk5�� �D����a��~�@�z���6 �D��*4U�Y�����$vEn�g����)��>���)t|M���~��j���+��K��M}?��o���Ƙ�/�<�-If����T��ŋ�b��+�$����}@U�-���l�����^-�d�q�6�f2MƊF��-"ez��X�<BMY�ߖ�+B�q�͞B����xg��/�̼]D�D�QGV/cOٝ�\�^7�c^�lr6T�uE�T��sE���} �)�S�Ȫ�AR�9��;��!����T�}����_㑙���J<B�R���cˤ���voa��BT?s(�aW�e���O��~�z�7�^��)�ً�L �6^i�+ذ�T�p�q��¦��Hv�mPB���~��>��"�)���T|Gƣ��:��H�W"�Mo�b;���l�Rb�m�����p,pxq������t�v89N?s��-��X�}��W���$_xd��z��F��E}�o$?t���&? }�gY��l��3Ɋd��ֲˍ���DVDP4�{+T��9��p��L� J�Ҭgu�B�|�>w=�blm���w�vU+��t�=+F��O����3#�򨰸��{�Z�Xg�w�j�E�|�<�ކy1��|��h"U�pE'W�8�{��	&��Ӛۗ�]��JR'ҔẄT�n�2�:��w�f�'�47����Ӹ��Ւ>z:g���W�3M-���Ֆ��m��U�{��q�O��b��qK7��Dh7������@��=���v)Nǰ?�%5`Z�zG�{�B�h��h��C
S���rh~�v�ӝ�MuD2L��o�}���!s�o����:��/[r�q(멁fj�ɼ��H'�Y����ͭ�
����v6F��*-��C ��T��Fn��:���=� oR����N��ls��1Wt�uk����2y���G�{.�F ��)�5=� (��ɴv�(��%J-B���rdICԛ�������Ijf	
�����@ń�w�U�U?f���3v}��OC^CS��G��Ȥ��9�<O@��?>>�8��8p-9<����y�&=�1��c�X�[ɦ�z�ͮ����rKf�l���A�{�o�&P���IƆ�b%7�e�p�:�6}���P5��G	�n[[$c���$'L�����0�a?;?63�$u�}�\�\�R��fj*�B��y��lB �.ui�j�>�tEWI��[���Y`����iW��4AZ�4u�t�a�>��c.�E%9NY�XO1�$��G��`�@U�*��-��ז���d�]���J&��)���a�&q�<Nb���3��>@��A|��YDcq����d�!�h��m�������V�}+�w�[l+��j���O��9%@�pfg	�m�����Bl��b�Cؼf�c7ʈ��������`;j�=��8Ȩ�I�w�7N�jk��j�k�dc�*i�P,cpH��_�iɝ��('�e���饈!���C��j�!�*a$!�{�(h�p�K��-z
kq���Ne<�f���.�z�����Ǜq�FE��ļYɒG^��X�	tŐ�w�(����^43r"��8��w{���ز��몐i��_L$��4 �Q�} G��'N*��{����<�+攎�Z#c���ن����\a�ր�;���C�2\���}� ��H��XӘ_��tjq�-o
.˖s����3	Ɇ�k|X�x���ALc�w�zN���:�����=l�q�⻉�5ґg�[�������S'�'���]�ԫ�ؿ͒�~AY�w�ԫ�O��ݍ�7�:K;l:�XDnrY��[ 	�Grk__C��)����͝97� ��ȏY�&�R�zx=��HI@�i���D��4�������r�Q��T��^�j/uy25�_������n����P_��%ࠡ�$�ҍ����_zP�/N��Z!f�;���(0`,�
�ø��|����!���Vu� �������
��gn�DR�Q�k
%54_1�)�òk�q3Ol�p��2�8�"��@��c��|�Eׂ}|ͪ�{�a�k�F�M��o�߸L�Ek�4�Q�}�/b��J1J���IjޒǱt��F��VL��X0nTN*	�ቇ|^p���0���R�=��uB|A!*w�q����7qG�zT����q���X)�S�������1�:����b«�x=t�&���W��r�\�AW�=��mȑ13���44�@B����\����{�h�^"����Q�b��]ɇ��f g����`��C28#�h����j�՛��x�~c�l)Hq��ɴ��` t}�ky
)��Hn�j���	 {t#ˋ���)ps(�9���q��b�˧�:M���!�$��E�}U��p�#�$��	�c=�d����g����Q�V����h�9K���'�1��>`�$=�g]�0r}έ�8it4���\��R�}B��(�x#�����q����=�v�T,9ȃd�̯ �����o��T�H��?�.�!{����DI;@���
����DK�O"��d¥;'`��B'��=0uH}$��K¤���P��`ۖM���iT����U�l����'�Lh����4��O�)ǝ[�h�|�组��>��O���W%����|�$F���2�9/��{��5"�Lx�5����>B>��u�Y�4Tۛ�b��}c���f�9��s�G�M*-��:�
�\�`.7%艢-��y��l-�����o+�q�� 5��Ħ�jฒ��.�����$��%*�g��{���z?[�����(1f�"�"a�mH��<}��/J߃K��	`4���YU��G�dm���v�����ɡ��M�5qg�XO�J%i�a"bN��E�G�����*?�ʶfC��	h�e�HEL|ԏ�N��'E>K��0�)�;؄��6
̘"�UY\���/eܜ©Fw̬]P%��t��f)�,���V�{�=��U����קbd8�j��_�l>!���%�$Ɲ�:�?�*0ѭ�ٙ��D���K����%<�ox���բ*���PCW�7D J�cI��z&�ρ�_��iO� t��'�nT�u����7.�ۼ��^g��;mfIu�3�Ķ��i9r+�B��,���4�������F�Kԡ���ArsÒ���M��ˉ��>���"�!�X퐍����?T5���ٞ�|1����Ꮮ��?�?D)<EQΐ������Hu�5g�Y3D����q�e�UoL�n��S_�I֕)!�vֆ� .h�=��D("���[Jؠ%�HS�|��_H ��0�D:Eٷ��Ks;[D?��tN7Ĳ�������L�ፉ�Z)2��KS�W,�S�Dv������S��MW	�����(���j�Q
űO�:;!���l�G�fT^�~����7�p�c�x�>�'��4��q�{VC�.��"1�Ja*��B]�RM瀈�'�*�����$��� ø��Hcn*�gа������wr5?��.Z�`OM�8�TH� h�p�kb�>nNoZc���d,	�tb�ʘL�{�I7󸲉��M�Zh�Q�؟Z>"V2��F�R�J��0��s쬃hbt1K�>��8�#�wK��rS��m�x��0ϥ��W����	}��\�ʸ�XhJ�~��c�V�����~3��Ӕ�:)���b��M8���to����K�"q~�%�)1��1D"�C�T��PN��6��j ̻��-���S=Zܳ���������U�h�o&awmXɦ�!jTQ?���S��������� D�W����x��0
H3��.�6@�S=mk5�(�/
�+:��\DC����e�_4g���6α�L�r�@9A]r_�3\u6Ŷ΅u�o�>�T�z���PH��cC���@�yY[�$l�ε�&*�[�
�1|��ZM��#<�bMJ�9׼�D�?R"4�����U4X�� �qv{=j4��]Ә�[������)42��X#��wt�t	uY\���˙�뱷�ۛU\(kz�XW�Vq�i��m�5%��D��[��߀�he�ل��K�X0���� �&�p��p��*X�߲[V��ㅆ*�j~~��}�t3���7�U�$H�RF��t\��'d������'�]=��4I��`�U��V�a�VZGh�����`Ӏ/*%׈�<2,��q��j�����K�g#�^�7/�+�oO�>Z7�t��՝8����B�ޚ�:��t�[�n��� �IE+�R��PX����tr2q��ϵ�0Y�r�a�;U�:W	�$e�?��9�n%�&%���ܭ'�9a	j����T)
�V�D�c���P8s�w���k�!����1ȱB(T`x�i�߫�1�_/)�q�~t`_R�ژ��N��3���
�{��qL��X�cx1&�	Z�Ū��R�!V��z�*���;�i "�����m�ϪVqT?�!UC���-,��0	�G��Gm�&��Ԥ2�#�]5�ݓ W��N����G4ÿ���d��Rs�:=�-h�v��}��n����F��aS�w�6��QPk�m����8w�W6J�1>a]wr�K�'�UI�C/i%�6q��Z��5�;lB-k�cU�Ls}��u!����w׳e�go���8�V�C����H���t�zZt�t�6/��r��Í
��#DQ鲠}FDɯ0��0�*��&k�SL��Jy�[�rK�2�ؼ�v�]u�x�5u=<7�<���L��Cs�Z^H�yQ�i��y݄4�x0`�-:P0��0T�˪Fw|Z������C� \�_9o������a��gJR�1�s dtMp�@�8��)���җcȬI�?U�����>	r���*���L�ׁ�]�8�pYU��j��&�)�7iV�=m��a��GP��)��O��.�z	��"	��e���X-C0F)_��?��C��m�P
K�yL��Bn�rʢ��hN�{���¡��j��#��d3�E�=��K�_ �;]���}���_�$�A���#�B�4_�_���)bC���|�D�$���'���b9�?ҊׄT�����]8���C��t񓠣���B��9�	�%���c�(�Cdǚ����
nx¶�7�� ��B�d�DE�X����}2��$����+���f�/��ُ+� ���ME�:���\\ma�¢5�y�<�<�Ha &������bP�X�I��m���BV,��;p3�v�I�|y����'-/Ng�$%x?�}�#����mB���Mi$�n0�*=���C�l-�3[��5�i��1)g>��_����l�E����8iRP[u9,C	
̀F���<�lN��Rn3�f~wo��lkf�Y�H�L��?0�^2Q ��lT�ޣ5F
��AC���!渴 L�d�U�I��9���=�R
V��x�?&�ʿ����ʿ��r�?-���Y�G�K�!��JS�	S�G�x�z�Sd�J���B��[�K�A��B;/��t�]������}6�B�69���)
qd��w�s>F�7�߬�݄#+m!^�Ϸ�K�?m��.b~�c�ͫ`���H$wªX+�kjg4-��W��IL��me�>Zņ�3
�7��s
Y���$�Q����Ж-ZK>�# �$n��WS"*U���·��7�D��S)ჽ��E���a�0ӳ\e��n��5U�ח� ���zr���F�@��1p>��^�B�%X�+f>��{��V]�����ga�O�X�����.��T�2��&�Q|��l���]��>���z�!gP6Wď��J˯MJ��{\*\Q�G���A���Z�֛�i��|*h�k�?�x)���+� �&���&��1�A�"�N[�ڠ��.���Hr{��b:�[4�Sb�]���g}_���@�E��I>���������"�L�i�����0e2�[+Q7 �޹]2��H�'.�n�E���X �#�.��=s������i+�64��� I�2��9\M���h��wl���!7���
ur����6���ʾf��wt&���}r�����7J��Vآ1��T�40]}_cmO�8��ܼ����ARe�����pӢ�*���QB1�y,����Lk�f�hA�0ro7֍��򪜝�Xc��p���{�R*p���x�{��8{�\}o.��|��ԛN�`M��G�SO!��Xd;���Ǒ{���3&m�B��0:o�o���m�J!�^�s2M9�h�l�E��ppl�+���Չ3�43�lwH��<����K��N��BGDǨul	��l�=�p����q�B�
��[!I:}����
����{ͩRl8�,�Z�X=Ҥ+î��8�Ő�#���:a�Hî=�$)H+�8G��>r�s�#~�{������i�?�\��4o^���	��������ۂ�Z�J+t͂�!�h1���
ҒK��4����Pg�#�;�(m-|�aG�I7"�[L+�Q}�1L��xa= [�G�����?�H�&��ʸ7fG٪ͧ��	���j��J��P5:�r�ң���H(��&���V�c��<����6���ȭ�oɋ@��M��/`s<x)�U ���7��CEj�l�4?� W��I��Cؒ)��䬾�7.mb�J�6o��e��\�D��,���9v��]�a#��&/ǆ�׹f�D�'�HH�Gt'm�����	������W�hح!g}��C�؃[�Z��$#�j�^+�Z��$����4l;���t�y���jN�鄇��ӂ,����K��,�!���nC�8��3A�/�/ p���N��;�`�����$�ݨ�vcd,\f��k��\y���^+\��$w�ۻꘌݑ����$$l	d�i|��d�����Z�B,d�3�:V&��vZ cY{�V�R*fCĥ�y �: �5���s��M���o�+Te\¦�/D-���P�^;�چ�
�I�7]$�ECL�A������:�d��]��|�F��ͻ����[��k���B���6t�:m ��A[�Į�=g�7����R�Z�ǔE�hP������F�r���\�<2h�����i���O�N��O~��j�y�@ܯZ,�R׏� �g7��e��3s�lE5%��p�W��[Bu濏�T*�&�p-RFCH�/cܕb��}nbzP����Z#X,cy޶*��tE���x�(7�р)92v^g�YX��zD���|K��-(�)��k
���:�r��F�Fi�� ����c���C'�:������,m���V�����BR�:8��b�T$?�[M���i��x;�9".t���	᡺e����?�:Aٺ�!4���b��I]X��#�V�A�V��jǏb�rTF�ى���Bn@�
q���%8����6=Nb����8X=|��'��n�0b�����{R��
^�����=���_%��T�f�/$Pq�E-��r/�zy�}�CL��H��?K@��A>��_&�����t{��Z8�0�]��q�����ge�R�d�O�m��|d~�8�5��u�Bhju�}�r_�v8δ�F�(�(��LSG��8�r�k.�-߰��[*��}�i܍�&�sm��5�Z޽L5���E�J�F�CF:��I���8�)G�p)����>���o����:�b-�j��4�G���͞����%�[���\w��Cd	qMib�m0���YB�hI�^ȱ'���ʺY�8�� e���%7 �S��
n��Q܃�,�������;)i54�B���9��%�?�IV�H�չ�E��|�1V|H�%:��851����TA�;Z�|��шk���*���#�X�j�`�֬^!��Լ���}s��թ��a���&H���v0hk�z0X*�J�/���� �vWFh ���"0�l�Z��S�m�5�^B��󤁭^��z1N��}�>��=�"�f+T�1-ڑ�2�Z�~eȁpRbʮ���a�঑����h�vԙ�*��j.���'�%f�+nѱ\�����iDr�[,���?��-,g�w�}S��w s�D@TxI���Q��+řYw��:#���$
�����"���GT�tD����f��@x��y< 
��.��p���St����z��>���cͱ���	�
+Ý���̈́@�t�Qɍ?��ZRK�$Z./Z�?mj��Q�Ɉ8!���	M��)�R��s���	*&T�i�03\��?��Ϸ�P��VP��X쑟F�{ yf@�0]s���41`;��X8�ʉy-���B���e[��� =��qpӦ�m���B��}~Lm\<d��
f㩠�:�D��rHѹ�@����%�/�O^0\�DG��p�OF�.P�f��:3���Y�SZ���m~��l�P�A���p���k�s^��J� ��V��~4��x�f�皀�nx��+����.��9�l1T�$W�����(��^�D^%�#����(Ԩ_/U!l1y�:�73� �0�0��ր��\T(l�V�"�
�9�ҚȞs �<��E����D(�v�)ػ!���m����-���Cb��pJ�+|I���M�|xL.�Ek���͘��xh�ɭ ������0;8�<���^>#@�nU�&�"ѳ^�W[��#�';�V̻i�
���8���,fv��</�0��
��R!�����g���Y�xjO؁./��?�}�Ys�# �t��=��ͶH*k�7ι?���%*��T!����7�/��.�We%s%z�
 (�>�ka���(`�W�?��<�ڈ�K�K�}�Tt�d>��Y	6je��?�dD^�~'�9�u�$�WIvc	�~����-pa=#-'�(�1��4�v��m@ 1w���Z�����-�^%��1��0�3�K�T��*����z���ض��ϏM��u�����ϡ�K3��λYE���>vE�$g��;T0�c��+<R�%�L��y,�j�vh��1�m}Bì�k��}J�>P�J�n�v�.7^�S����?�,d����ʨn���k�N6
ō���3�6�V�+3�2��*�1aX��*�[�%��8��O�	��2�}@�q�t�����#uu���s�7��}Weȗ��u����~��lm�����NZ��ն�*狐OD���߮+>����qD� ;R���w�j�L�_����2�q��vQ�WɰƔ��t+ml|������h6��(�{���!Y�:����2�0����h�Q�w��H�b�u�t����y�9��V���$F�\5`�t��0l�R����f)� E
�z���~d�-�KNٍ���$��TI1ίc���#A}GF�ϕY ؾ�@�I�E�Z���)��p��)zW�3��P�A݁yvi���莉����{�I��.HtBߙ����;�=��+|���j9�IB�կ%v���J��^
-W��,#�ѡ������~zEu9�c��չT*ȼ2�C`EC�|V��w��gٌ@E;7�{���(�To��g\c5S���n�Qb��8��Ǒ�;�^��w��;j-��_sg�X3�]�SC��Ʊ����e�U��ZgCR�����Bϫ\6��Qtμ�����%P��iT~
���Ɵ�+CN2�M<�L�=Q�_}+I��ĉl���|:&+�iIv��#��b₸ۑ8�J�fw�΍~�'����8�(��0C�n��[4������L�|M�6�H��=#�5�_q�\�S�7�;J �l�M��7�[8G����'c���M��"A 8�R�������ճex�)�w�8�';�4���8{ �8_FS~A?EJ��m_N;��!�I?_�����]iB�!�@�r� %�J;&O���t��K���j��ϧ����*H�6ݼ-+Ws&y$���������`{���J�>֔�(��I���~3���@�W7����mV�I�`��H>SHb�yn^(/߾b(*���)9n{���
��[�2a�[˃�>/\}����$g�6L<{q�'���4�nG�;��2-[�>��l,�30�a�e��6Q�E��Yw67�t�7�� wk�$�S��BhWp�S�T#]Ƅ�VJo�C6�J*�Y�<�WO��W	򪂍]��I��a��8Z�����K�$���Zx(ߜ2tAs�t�xw�#�J���Ð�?3�[����S��+�j�O|!�߶���^������	$��r��T Pl��%�i9�a��Z'yW��v�������6�W�j�)e����P��ؗ����{�?�m����aə2���%�D��)s�&��[��,�
���XZ�;�[ޛ�#g"A=��)m��"���bA$H��G���!��jg����ap�碿QDt6�|X�焖�u1C	��E6�lc�%n<aۦP��`�/"=����^,�����Xi߷��.{r�
��`OtD�^���M�+�Hm!��兹 l� �N|Ȕ��.���Ey�u�f��E2����R� ���ρ��ug^��������x��^Ī� ��U����:[eY,�6�zT�4���"JU��	H�y��۫.��ʆ����!T[�ذ&c4����1O����K�Ț_��+��J��4@�+ɸ"[��H�\ǯ�wn�m�b=�C�}G��x��^���>Z�yQB|�/F��s�#?K�0�f�d0��/g�&�C��^N�.;a�.C�(��'hh>���}�w��H�&L������,�ˆ��B�6�PW�|�&;�������xFU��1KV"g����Ih�)�?_�b`���j����EY}l$&��Yb���E3|��t���A@_�o��a��6"��/+QSx���y?�ѫ���x�;I���Z���
g�����\@�E�-^�{Nz�܍�/�K�Ì��Nad�*Un`3\�޲B>��h9��{+4�h�]�f��Ό��ӛ�b,�˲�.H�z8e�%$�%t�
���n��7��{��9��q�����xXT^&��Z�}��
��~��u%}�"�*���VY����Om�wf�m�/��θ��g�~̙�n��&���#`�i�2@X"�����]%JP�n#���Yəg3ֲ���Fh�4�M���m��\���a���Eg���rݓ�
eS�l֧ O�M�2��`��`Uy{�x��zSJ<i�]���k���`���;�e���P4����w)���X7�u���ei�F�m[(:��./e@�sa����S��� �s�H� ��<C�e�	���2}�N��`�7�����Vg�=�!��RD�y�( �޽�K���s��x� ��C�h�G�n��;���:��5E�؛"C;���1��??���- �ܚ�@�W�Eo�IS��� ����Ҟ�I�e#ҷ?��������6�Y�.JX��8�^����J�m F��#��2�\Eo�^���j}vz�t���	 �vc(�j��UY�\o�+���>dD�$ޢ�e�sq*dR�Ȱ��i)�e-Cuĵ3��ʐQ�Ҷ��-ǧe�8�݆OJ����4{/'.�:
=4/6�0�����ɔ�!O��yn�iB_�hSg*�qʑ5K%~����� }���s��xy*���q�us�ՙ\	�~�[�60��nR���^V�n��WWʦN���cԣ#&�� ����q��>'��dA���'�Y�ߡy�B'����������𺴯�RZ�Q���O!�j'�r��_�����������{e��~qt��lU�A��S��?�Q�}���`�� ���4�<�ȳ����tdt�<-W�:���-L�P��F��B�T݊j���`�a��7�y�mj��3����pi�Oy�b0�\=�9p�X�G������=?[����)�,��Hr⹕�����Q���J�h�%�J̴7�C�T%=%����-nK���@xb���;)�z��Ӧ��74T4���{��m��".�޼
uG�z�Z],o��ug��;J�V��[:W��?e�S,~��I��F`���������"{��8w����Ο���U��P�`��I�7�ئ��d���T��'m�\j��x����#��w�{�#�)*S��ф\a�8f��{�ݼs@��Ob�a�e��	�)�b�\=�X�o#T7�>O[2!`�9L�CE�/�NJ2���xl憚`/��GQ��/�eAw����h^|��Xg\#OiU����_�fI���*�DV`�$��UY��P�pً��y�x���&��:�j��k�s� �,�%�����*)�rP��b-jv�! 92������7���skh�	�,�ľA�Ɂl�y�ڟ�{�Z���il��e�ﲘ������U��&K4S,����l��S��� �@����ՙz� 4�D[��wj��9��u0�1Ŀ�����PnǖI�X.�5��?�e.�-]M�[c�m��'<�]5�*����[�@4��Y)�@I�Q�8�Ńl�A���UZ�'�K7Hɏ@�qH�UO�Ό�$�)I��u��Vs��ˏ��:����V�?|M���l"��<���Hp����A�ۅ>�h��P!�����ۮB�mK�>ۡ�N�Tu��%7������4a#ڷߔAH�v�]K ӕc��������D(�w���˗��-d9���~.-��<,r�7��3����y\���۠$Q�N�E�O�]��F
��	��?�}��Ag�$���4��X�ml����sW�ِϽ!�(�t��R.���u{+�:����h�ހ� ~�r��
�@g�?5�0�v�T/wOVɜ� ̏�ָo���R�-02/>�L�-J�3���;?������$ ���޾����E�{�Vq�*IN����<��������Q�����Q��L<���($t/����,�
�i����*jI�w�՗����������?��t��ԔW������ł8������m%��.v�u��mNeZ=��*Z}�Kt�
���7��)n�b�*&>��6{�&;g;�Ą�M�0�ް^S��}���؍��k#\ >~���T#޽d�� ����BH64[	��M�R�\�-�j�,;'D��[�1��J���
�FvK6�v��cehp���o%��+]�s<<�t-�ԫ�0�<��;�t��d̓�n����Q�h"A�_�g��H}��ZOfo�d�R6�͚�R��Y��I�(�pU�Ϳ^��E��@~��0C�o�B�i�Y�x�
-@�ݧ��Z]V�[��������:����[��&��~�z�eǑr`;���>o�1	���B*�m�:�):lA\	�qu�?�3�5���G��������/�)pЈq埔�����L�'�3oE�NU?�'�c�R�)��"	�71	��i&L˦�N-������,�s�W�+�W��k+�ʘ��|��&_����6z�ٙ �N�j�����k��E
z�f�Gⷈ2��e�d�Sw@��:�.9:7�,H-�����5��ϴV�=)rGvy�'����zsC�4d��^,�#+p{ps#��������<DJ_�'��[s�{��vG2���Bϒ;�I����}�@
�v�+:YRQ���uL�;)��a��x�L�L�qb��sxQJ5�Q�:�z�3�A�L��$�΀'�+�Z��Ԑ	-o�-',�^]#StkKGl��ws:^�p���w��~8�[��Cqo=7,D�t�2T�Y�p�_4?��]�U�3}T�C{�z�I_o&��G�5�(��8�T�O$_���~g�]�UY�e��SĊ}]0�O�M{�f�4��eb�)n�[�s�w	��p\�K�.�����"�'=��9�)��}+��}�C$�(bY�ŏi��W2�*p��� ��!I�������D�$�㈈���wE�V܈F�<�w0`\GC$�A�vª������2k��?6���@�[�)�������]�������D<ʦ��@e�B���
�!!caaVsr�E��j�-�dߠ�[�����Jk�?��I-�(�W��Ʒ��X�H�?wR"x�O��J����tZ���!�PI=���o���p1�zd<����?�
Pha1�Ld��=�N�kȉ<9 s4�<c
����7�����(�Y@ͤ�ww��T�q�6��-2oS�I��J��|�萛A��!	��,������7
�c��9�PJ�U����s����IR����2�T�]#r:���*�N\wG�Lb^NK��M��2NT��:�<Pq���]�G����&��%���>d폴?�=��Mk�������p�y��7Z����| 	��dv꯼���!T�}d�G-�	�����n˶���|��κ����[�4���v�sGXsB�R�����Ѵ	}�F`QD2��^/#iS��sR8�q{j��T��&\� R�V�R��7�j�s�<�������n���.p�[0�w댤u�/�`,���x�2Wެ(YSA��+r��1]{�����PI처vG	�j�"���f<xړ�y}�yV�?�ym�E�5p�K�=�4�Y3���{w��7�Z����q\*��G؛�M;W� ��O�!C����`�]�gj���
z��o�����h� t�|�'�� l�L([+۴;��BK4� èfpu�MF]�� ڽ���ĘT���P����X"��G|.�H�=�h�N���� �uV�q�{�Ͳb�V D$�7�3�jӊ��Y�lR�M�F�� ��g��p���H%Z���.y�y*/�/K�����	���i��x:�V��s�]r4�C��&�j�^�`�;�0�՞�@F��%�4�ZQ:���r㲛X�$w��q?��?�c�KO^)v�xW�p��Ӡ[(��|��g����=�����-���w"�V᪬`�TW�ܲ�#���wf������x�l2�CQ�`�'m�����<`����	ͻk�� C�S���s3O"�E�n2��r7ǲ-!��zqW&�vd����Dر�[�%���r��o�*��h�5�f��b`���?}�$O�2Z=��qye~�-I{o��ej��1ƍ�΁b��������FեH���I#YĴ&O]y��둎jܻ���2�ù�|e��èn�fV�e��i����.�����x�Ϙ��#�A�ΰ� ��H�'��ڛ�盶m2��T�Y��n�C��[�B�euz��P����ѫ�n7WsW��3���8�?�&J��N�!#6��	4���T��7DI���&6u-m(������%���N�����ڳ,�l�s	�C��]����k�!g����~�p�
x
	�$��]Rtt8��螑��|C�>og��q<��O�N�j�!�ym�଍����R&�,�z���I9C���1��XgB��c�-5ę�>��PbrΙ/��ܶ�>��z 6�o�C`�r\�.�C�)�	�fy���W��t�O�)�K���"V%�,�E�e�T��V�8b;I!�As\"F.��N�wX�ZM��^n��$Y��CX .6z��Z�^�D��۞��nc�������B�<�<������΃�N�$�U7^�<ˤ�H������"�WG-eDB�#տ�X'�z��skt����0*�^I��zO������o	�eYm+Yd�F�e�������c2�Jml��E���Њ�c���C��)�`G5���eC�3ٰ��k�����ч�E^��b"o�����|�(��{;~��,3|�U�(�;5��ΜZQ}��.#J�Q1�|�[�7�q��~0��$ߌKE#._$�c��X�TRj?>z����-ɜ�V�5��	�k�YPrX��绞�#ia�х��i5(�}�Wmч��H\DS#�����]Eg�/���{_RZ34��bEH��/׸�oOv������_��5d�5�d��M��Q�k��_�Z���f�+�� �=9�6�����t�����l�Q����A��.���:�m�}�+?,��>x�按�z�V�j� n(��m�@eq�K>����9��7j\�4Z����O+�ػ�S����2�i�r��T��9�%b�O�a�h.��]�ȓ� 2^�b�Q<� G�tV:h�2��7��,�ԧ�����q2Z�|��u/���9��Ќ�O
�d���(ܾ��Ȱ}�(�zx����cM����2"֯��� �O@�~����_��TSR|�Of���r�����\DK;P�ř!�l�1]�Ic	�M�<���_��  E^X�I����c&x�y��I�_��_ t�Fң���+>�ɮ��렙���I qL��Bu��*����$����	7���hkm�/��:���w1Ps��Y�,�����v{v���
YK�����BM{�Έw�Ǜ3Ց����E�#�V~�}�\��/`���ɛE��Ò��6�-��<���b��_���L�R�<�Z�u�n�~�HF|J�n�T�� ���z��IFu��;HZ������̀m���O*�W�R���$�.L-�f�-�is��C�yp�̘��0Շ���*l1dÑn:�7A\��}5?��H꼷���M�y6���X����S7���:��Z� �m����W/��l/���B¡<�JU�4n�f�J�	�caG�Iw+��y����<���RY��R���+����_īG�b��9��(��U�"q��~���%l]��K���Y]V�1��8����iF�Φ��:*|���}����˪���_x�����%���Lea*����P���(���#!;Vhn�uCȸlu�.I^Wemb�B̋Xd�kײq�Ү1/�j�?��[iW��q��հ�ǐ{�)�=�c� "��TV&Z
23���B�p��ה횫����Ac�:��:OН�]���	R����m���vHX��f�ܣ���q�p-ݖ�LZJ�i��*��m,��g��Ľ+gy)�.�(~t���xђ��7*��)�H���^�k-��;�4H��]j�9�0ބ7��q1U�+w�(-w�5��ݽ.#���-��7�� �=T���4�B<���������7@�Y�V[�3�*K	���eI��t�Kj��:��[;�d�^z�%o�m�<j��yz��8x�;�bD�C��~y0j�`-N���2�S�G�����سa�JC\'4���)�e���B朓��C�k�ss���V�5�V�Ԕ���e��o+*��>9|��:kL�<Eg�[ᚉ��#��s	+�$������RHd�G��IG��ʷq�k�M�d�z�Ǌ����'3o�h�?O �V�x:��c)Z7qZ�J��_�A N&5SH�M@��1	�sX����I~�$>�� ��Ⱥ�_d�7&��=����Ϳ���
	��o#�%L���5��0�r{P������\�1����b�Ng��٠�C=�0�dxy��蟐��ّ�f�\����[X�r�� +�z�9��n��䌭3�
���zV2~��/��+o�dʻ2nBZſ5������rI���� 
r(6�E����.H�Ғ9�µJ��ʓ���ZV��0v�b�jc!����������0��-������X�L��MH���y:";�����{4GJh$�f.���d���a�ҚT�B�j��X}�ؼ�'j O
�Sй��B����D��t2 �Q"��І	@�BT ׉\^��2	�֥;� ������Vܺ���$-�#]�@�9]N"�a8�����ɒ�ղ�8�n��E��=m�b֞�dyKX|��es����D�ݶs�@Bـ$��w��,�8��� ��4��)����7���Uu�;=�zt�����U�G�� �K/�=x؝9d8(��t�(�O�%�
f�.�8�Ŭ�tg�����Yl`�LMH�<|� #��-9g�mԀ!Z%ȩ��ή⡦p'�2�1M�1I�hw��w�ܮV�B��\ ;�5�����X�=��j�z@L��G��`
�\��9�.e~:*�gک���5�φ�~cp��Ջ�}���S����J�C��T@,�;�Úo����Br�x�U�De�4����'��v,{����g��^Q�������t��9�'��hn�����V�ƛ�5�
8��4|�
�v�}��%r�Q!נVuG��#�XE4�A�9�P�M����(��)d�k�w|_D���H�n�1�Yw��A�F�
��: ������!�8�e��罄��y�L����Fqf8��Km����{u=ԽIqzx����t�֠oЦ�ex��K�דY�H�0jJ����CK�v[�9�Z�7��9�����HMK�1�u���^m��r�`��g\�9����\��@
���}�*�`
m���o�tK'����3]�c���W������r����ag��ip�Bڊ+/�	�-�iҸ�� ��%5�\��J��u��}[)��#�u����!�{����Y�0rK�;D�:^���D�*�e����3��:�;7to+�]��m�N%NUW��-��n��x Β��Bg9��ہ��O	��B�y��5�Dl՛ax�#j�g�L�"�S�����Dy�,S�4�� ���e��	����4m9 1P�ȿo�#[[i�gZ1	˯{�'H]\�0��%L}�+vT�Z4�V���D]1Օ�u��T*�a~��������t�Eʢ�sr��&J�>�HA�͊�f�.���а�wG�,F� �.��12)֯�%9�,���>Ka[��p���އla��ʠ�o'��g�	Tp��GK��u���w�|4���+�T��pt"��ˊ�1�'��q��G7�
���#�`��)β���1mf �o�$X���P�1��~�.�8A˘����J�Ww*��7y�Ҵ�n=D\�u�"Ɠf�0I�-5��S��Ջ�ʄ��t0#��)��Qח>��X��~��R����RO~K�EK�HTP��i�!��@��4�zr&���3��'p�7��7ݕ5;�����UM7G��(�C���s�;�M�T�]�#vW0��3
*��1�&��L`���'$�;�
O�T���3H?F ԉ~"aU�
Z�	��\�ƕ5���U�������lj���z�	�ǆEQ��D1��f��&-D�O�j4yo>eb�ib��dx�b[6G�mN ��D�����>(E6�n���Cڋ��88eC�EZ�s%��yR�C�Q;�@=$�UyE��صӨ 8ֽ��;Zx�6-��{s��oFk��M�<�LL�����i-�I��e:�B��x."ʔ��40�)�	���"�Fp���0��V���d�������LWN��z��A22:��k6�m=O��Ł��2g-��m��=��&�M��T�.��p�9���>��:mz=�������t�m�^�F p+W/�)Z9ś$�0��������;�h�����D�W�"b	c����7ߴ}p�px$�FaB�ي�n�S��~�t���,`o<yF���Bc�*Y�����ÂS�����=[ݐ���
ӱe��kW��H��⣁��ּ^�P�^������]W�]��M����둱�{���M�T˃����x1�W��bF�!m���5��Mz�pʢUz��k��Wױ���T՜Mk���R��`�i&F�tH�˵�8��s�����R�3cr���c�N��G�G�&��%�T3� ��L�G��!@�O�O��4�����K7T����Y�L\�{�Wc+T�a@���7Ւ��� ߫��l�֑_�1�bT�f�]�.�<R����Kt�Hk3,�9� ��S�(K.�z�R�i�3:����@ÿK���Dv������1F��i4
ϑxKq'�+Zd x9�����hn8�$����_��|��@՟�D��Q��Vaߎw����}�����n��\m=[��Ԟ��z���i�(�(5�l{�ɞ�����g�£�������?S�#����r�9)iWb\��VO6�,N�����r�"��G9*�*6+(������P�jH��.��9�}��Ι�!��O"��;߶(�/���9º�D��?+�*��s�д<��4�g��v���@��QU3���Ug�k�K�C, x�n� 7��f$9@�<k{�J�&et,�¸��a�[y�C{]��*b����v��,��m)'�Q�K2Kh����yLq|��so�mj�ۛ�/�-��`�J'K �V�ގ�><�e$9��M7��԰@t��]ַ�L�8���D�?EB��sĸ�i�B��ᵖ��P���.sl��	s��� ���j�?Dv���Ι��j����T�1V�a����3o���W��$4�Wi/��҈&߾�5�+B��=��4��
�Uox/#�����JP�)�FO�|f.�s��
�̋[����	b��ӵSW0%�x���-�����/1�`%���,�
|�	44�6�l���LK��^��S��+�5˧��:*y6Q#��X�%忉}��e�mji��~G�Pz�^�[�i��U�/)��g��R��q�V�vm����R"b=N��5�8tR`z�����=8�`t	���}˵��D
q�NL���_��3�r}UZ;���������@�*���h����!s�B��a��!�	�����a�J	�� ���{	4UU���F����*��I��-rA��{HU�,r>pZ����]�?�͉>���Bر\�Sx��#Њ��_h����6'� ����qK��'�>}qc'���9�%���#>Ϧ�
�Sq��~�����qb��d�v��Ng\�H!ت�sX'5���ڥ5���;�*�6���m'��>������B\tH$�eĨ`��H�5涕�Q�Um�l=^`����^�#7�C���lٻ���l�G�0apwCԜ������C�K|�������6�|�]d����὾q�������+��4�b�� ���)��M�ĩ�շz�������?�E��U�ƺ�%K��?V���>U0rc�W����	
�������t�M;
uM�����ښ-z(»��Ri?�}�f���m�%��t��ois5�h<��Ь�:J�ǭ�\�>�ިd0�6��lqQ�vg�jJp���LV�B3ʨm
U���ԈBT�3�nM���×�2����w��p@hb�[�a���ػ�v�er�Цy��K���xe��l��$�<5��_ň�AR�;��"�pB��X&���,���Z�fF(<��Q���Swf�6^*\�=g�s�Q�x�٘%��8#Scݫ�*D�uZ�M0K���ɓI%H�.~�&�V�N�I
0)~�C2U8���C���
�-�9�.���h�A��Pr`Gt��q؅X;�dv�������۱+O�3a�V@�]�iU��󯦁<�|�5��(�__����w��^�Pz��ᙗ͏�5�C1�N�E>�y+��(����x/��"`����������M�dTSq)�SNP�s�r4%�ȩ�@C��hI���Y}n˞_������q��PO������12~mg��{�O.�ĥ$�lT
�~s٫�/0��(��a������/)�*���1�Ʋ񕣕j ���8���鎏5�
�ċoB���ŋ���0��*X.t��E�{�#����*�)ִ�F[� ȇ�n�����������Y��jv�J41U�vuC�40br����83�\��+�÷�Vy%�Ľu����4�?�2�u��D��ʲ�u4֊��US�#�J,"�/���E<p�+�~놮��F$Xz�Ԭj�6b��Y�1;�-�b�-cv�J�Z%i�"Y���O$$<K��@S��	G�8kDx$��י*�@z�!��m���-&K-��0�E,�L\)C7RlJ��kBӪk�;�S����m>'���2�$FD��Pi��5R���`j��P�0����t�#�y$�Ӻ"3;���U�C  W�s��{����{�䌉O(@7��6�Lc��?*�tㅣBF���Y�i�L���q�;mb��媊 x��Z�ɋ �q?��;J��3Q{�=����6���C͘���u�5�/���1��=w ��!a�Ϊu��˚�JN�ߵ�v���O�tS�^����̊�%f�o��7��{UU�*�c�ܤ����Q�G��Y��$��+��A�Z��������*�RE+�a���b/�\��qL>oO�@��x�&|�����ڷ/h�޾C��hj&����3^�Rs$�>��g�G1��T:�h<V���'�r����#��N��q�T��"I��ڴN�'z�	
�-���&s���AkɁ���G��J
�2���{[�L���M1�V�S�k���ʲ���{+Ji��<V�~��?��x�O:����3?-k�������_˃z�K.���*Ɋٸy�ҏ�b��j��a���ŋ#��og�nڧi�XzG}�n����3N���5S#^�)�Ķ9V���j���T�ht�P�,����P���#I����Y2��!K��>��]�GH�/�v���ߜk���Rc<d_떍��d��U�b�J[��1�#饥��D��P8��j���� ��B��Gdj�$߲��}$�lX�0���jΊ���e倳-�P�Y1�oL����ں&#�xS��l?� �	�`Ƽ�7�޴	1`5H�b>�o�2J����_S���w/�]�a[�/aC�܃�Ϳva��U�Q�C�c����<o�^�}8��m7��É]"WY3���Q�����q[~B��ծ���ݜ|=ޚ i���4��Q��ǲ�5�w׸�a)�C�D)��Z!4���2�� �L�K�^��'IuR�ޜhN�u~�XjOܞ�}A��K�N�$�
m\1�%��4������	��~G���"�y�g Z��{/i09;�(|��m5��z���С�V>��S������="�)���N¥ ������a��E[]3�2C�������}�?��d�������p�Tz��3��GB'�(X6k��yp���� ��?� �ϱ�ЭĂ�yHǡ��*��s�t�-���`'\:�=�X*�5��'��zk��.(��v�b�!�=2OnwM�>�W��*�t����}��YT�fGT���;�� &�S�h6�;e�}L�nJBC2^\K`?�l�iY�إ=�p��r�Ĺ��Bt3"�4��q�#��Y�U��!d��E��
f�ϟb�@�;A�2�ʺ��`��	z/9h�͒�Z/C����Ap(l�aT0�(�4� �� �p[h%�Z�umD���p�3�\*�a��枷���M]��i�����u����2�eUO�lO�9��k��z�5�_i,�E��:U�n��0��:}&jB���)���#q�sL��l��CL+U%�����a�4(s��k'��h��}b[M���ݮĢ��R���� 4*�B�q-����1f��7
ܜĔ�M �C(�^!��:Z��Fy3H Y���ڱ+��5��E���l�(î^�&�䣕��Ț.�fhyo��N�\����p!Zѡ( 
?-��Tv&��󋬟c!��>T�ۃ� �{��*,ϐ�_���-���^�J�]��;"�d/;2���;��]�A@�I��z��؉�k�#;fz�Q��4��𠶚�o�NKO8���"�[������e��"����e� �d]���"�X��E��ܰ���r��I�H%�I�@��o^�[�G�ƃa�ѵ�2��zw�f��*T�_;aJ�410���S���(e(�_�C,���Сb�l�ȳ�P�PxMr������U�7��)�i#=���o` ��A�(Q��d�n�&t�9S��n���J�L�=�֕����)5!�gz���~c�S�U��|y��#��\=;iAO�������zk��1�����IK�_'���]��9���$;(Q'��Q��L�K��� �x��?����C�9�z�Yy�m����)��BT5��@��^�&����y0�_���4p���ؖQ@|f���ȶr���3��R�߬'ɴ�
(�0m�w���m�?���봀6����D>��y�3��0
\gb�[�j-ٝ1̀�;�n�?��F8AG����1�m�s����3׿h��N�!������Z�]�Oa�#�x*�s�r�1�b	�g���'���aZ����l|4E����F��I�߯� ��}����
 �WRW�1�Y�����]�����&��#���N�To�!�3��^pxh���F,��P8�
k�f�~J����:�� �q��cYr��z�%�,Eopj;6��Ţ�V�;���T���H1W�Cʿ� ʖ8���������{������\\�<iUj(�~��LmZS����~�[±Ϳ[�Ve-ܸ`�Q�A/K5p�=���}���v ��L��̊I��P]K���V�P���@Jw��EW�8��e�R�=��~�v�SD�t"鵆FI�]N�b����#p��Z�;�Ov��K;NS�t�m�c�jR�ʃ�?x�ao������mn��1%����\�fl�~\WHN�6��>�I�.!�������{����;���/���� �\�YUn�F uf'(�@Ǣ�4�����T�.a�Z���sэ1W�����22K�:�:>�`07�Χ����DY$�*�N���w�Ϣ�h�bW"�Ū<ks�#��s���/k!��� �d+;@��7y�D�e����9��uR��h]/g0p�,}K�����ộ�R�f�����3#x:-6!=�sL~K��+�R?�͏{8\�� ����L��H�����x$nX�끾qhF��so�
2��E*-iBT,�Xh�F̒�sȎv�/����6�ޒ���siƘ�r���k]o�mڶ��n���r��ѹU���U��Γ��H�*�Nŗ��M�,<K�a;~)���!2��5M�"DB�@+ M0�W{��r�zHjG`����5�y��(�6����R]�
����0N���ބ�w����?x��I�r��_b .���3���p�6�������v#�� 	#c��y��%�R�wQ���V�u��|�\L��x|�M��(�{�2{�g��#ʯ���2ߔ��.^2S��n]��g��C,Hp�s�\:S�L�g��3�1��;d��(�� �o���\���]��g�K��fo�r1�M���H5���p=ʾx��簋-�9y�b��''T)(�j��+�i!����L��WFVx�!;�M B��ޮ�q���K<����&��{��t����D���{�XS�0r 	C��QEB_у�̥M�Yf�*ŵ|B��~=�k�Ҽ�M)$�jE'i����h}�!�A:�Lp!�/>L��jе�����v�n�IDCE��^�̌�o!��^
<��޸Ĺ�b��'�+��X@`��D��ڊ}�?4�O+�g-����Cv�j�F��g��Ժ��-��a� �BC{���k
��L`�C�~�b�ɳ *S��U3W�)�� ���/bZ�(Z_|lp��`0����%-l����8CD�`m�\��
�� :����
���vvϑ&�e[��td�v����p5,bj�ČK|_uH[�á���ʩ���K+	�\����u����G0
o�(z��R^́ū:B��S�M���"��F�MC�畡���'i`0��FLU��N���	������Y�O5l`u����hH���a'v��#�9ר���V�0�ލކ-�����6&��<B�ʰ���������<`���b����i�x�uN�B!�[�	�X���4>ֵA+S�z�<X�,�J]Y6����l��1��~&(R17R5-a���D�ղ��#���o݋�Aa�y�g�QE����t��H��"}�4ݤ<�`篆���U��<V�+�}Y̵�V�i;
peދ�6^�0{�`á��]js����*�G6y��a]�MH�{�f'�|�x��%=�:xr�"�0�=2֏�7/i����-{�8���?��ެm*�Y.��W�k5=3�B��Ý�ϖ�3c%��wֵ�s����?��S�������6�9�U��#�}�g�o��E�SB?��ͳ�� _���	�K�W���ic���(
 ���3 D1R�k���%��w�M��k�[�I�ܗǭxF�ܧ�f=��'ٮ�2�����`�T���?��WJ٥4AZ��=�S�Z���7�Tol��vi�f�V�x&�7`"�Œ���7ȿ$��r[��	�'����TG�_[)�0���W�9�g|�;�h���?r��H}�E�p���p��z�3e  A.��Q�>ie����wK�DE
]��A��KAN!a݋����jHn���o:͊+ر��;~��l�6