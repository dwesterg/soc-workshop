��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘ��g�x�Ў�+g�@(L�=�еp?j��ބB���{L���X7��o">W��D�d6T�0��:�X-�TxE���$���Q]߸����;���Az˨="��_ٹ?�&֪��;�*u��},3/>W����6J�ngn$X3oC��[�!0g�@��)|�y�7��ϯvf:���?lG��3�Bb���̓� �j+΍J�G���!��aO�l�;b�����Ϻ�r[|3h�q��_}���˗�x��l�!��tRD`h�W�����sR.�zO�Lc�U��*��4��#A֥�/��(��NT�!��ǣ�x���QN�=���$C�-�]��.�Q��<)'��2��
���T����4��\�@�'Z��Tr
��i�7?@�U]6�G���P�*'�VM}Q?w���B#�=/#��DǍl�fV��-��nc\���۳��+�������<�	;|{��^�<�k�B a����B��h�ks��*o�ˤBp�e <9�� �)Z��e�Fm���h����c���Ҕvet���O�Q���U5�8�쐕��a�Ni�&�!<���j@�� ٮ��5��s맴���!1�N�e�?z�,�
  `��G0�YT[���J�U�,�M鸻�os�qI���e�#⌎h�Q񏠳vpQ%��S`�ӒL[�0�:Q�(+U�AD�k�	�ӽ�W�NH�P���e�y�,G�!��bsD;�{wБ��x���Ԓ��!�=X�B���OrI��bg^7��	^���<���VJVcn�@FW�%zĺZ�W��ƀޣ?��VT9���"۫¬���1,��?p:�[4d:���6��N١&1��9Iĵ��	�A)�7Ii��GM���l�2�)�[Զ�8x�	��z���t|�A��	�/x'��Ӿ�p0�%�Me(:e�@�D�P�Gɉ�̍��c��Պ��^��ω��G;�?1|8vP���[�B|��3K��҄���$���K�5�%�Έ��	�J�uf�����Y�j�m����Gl��Y'd���Q����q"$+�W���
a�縼�=BH�7������}g�����0+��x�>�).ES����ܳ-d�M�έ4m2��s"/r��WL�R�{pD�,�'���>j*!4�h��E
�Z��-6����&�����|�R�UW��M����}�P:a�}I5�T912�.o}oM%9	h�u��NXG�Z+�6�#bI;Ӯ��dRs^��.v��jŀ�Q�i�yưt�O/��dI��Lr�b���`Ձ�DgF�Di�������6C���!���/ӌ��y�C��D�r�|/>�Y	��-�R��z@��#}�߿�&�BX�:�
�M>����z�1~�"R�֮�d�I���M��1ګ��R+����Sr"
N5�"�3}J�k��T��aw��ߤ�����I&�BH���
I�"����
��f
O0wn5��������-��%5*�]��ˈG#1$��d[^o�LF1鱴w8\c�����	�s}�چ�S�)Z`��)MM�i�r����Ő�na{���F�OZ�C����$g�kk���:�f���aST�Uo�J�%��9z���PH��ΰ�t�c� ��1�,y�� ��;T�?����"�d�����{j��R����hN���)p1�P�фT�G�F�g��L�����q)Mo�-�H~PZ|�����%�BFA���.D�UF�{DH���B�\
��|Ko� DK�`~Y�\9�R!�(������L���dd(!����n�#N~�$>����W����e�C��6�n��
$VA~�U1�����
�KX�ʲ��se ���`t�/@�A7��05u.}��j���MV=8T�>Ddz��bW7�9�q��(��q=���^��^{f�ѵ?� &g��ٿ�����AԨw./�e>D��-�_�84��h���/�/&Fk��F
dYCx>�Z�$C������UZ�1�47�!L�m�t��������n�mC0T��O��_���v�w���֨��e"�0��23!^� �,Rى�7�;�ʏ7U�l�*�ٟ�x����q���0�=� k�6lj-n���ʚӢy��@���=c�Ƹ�����Wc2=�M�ٻ�����>vJS����2�gH����뀫!��s�Ɩ��� �)�E�S���+~�eku�
� �^�� |:[?:'��ü�уJ=�#���賶��������Mvr����{%H*3EK�@��{?�[��$�)>7�����a�=���g�*��	�e��"KƘ}^3��ʌ"���Q-��t�c�:�跶������O����Ci����WA�;[���W��٣�o�D��lֺ���i�ʟg��r�<�g��GM\�
\���ނ���r�g�A8Y'�������B���O�҂��WYȴx1���imRj|������g���э	��.������>>a-����
��Z nx�wac���p��y������l=mF�Qi�ų������ϳ=6SE�F���Hણ��z/
M;|��R�s`D