��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��%��-��p�g/�3��mC�C�;[ah��g�pk�˂��l~�<���]��DC�t�M�E��5p�� ��ֲ(ʧk&��q?�������N_�;��J,�fN*Q��I����*����W��}�($��V�����N���5ݕ����I�YZ
���y�ފ D�$�ih�$޾� ��kh�)��t�	��gMaG�~�_v�(w�vk���h�Kɚ���`F�����:Ϯ`<�~Z�f��"{&8��{G��͒�t��r�U�yS,�� ��?�������N��ػ�v�*z�����r�|(�+H]��ve�-7i��`�A�Ei�|T��'��N�'�7z�>��K8�ұeU�3�6���͢Uk[��($�6w�5`'L8�=YQ�y�����j�GaQODT��A�]��Q~�5��v�}=�C�Ӯ�b*�Z�z���+~d�"UC�Z�G�u�D�g��(�$���>�D���!m&3��G���:�����wzl�ZL������W�� ���;�޵��9��Tgt�h��&���������͆j�+V�f���J���fȊ��(��h�,9�����R���f�z���@�5��s��A�����@:W��!���L��Dn2g��d�!`ia�����"�\P�]���c�j?.��i�قJ!4�.0h}�����[X~3#�T"���K��崑NKZn���K�`�OID�>@���UuL��z�C�p���llμ�ďH����ͳ��	g�����	�X�{!�Y�x7Ԯ	��,�a�(��B���aUɰe�̕������D�A�Gr}=+�" C�JNUtfTdb�&�׿n�gx��(oR{4\2�����6��_@���#�1�4��vAy-�/�T�׸`�ɳ̉n�0����g�6�M?�j�tX���oM���~c�2I+N���i����R%&������J�Gð�)4�p$�(�Fjz:蜷�1j����[2^�q�t��5�<�5U�v���5-w">3#�mp޶�l*��"�+��� �=�i�Z�'BZ?;�������������m�N���%���t��q��b�˂h^V�ۡ=�z�9M��(@2�0:��i��T���3i����r\:��v��?�u�q�R�$3jhq���(V��[/�f�q�;�Ǳ;2!+$�PMj��LH\E��$��
�<�zxl-�'���bG�m5�e[�QAHw���q���
�ޗUE��q{%>�`v�߰�l/�B51&|+@�E]Re�����q|")�rB��:��fY�t�d 2�qh�T�CsnI=ߣTK�O`Ɲ�s]�}����[�if�HC�K�Y?����hzD��4���ݾ)��N�>^}��}�n�f����+���Dh]��qmd㽟w�>�Rg��rGCA�lʚ�{c$@�br8�G�@��/��.&�1ҳ<:�u��>��r����/���S�C���V0ǯ^�D!���e�C�daM���,�9���qT�V��$S�V4xb�&v!�-\�^d�<��Qʝ��OY�����Dz輻�f�fO��@����k� 5���S�NMM"!L��^I��l���m�v�(4�%� /㺆�g8'��x�k:��q��+E����^�1�N>/��ǭ̚��ɇ.q5���)�GF��Vid$�Ո��ZT1�I��j���Vdo�7r׵C00�3�u�q�F�3�9�5�̍�Y�Z7���꼜��?�Ձ�7�vAb���v㾏RA��zYZ�O���Q� ��F����@�x�c���)=��9�,���=BfX��(bqa���U�<gD�ܦ7j7�jt(�/�$XpOkQ�：4WC��8n9�i��2Z�tn���OB�U{ ���ؿ��P�/��ijG��:t|xuA����e��
~�!��l
���< \�f�44+���R���{���u��^\�����Я�rG�+�/蹋��V�"��45`}R��%��p���+��ΰ�_[��{C��iz���{� g���߿8�*+U2)��ˆ id�̑-G�v�w&,Kҧ��&�y����Ȕw3��EW��[u�&,(�t���	�:��C���Z�7� ��5M�q�ŘJ��G?��)).K��a�� [�w�̝l\����0L���l��h�,�$c��ë�9\�ޭ8����G<M��IR�YLKA�3��d"-���,&X�[�p���ò��,����Ӂ�Ӛ�5(�'O�X��C�zLWTFչg=|Gt�n9�֠���E]#��z�>�W�޾���A����oL!]eo*�ϗ�L�5<o��X�g��u�c������ܙ���l]�
��`U`�1�j�g���;�&V�I���A^F�6CM]8�YxUηp-�
H
q�Zo�� ų�uQ���er^g���kI�bbR�s?ov�Q�#V�z�/-�����J�$F@&}e�KN)�c�?|�����Z	6?�����f6/��B�/�02�V	߲���i�{U��%qʁ���:����7k��m<Hԏ��o�K����&�n��/Jp���<p������#��h�j�������7>Hdv�UX�g��c�>�#"x��x����1��B����]�D��ᛲ׹���uwdguLd7�$����c�Ƙ��BF���6<bcFd�P���nrDl��o�ڗ�.�c�.��.p&��!����7]C�� N=A_��~�$s�ӮR�F�z�+��,˪K����-^+�c^�H2� �b�0��%7<}���T�L�����U@۳Jû�Yp=mAfH]��(l���Q5���n�s�#g���A#��X.�5R�jFb��$�+�l0��_��z��-�6�5�Pw���uP�8�RMt"�����^�J�N��S�/�U~��?�&���9]��M����0C����WҠ�\�`�5�<��K�8�d#��`����)B�͵x��o4��qĿZ8������d��O (n]�b�+;9j�_��I!X!��X(<�O5�q=���c
+:�@T^���84��"���B�	�+\e����~��o6�6c�5�㚥��Ȟ�1�����q�(Í���#�(ѣ���5ݡ��})�ЙZ�B����PDf0�d_3�}����ԮGF�_��F4�U�g�
�1�*״F�z�����G_^���R^t���+�';S,}�I�qZ��������J���C�@&< ���A�!��w�l|h��f6oɰ���z�?w�d�m2ѡ@�J��H�~�.|���!�P$$����h���rs� r���s:����7:j�L|Gk��ݓ_�M6��5pHZ�C�u���pMי
��+x|i�oPl��5P�pg�lu`�m�̒�PƎ�0ũs�AZ�+��FV�0�Z�����I\z��V��o�E3�O�7(�
ڽ#b������ֹN$CEN��k��ȉ�&�c`\�Rѭ���U�
MI3�O0���S�$�Z\�Ne���U��{�Ŀ�@��-�>�,t~���X*G�k�jsz���E�܎*�$���Cvh��ڛ]H�-iKP�/���p1E�
~�+^�b�3����Չ��`#�t"K(L��%�
�y��3N�י�ӳ�Х��'�2�%�1�H��k67(�<���������xA�~g�+�t�\[sp	ԩ���q���ԥ-qy���d�v��@Q�~�"f�+y�qY�'���y?�[AJ#<�;�� K�dnNݜ9:9��,��HGyx�q9�CtXƣW�?v:9��o����'��<����	|y���4d~����]�X����z���Em�H>l�؞��[�����$�ӽN-��rU'��ݴ݆�POb�7~f5������2���D��L�Oѯ����1��U�s�X���#�f��o"�ϭ�����d۲����g����~ۺ���6�} [m>�nպoј�TT�k�îe�Mث