��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P���<߸�A��4��qkl����q.�7o�X��ږP�6�B�w���tT� �m�T'�b�n� ¶p4LB�$~^�c�۫#f��!�H��9#�u((�	���'��Rsী�Bg����ω�a&e1*���a����m�T��!@?�iwS*�����a4�l��8�Z�0gB������9tK6��Oj�$*^�bqe�yM�k `���_�N�X,�u��_l���i��EƵ���W�⒌W:LU0�:��ɔ|��EX��贱��hvW�}*8�� <X0FH�S�G�7u ݔ;�V��;��*� Nbq*;X��צE6,��+�o�J�� ��Et5uJ%2�5�UL�&4�T'@.*�z>;�_+����*�ن���.�L7��\�xQ�R����1��_g�o�A��N<5�c��8�k������c�T*�L�t�g��6�̼<�<�'D60��Z�{~/q�=� �Q�h����(�hr�<����+ad����� �w~PS�Z{<I<���C�֢ͅTl9w�M3@;�� ��=]�D�n��BI\:qM�uя|�`��K�����`������z����"�|j�OW�1������[�+�t!��OtV�3��|�9�v!�y�P;3d�,�_�gg)���x�7�.����Ҝ{��c�0̴8�f�/>Gy�
�"���6�K��βX��L:���`Ȗ�y ~���Ht��e�N"I�#�E������q���2ʌ��$.^��V��Mu�S& 3<�9T�Z�I�)2�@��5�`�'��ͽ�~�� ��d�Nˇn��
�>e�R4�u4�$_���a��Y�p�0���ۑT�TKW0Ĳ4�Q�S �����h��g�#�NF�sT�kyIX�胘U��W�1��#DMz�*s�1�gat�7_���{Q>�ݚ�d
n�]�\Ǖ���Uo��������B9�D`5=Nm7�z����_�hEOV{&����o[��n��&hg̪'�f������~��y����U�t=��Jܻ
:��8�q�t�l��M��$��j��j�i����x��BÝ��|�����$�ߔ�%cAx���8��ώ.~y:�����THPm����bc�-�%�{�KB[���������A׊į�riGQ���9�B�e&�Ϻ'����@�T�ݭ���]�����8�S�b�[쯻-�(�rT�A���B����G�گf����"�j���@zl��$e� b�T��=���ׂr���P�g/*x/ظ�a�q���Pz��-@W<�Иb
`*P'S
$�|L�)�1z�S�wG�~R��R�"7��}�nb�|]�c�C{��H���
Z��a)�y�v�PҲ���<��>���N h�KWp�!�s���^�U��ܨv`�|�\A�������Xw���4T����S`���whJ�l��~���ye3b��,�T������`�^��&�ɞώ�ѭWO=������;EQ:��8��a��[8�+�]��<�l��x+́��rH��i�g� 4ܦ�jm�&V�'~��ZoS��u�>'����f":-��-�5�Z��[˳ET�(�	�Y��e�a�q�>����p?��L�J�*�ؓy��B���=�Fym����#[u�|_�R�F�ߣ<��������Ҹ���)���?�%cMo�7�4�qB�v��#Џ6��ysu��R�폵s�F�(�ֆ���y���榑@�{`Q|�����D�s%��H������3�z-�yq�z�Z����5x�ʹ猺�QwBY�u��e4֜ړn�v�.��wZ,�c��f�OiL����}�^���r<��X��qա�?����ˤ��}��H�c�����l�97�y	�Y��p��/նQ��C��
�)z3=�����QR�/��!"ݲ��rWJD��]��ǽFlw7���_�Nqr	����q?��φ��v q���J�Sf�����5�ʑ��z=�jз�N��ľ����4Z��%�xf5�����k��9:d���p��[$�-���߂�Ï�L%��9���S�\.�+����p*{���I���s���ޤ1��V=m2W"3��U������;�Br�`Q��/���G���6�C��҈FV��>��W���^t�K"��5B��$��Q�tU����i����+	�KE;�C�>��Y�E���в�2/>�9�K�mz�c��y�D"[; �˼y�$s��MΗ�ׂ�%
oI�w���~����JO?1�T�m���Y9�rt�'�e�ԇ�f ��܎zkȪ�0�]ܹ��&Rص���E��/���IOj��5S���I+r�h<����g��$!A�,�L���jUd�w����pk� Q��I�Ȟ�4 e�Y����(��W�42Pw�.!��ҙc���g�r ������cR���X�|��-L�h�8
Z�4J�hK%�߅�,d8Ydrhޱ{�/��O�}�SP3z[2�Y��=�7^1SA����2�Mml0�n�u;�V�H[hy���ô|)jG���5�.� M����-c4�_{�D�Bp��ͯ��4��߶:��Y[˄����d�Sx�I��By������z�{#���{Ȱ�s�6�׳fG�J��%�J�'�8ĉ�]UzcK��+9�3��e|����Dbt)0��  ��F�����iL�Y�e���V&�ㄶ�km} �u�fn{����\Cj�!�X!yqN\�G���sD�]�������1���Ӌ�p�������!�2{���#��~2���3��6���P�y��=!R�[`�%9�@�vr�ŉx?�*ڔ�m4y*�l�I��q>�$��x�&�(k�}D`)������r���L����RO줥�j%�ʐbi?i̢���:{}�\*s�碏q�\��3���wp�N8��(�r��ʛ��8����:ʶK ע�)��+	�/���

���Ke�����^��SnC��G������*�3ĩ���>${�C��qV�S�Y�u��K���#@�t+Tg?��رy�le��}�u��n��&��앯|
#\�UҁR�tӵfa?��bn��y�y�I��c���U��x~�ט~����a%�h^K��	�4��#���2[ +��I��R�3B�h� �k�x������:�tE>��2�6�A��uG�M��OF�&�3���1憓����<h�>�sǽYR��t��v���J �����L@�*��V�k{9)ǐ�0+J	I�XT����FMa��a��3E�ś)/EϤ���������|=!����`Ս�C_�=;�Q����[��_<�z=�C��6
~yo������4ȪcE��� 
	MF��3��d�X�:mv'B�Dz\5l8qAa�����>t�	c�Q�D�P�+f��K@p*O*����(�m�qQ�,*��\J��i(x���u&i�|�c�yL��j�Xr�$9����D�Q���l�9ݷ:��YMJTZ�-�%�F]������̋�}ß���N��5�H��s�&_¬	��`xnm�)���S�f�C�lY��f�c���|h��'J��=/dB�[:}e�$�@<��07�q!>nP�O��'��c_/���R:��U����W0���������+�2��z����	�{E����D\�����ڶ@��ÏoL�-��O��QA-�3X=�'��9���M��e}ށ��c�3� ��\˹�SS6��e���̱[>���b�3w����b2�ιއe�y�~$��j�<�$�x�`D���B�J�}�Q��K���W�JJ����s�kK�����񀢮Bfn��rnme�[�[�K��bc���*�#�/�z���p���MzcN/ ]�9�{��M�s/ʘڠ��+��Z�yM-0%�ts>����1��,G3S<=	*���Yh�N�Y�UP;p��R%޲�_K��ok��f�|-��u]^�!�)'�L��m���>�~�K*1���7�(�����ڼ]�v�*��q	{3�U��>�62� FD����^��юiI�y��,��v��Q�(Qx$�i�-k5����`���9 @����&��*����CƬ�:���c��!�I21[X�	Z�c�4@$��bG_,�]�����\Y,���>�k�������ܾ���=܇�֍lp3-Bw�hP|��=��>A!�g��h�Sm~V������TЙ�{����7��f�­:9��3\h'@$,a��9��g��|�T�I+p"��K<9�����[���vQ�Ÿ4.>��uP��[�๧{;�w��JY
֑��bz���mI�;KjZ+il.�V]Z&�g�;�Y![��t�w�vev�~U�K���LD��Ȳ
9���d����*�XW(��A[s�����A{Ȩ缠�-����j��\,w�:��i��B�?��,&��J�@�Cu̧�kvӪ��\�a��Q�2�k�Y�F�Gi��4�'k���-�D�	��q�1�h@��0��� )`S�$���&i^�/��M���l����>,E�| �L�4�I�_��hf��j3�;�e�%T4V��%� �5��'��+��&�\�⎸J�-���b�z��m��R��]��W��!.�V��w+:��I:��rHS���t17�d�gbD������(lLd4._*�ƒ�hv��z�l�T�����B��ɍ�T��R��8vY^jsi�?�;L�w3T���B(���*���{:�(P!��ܹ��QAF�ʖU�;�q��f檀��0�A�l*w_���k�gi�n�r�G�~�|����}
S?d� i��t�<i>�M��X�U�Ipzկ�I���V�:O�QU��k5��iVuڲ7��kgk_�g�Vi��ٍ��`8�f�M�5�G��Z���q\��].W~�P�Q'��rZy<B�P��A������ņ����UO��[B�{m�[��h�|,1�y�b]Ls�Q|/��EY�M�r�f?st�G�)�&0iG�v��;���&S��rj�:�o/�5��rp�����DP��{z�"�M���dķ9�]·�
|@�< ����fP����`�_��S�]3�L}��d�-O�a�������C��j|Us�h�k&��(�)�Yd�nᝎ�B������K��#?�+�b� ՞vh�"�v�q�M���<M���Ȍj� շ�]Рq�%�Ţ��i�����W�pd.��5z�%�Z�L�4ܳ'�u.^N�D����=u�ͼ�8;��,��K|0�+��1��
f���P��-Td�U )�t��_���& ��VZ��w��*,N����%1e�Mm�
n�@�  ���Q�z�N��uRc{��a� "ﺎ�x�`����a?BY�fP�ļ`��<'C���V���H�Q���B=/� ��=n� ��m�����L%�Vջ3�.AGS�&�&3J�W'-�f��H�b�_Z5��}����KSϳ�$�0J: �pL��^|>�EC�yả	�A�&�D[E�D��JG*A��@5�j6w��}���������nD�%X@
剭�%�w������+�V��<r� z7h����&�Sa9{�!I(Of�L�ڹ��AE筦�Ƿ~�+�FNt�ۯ�F�
\i��k�~�� ��L�q��N���vs�	MIpP� 6��Q!CE�Dm (W2,�	�e|�����K�Y��R���֘�|?��{�x� ���ܬ���=S�gq?֡�3r��M �2<Y�#$O��[w�O.�8B!K�g؆<�=)���S����7"��"���[Uy8Y44���qj��<=pjF������V�G�ӌ�|��:����1ң���-�ݟ�i��R�-W�L�>��ċ�F�҃�K�(�*�c�bߘN���U����]-�v$����7�
%�%o��F�T�A��W�`Jh+�~��֯�� kN�k
^ AB�j7�ʖ���B����4�[bwߓ�غ�o�R>�?���>��hOi_�a�4��c�@H���N
;
�ތW������i�4N9���6qndc���G�4h�6[֎+�b&�4`��۶� {	���JAnj�K��'���C�!o���0B��'��4k߅�`
w�a�'���c6]!�C���7�R�̀�>h=օ��U���q����E�yB�;*��wu+wKzl|R�H(Q2�5��r�Ү���1��׳��K�Mm^I���B�9��s�4�r����Ϣ��H�B=�"O�=Y�'g�k���Uǜع�K�SE��Ζ<����M��<
	2�߱ϻ���w*���̷���<S����v�<�3�n��������巜���