��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>�����{I��v:?�BÅxJ�B����f�d���n�,o4ʣ�Rd2V��&����q�B��$I툒GM@�m��O�+N���K=��~���y7���{<�����(�Q�4�.�����BbLS�K�,�ݡ�&-��-��L.}��7I��L�p����U����eT�O`(+0�d����GK �<V"=����)��*������/����PY[I����n��l�è3��ML����59�ā�#k[y����%/�7��� �>��{��*�hv�&9n�G�OO���{�9Oo'1#gP:�S�0�z����?�w�'y����_N�:f��0!\���١�rJ��nJ��~
8� S-����L1<�Cj�,~OB	^&��Mt�t ":]Ej��$������T�z����Q�(M��<qv�:����E�uje|��lg���p�6�bb��Y/m�?�de�Q�'�ȅ��-�J�)\�Y�jR*G�P��	GЫ�f/����rW8�����I_�Tt�p&?ۙpo�3�O44d���@�qu �;̥Ȁ�.K�v�Q�FZ���BtL\w�% F��p��P#:}Ȏ4i�3L镦��Ѿ˲op5CF�n���S̞B`����V�n$�@w�W�aΡ}�$��J���.}��[����j�h�\���7����/"R/[֠�B:��P ^N!S9�:���S�����w����>�7{� }��Gf�+3��~�8��]G�i�j!�*y�O����K��� �$�u��V
J92(����4,r�(��"F�ԡ��U&e�E �`��F����:��"h��<!n�&����n���{7�����l������g��?)rz�f �Ǌ�Ğ@<lJ��#�c
��d�	�ЌFE���]R���&#�	5jw�Q���Hk�u6N$Y����ˏ�^�̙�5��5� �Z���s�/�7��yw����l�Q�T���?�g9:n��b�
�`�T�څy���.ʊ� ���j({��&�aS��}*M�p$�{z������}|t㕊!���)���*hT���?�~7��PWi+D٫�J��)����FZ1EYg�;,�����>/�&B���|?��ŗa�F־�f�aA&
���<�P��y�:X���P�I3��:��LR��}Sp}ҙ�����BޑR�V���,b�#ٞ��Y� ��=�CK��05�45K'�-2`3n?Y`$�7>����U�K>@c�0�\1f��/���)wwЮ�F��4�-��"�B����e��\���1|�T�U���"�=�K�4��ӷ�A!��?�娜<�ى�E}l�4��P^H��Ty��|ְ�֘��J����SL܌T��9���yJ4�M�pȿ��50�{�=�3q����۳I!_	���e)B��$���\���QP�%�J���w��=ڧf�k��{����/�Zi�V���t�G,*n�{�����?9K��ZW�Y)ath�Ɵݚ�F��'l����/��V|<Qh����&g�[Mb������aq��Ãum�7�Lj�g仴-���G� �Z\k���ȟ�Rm�am��ݩYY@���9HϬh6NR���m&Z��@`^fç�z���C��$y� �qZi��Ȟ��K��	�p|��U���.P1C��n�����|W�;.�૿�5�'�j���8��WӔ��wjg�(���֖9�^(�R�m 1�1�X��c�h�Hᾥ
�s�:.����<�{��lL"E��eF����O?���\4�:��M1��+�����A��%�P���H'kE*Ld�.ֲg�w'@3�g�7���p�$�[3
 γ�F��]��V�(��T���ưp���6�{T�b�#O0�#��4�$m�d��MgM�m���K��l�	L�8B C�='��˟�fipej�)Ή�~�������~�!]��p ^�.��d�]�%=�!R�L	d\ˤF�p'����p�9��&�=M©���Q[�A�����2r�"ф(ߠS��	\Xџ�f�7i�"� }��7ו|&�� ��Hiu�۾�[u`�*j��tM�R���Jsf�͏2V�������
t�j�P�H��8XҎ��S�R��GR���tf�f������ibA���p>����YA��q�b��3p�S�@�}J����T̛�ˍ$���
!ū�E�$��!��l�,I�e�8	��)�����A�^�o��@2���s�;����E6�q�e�(a���o�\+!L�����}�	�<]J1�c�'
:�)(�3?[ΧgGv�\�@7�٩/��ӱ\=���ړ%���]k���A���#��(=�
�a@���l-�tE�j��w���E6a[I5 F<��G���l�X��%*��7�$����[2��A������J�ʘ�h�a���K�u_K�⭭B?�	���%�Wt:�Ls��rΖ�掏v��0%�>"J7���Y �Е�u��+	gA K�M祔����Ǐ�{Sꐻn���]>̾�12���'�ߠ�|M]`�_����y&7&��P,KYG�#�������Ԫ��؀�e�F�Jl��8OI-�}�0EzЦ��P�wf�q��覷����K�oP7�ޤ[�`�1L��r�M�"�V����
e��ib�7$��qt$~t��r��,�f���$�!C�����fvf$�����pq�r*�mT�
@���}��*#� �s����w���kZ;�m8a�\���R�G#����c-�X�Yݐ]�z�LH=I��c!�;�CQ��%y�.7���"�w/���[�)��ml��i�Gh˕��wǶ���=1���{����J��X�&��9�V�r���
����1�V�W1�ϳ����Ů�P�Ԏ���$7-�Ȉ2�{ٶ�\z�y��{s9N-��	�������w(n�Tx���!��k�~U��wb�����T��x�>c`}4�g�������0 BlϨQ��N�Rq��l#a��λx�����;�_��Y�TC�S�F��Τ^�~#�'v�t��A�
QrD��̖��*w7Fs� ����������V�������0f$�5�e���F1�7��t�ܖt�h��|ziZ��:K`l���Cṋ+�#Eo�>`L�� 6�P�(2?L~����\W>#�x�ª��G���ʀFA�Ф'YWՏ��7g9�~S���)�]i���$��O�����uJ\�G�1 �F� �������d%�3�(�2K�SyQ�I&$��!ә)��J���[E�|�r�?l(:��8�-E4��w��8��������]N�$�g�!lW�k���8��@@^_����L�DQ}�_�Q������[��ǣ�y��`��A�������es��/P9��\�ɩ8�k�]m�v�gXf���{0�`���r?Www�r]#�i�skv�yu�Z�ӄ-ʽ�v�~����4)��A=��v2�lr���c�ߙ��,�fR���,vyj�MPhY��������ŎiL���D�L�X�;�ͷ�?�a�|��g���K�ї�s�<z���^����Ņ���m�����o~��R�>��U�3X�ҩ���Q�2�Gf	�d����i�zƈB_F�"�������Vځ)Ar9$X�f�c�u�~!Ԅ�?\6��3k���Q�	w��mA���GX,�g#�ٞJ�
]�i(�v{i���TZ~e7�l�l�f�7�k��k�*�y�V��\*C�)"j��7�*��V�e2���!��,s8��Q55�%K^�,c�=���TשX
�ݛzw��
��@�A|T�6>s
����������p���xT�K�U�r!��� �s�d��s��^C�0?�2�51�Jq�Nf��N�4�R�%�'^?�.J�[��Q5��[�v��/|�-�WDF�y1���h �\`���2�n�^k��f��߲Д΀X��XM�y�<b=�-l�/z��Z�߶�� ��L��6-1���J]���^����k�Uj=�����Ŋw�>��y�Qח���>M��6��-&`L�y�)�wBf��?_&�qBU�k�{f���I���1۞c�5Tǎ٦4x��`�C��?q�rL�4^ݗεeڐ��2D��P�U�k��7��ۜڠ����������>���#�u����3��(�ɻuk�.�j�^���Qqf<��	}��n{��&�yPצ@��@��1���ۇ �ɾH���d9�l��ҙ:��c�K*<k���a�+�歪�(��N��d1e�=Y2���Ӱ�c
�*R$а�yy~�𨼢�!/a$������*j�8��m�����G�w���B@��kX�F=��!,��P����(�c�Sֆ��j/��ԍ� �v���3&+]S���5��	��%�N ;�f����O<�?��5aJs�������*�$
��^�m[���\�3���5����TS���)����F�"������wX��s��`M��Dչ��>�}G	,0�9�cRS ���5�x�_,E��o.Z��x�w%ns �Ŏ���ٓ# �og8j"�,�!�Э;|Z�5S�����*�m�HW#�� rw��Z��������tq�|S�YȔZ�Z�i�/�9I*G+<u>eO2�NIBFxgk�[�g%��zY����R�_�����܄*�ѳ`>$�{���Ro�J"�1F�G};!��\x��b�̕C�
���c�_*�����~��<�Ӏoώ�`���ч�E�@9�pZ8�~�������Iyzϴ�1-��
f�Z�T�+9�2��;W�k��u�#�|��>
����Iۦ�D�
:��ZQ�J oD@���Y�<��33��-+X��x�cu�;$���am���.��!uX(�����{�fS�z1ep�eu���q��P6���a[���΀�0�����ک\�j�}r�N��.ӷ`�RԳJPw��[k��X>3�y�I�4\��{N��L�=X�Mbr�G�K/��ѐ�S����.D"�I�#��'c��Rw;S�bN�N�uwz��u�4�U$�s,3�j0`�[Ҵ�bz_Ǹ�Ҟ�3^˹q��AR�I�?�_,�@����v����E30��13pAw�1O�ݎk>�����t��n����~�KԳI�Y�s	?�-ae�o����������;ˇU�IY/��w�W-8/?���T�Yy0�ࠤ�`���<+(�f��`�(�R�:�֙��2<J[.+cimb�Ͽ�������>��+$�l"���΂��`���3���FX
>Z^գ�)(�dʣŠ���+ո�`.�O�r�p�7n��.��؍b���dU\df�X��|�R��)�_��}N�h�E���(�e�ɤ0�1k���=p�ݩ�JP��%�WzZp���&��ܥ�����L��m���N��(U��J-G�C����J�N��rο���OY�����䜋��a���[��/l	>ni�Y�lf�s�����6�vPjA���D}̔#�/J'���B� ��iK[�_�k;�Pױ'����\��r��Q}�=�a�k�<(t+�:	J�Y�M:�A�ǳ/�r��)��R�$�#�z� Y���:��?,ua�>�u3E�@���v����W���^V���bdr��,K� �Q��*'�_�qк�ذS���R8�آ�s���	`�'�'>�Y	����Fqlr�.(��~.c���kL=T����!H�kg�`z�
{��u��q�ExQ��j G<��		M�?Y��+_X{�%��hM�+,��|��-�;&P��U�չ����E6��~,#ћ�,�Y
�b�"eł�' ��knj4����w�����ˇ�]��[��cR]�i�R����ǣ�^!n��Nd�֛�7��l�(IJ9nS����Db	��0i�D��8��M"K;1Ɠ���͎��Y|\U5/t��ո�_O-z� Cj��?��ڳ ��׵%E��2�7���(Y�t��9�6܎H=c(�u�Ac�*�0|úA�5���a�d3�kK+Cf���Jidx�C�*2��w젾Y.��2끞H�0��Z,�\�T)6�QF���:�uH���la��!�����m�������z�}�>W�S��)����b�F"Θ�6�\���y�%5Nш��<v� �	�1��a)��(�����GY����[r;���~Q���
݊	�>�/�f�$O���V�Ʒ�K������oz}�C��a2z����M�2M��|E��ˤ���?��@�n��f�A5B�#UG
tͫXvn�Xޅ|J��P
��|
{>�f�������%�i��)6����ԜM�BK��	�t(I��干��-��M(ݲ�\�N3�~��ZAL]6����1��`�$.�GE�x����xՌ}�׏/�T�.Wp6S�A�����ΐB�H�%_S_�r�Eǚ����3��a�T�[�y��0'XC���/�S � s?<�'F���9�ʫ"��SgW�o5�R�NF���y��긓oG�шm�D�o�쌃����U����ё���r����?b�Km(�:��]�B�Gϒݶ# �X�$?�R�!Ȕ��Y��V4��%N�?�I�_�3|�6Ns�bJ�џk�o�R����Z�]w��d����E�$���eӺ���H �ɏ룆X�-ٗ�+��:���h�m������v��<@��xʽ�39w���d����B���r�BR=X(2��F�#�t�ߡwU�w݇T1����J���,f@�.&��o��J�wI��̸T.Ug�ɳƏ �X yJ�X���#���4�Ӟ���&�39u�J�K��}�����8
�4ەĶ�眺�!��d������ެ�`�O;��y������2�:OO�`��!4������Tw1�OCHJ�� �K�)�v���/���ê�?�a���L@�2�a6�S��(nOp�rT��a�\1䎑U���{�{1���պBJ��y�^9��Fx0���J+o��	GvD��κ{��ʜ\��� B���*��ǵ8��G��w �tq5�������?IG���6�u�g6L�Q�E�oo�O�\��� �ظ�0J<<l����t���4�7E��3���l߯L�v
�QuH�,��R?�k����k�-����x�|��m�諽R�����4��e|�j�k��NyPCZO��#�*E����/���/��Q��̽�;���Bo�ً<��5@T۟�/B��m�����,~����5�=���Ը�{Ը���`���}��� �eA�Fj�ڟ�[�]ND�>zؖc��t2պ�L�ă��<�R$~�xe�a�����;i �]��]��<�:0%�!��R�d��B�{��ͱq({��%�d��.��?��i�ؔ�@)���LMM���gG�=�n0,@w�~�a�����]jp����;���s�� 3���(��u�k�����K(�eRw��%(gE�����g�]��ݗ]h��n�E��o�C�&�ߜ�`�~���f|Uef
F�V�'P\����+[�	������d�=_�)F�Zx���l���?!�)�����ޔ_�3j�?߽09}f�c�	���Ag5ap�Ѝ�9��D��؊���ڢD�v�] =)��&��d❮q��d <U�h�hx� E��Yo�}���,���
�8�-��ܝ� A�=7�+���XX\�B��xl��FHsA\���+{!7�1���6Xcb��7�����q3o�ҷ�qB��"�î��8��@�[K�<\b1�s)���++C���|����kR'�ȼ�o����M�jpn(8��&Rߤ�p-���28v�%��$Rq!�:����� ���*�>L�۫�f�xٹ~�a	�Ȯe�t�y��7Ѩ~w����>g]3a�ތ� �sr���+=�<:"˅��!��e�W��|����Ћ�u��``���J��v��hY�����L"$�I�� ���� ]f��j��D#r��0�
C�n�;���;N��-�K8�0mkm����~��Y��HA�E�N Ѡ8gB����V�i�؞Z �G
u@��H �`��?u��c��zU-�w�fJT��G��!@I�J�]z���"��lʥ��Iw�_ӆ+��t"�p(~j�$T�.%5�S��A�H�tޑP����1ش�@@����a�����Dڠ|�����0o�x�2,�ŵ-"�ٺ�� �D�����+�'��i��<I2�믨<��@���C��D2��83�H��'bl�d?Tr�6<���j0�%)�����yqݮ-��]��~�ʘ��as2��T(�o#�/%h��E9����� ^����PW$\�*�)-;����7 ��;�܉�?(VS�wܝS�
io��E�<@��|Pߖ�eL�0��n�����Y:&���6�U��G�w-^�T�v�w�8�nJ�' �obhG�)!�I�#\��X�3�$RU�-h7�`�;+��i,�c���W(��#]�zgo\²V��H*�T�|R�&��`74��>G�A����Hy�-qm�;d��	�rEK
j���QD�,�$q��R�	���))
�m��4�<��eN�хMwv�����kg0sfJ`��U�KR"FĪ�Ŵ+ ��#��[zk�Zx?�՜��1����rK^#�sK� �b&2r���5�����]/o��m�d9���MG�t �(ES��z��;D�q{&]B�t�&S�-�����B�/|�}�3��5r�L=DD���\���s{zo�8 lE�:5]�C+���7�F�7�,�rg��oӥE)�rGu�f�f�]ks��~&�+?w`�� �v���u(ⓩ-),�F9�7�4y�\^����*���� :��a������;`U��J�c��W�s�њ?�/tY�LG�nfݒÚ�S�gV7�b+W�&8;%$�6�a���:^^.��V�L����0N-6t�=�YF���W�Xl�a]�1�����������]�(Î�@�V��*�lHV�]�{�r������16��
U����Y\m�#�d���h�e�Ο>���^ܩݸ�0ۋ���C�)����/Y`qa�>�j���q|�<q����q�;s�4��rę��Ώ��/E�?�����w��a�Pg]��Qz �`���wՍO#Qץg�D�����Kos��:XϜ�ͅm̊�� ϥ�ۦ=���γ�c����~7�ާ�u|_�`Vk�!��kH��1�W��JE-��P&^��=�5���26�m
*Ҟ����C�����O��M�ݓ��f����Ѝ�7���2��H�|v�sɛ�m��_e=�;�Ｑ�6�NP����i�O���nb"Ӛ�AR3GXP�ׄ�+IRmu�^KlE���˚t� �_(�>~����#��9a%]�r��3?�k1r��	� 2�Σ�$ۭ�nm!8�pHù��������_q�3�H�ä��{OsFW:ԝ�Y4���mR&�w)D�@W�� a ��w��&@�������E
adL������N���0�����XC��7 �L���������O�Zt�!��W(�����Ă��,�0�􄅎	���o� m+�qJ�w�1L�5��IK7�NP܀D��q~���ܜ\�IE�����G3U�{uz��0$�(�m��84�$FY]U�!�EIC;�Tf}��O�9Zw3����f�`�\����o8pܺ:ܚ�A*Q��%}z����@1yi��=L	�_��L�ʃ��!��3lG���A�ɋ�p��J�c(cms�G���O�����E�lܿ���X�xID��{��q�1đ�xq���]@�N��6SZgN4��$7~N��I��`UhR�e�'&��S��C2Z��;X���f@���������Te/Ѓ*�``����J6\C?�i�̪�3�KE�_���� K�:�pO�޶�����N�!�����!v���=B��è�{���pz��-r��x�'�|m�H!�����z������>��FqE�fK3�ij3�?hVG����a��Q��,�J+*��n����e1��`w��G��AY���oK��i��՘N�]b$�v��;Y�|��]R6fY������A����q��R����s�����v�rIO���s�k��;�oаW�!���@+�閭��ޥG�\�6,���O"&�"`Q���DE��{#�HPo����_�p��TTke:��n۳ �Qe]��	����J�0��W}]�6��E����+U����	䐆�]7^[7_�۞�Ġ���0Rl�U�8��\�Fc�L����v��(*]���9Ǐ��3M��~zU ����!�t�B������5��I�Y���c�&�a���{� n�QrVC� ����`�8t�34;���d�eB:F���Ǹo�(�{[��(O���d��L���S���ۼ�F���_����h�,��s���jw��<�X���%���@HG��Z�}8�e�1$�8lhq
�3o�=��W䵩��t��bXd���t(�*���C�%G5��҇��ZAQ�Î�.pϳd$�.d��GF:�k	|?8�^i�kU� ���'� RO�b����_��2	�KE$2����%2��4n5����W�����k̟����Vantd�8����k��0k �W���2��ϵp	���e��|\�
h�zy��'i��&�Փ3s��W���2�N�BaBU�>��}�g��ln�މ��������N��`�B�*����:�ȷ� |��#aU��8~}���M��e6Cw�'m���޶�qo� T. y&���O�r���Q�f̰aPy
rP���W.�=�0�^�Y>�*J�?}�K�S�����ӷ�ߵZ����;&��xo�)�㲺�>�v��M��s\7�g�T�30s'9�o4�th�<�s��ܸ�����4�t#�R��( !8+�&m{��!�_�gK~f�.���$�����@=m�$�C�(���)\��i3��k��nC`T����>k�� z2��g����e�~�H�`�^tf9���S�7��;"9͘B�|�O�6�Y�cI��/i8ɩXx�y�����&�>��YL�×E�"o࿔�W����j%����/�`'n������ �p�|H+<v�,#�9"a�}p6Ͽ�f|��gY�i�UI�U'd8n�[*ҍ6���'�e�t��!D�B�� P�@����c�^�����~�"J�>?�&��'ӓ~u�(k�N�xY�Dv^���F�S�?���fwJ�9
6��ͦJ��iе��)\4�;�~;#\����Gڕ�i�>=߇%�m���B���4��L)�H�S�%On�+��y�(Qf��2�����#�:�c����/`��ȍ�C�`^�Z=_��/W����sjc{j��G2�(j�B+�2�J%�Ұ���J''���Y�u0v��o����fd:���>i�]�{�N+]ڢ5��؞��d��J8�_�����~����FN�� M��%m��FÆQ䵠���\;�IC����Z��a�[Kb�\y��a���ڭ3w���){��,V�WEb���`��RGw���������"���5iW:�Q�±d�P[����k��g*�Ɵ�D ��n>����F�XLr�h�Sfpe��#�?ۥ~z{թ4R�&2�ذҞ�mY*�2���.��_.qL�է�z瀌��6F֤�b�A���� �9���� �l���R�d�XgP���1���bF�\�R �;�}:%k�T�2ޙ1Y.WV��dȾؚܑ��y2q�z_XVf5�ܝ���_��JC ڀ.HtM��,��/'���FrU��c����Yu��L�(j߹Y����چ2��P)�d,L����p����9a�f��w7C��Q�\O���/�Qv�E
�)��C�-x�O��e04�M��d�:�����,)&A�@OG�l���-���j��Ҏ�^ۖ�6>�3PU	u���׵��9���K*���6db���4�<o)J&����@.��勐�� YG��	S�����|�bn�����������j�����H
N"0^�v{3�0�����f��9^K�������.�Ozɣ 0���2G����%�f�4pz�'��9G���f�_	�*�S��0���ޒ�pC�y��6JJ�FN����}��g�0B�����Z��(�9$�0#@�5y4�_[�9�n��0K��A�%:V�j%�~������M	���a���,q�
Յ���:+ĭ�"=R?�r��tq�-��&P�;tlI��O�_�%��Xx8����ͽ����!mW��6t�Ȋ҈w��*��4�C-���^����͉{ ��MeZ�-s�%���W���^Ri��?���WN�C5���;m֑�5{�{�Ϟ9h��:�E�N,�K�P�����-�B�����U>��i{S�@�%~hp,r��Z-�֍��� ���b�aˡbf�۟������hE�L-�H��5�q18�S���<�X�,m�����OW�(]Ń����m�c�dA���B�$Ͼ0� �8~�-��;<ֲ*g��B�U�4�8Mؑ1UϩC-=�E�L*�*$Oc]�je��'�"a���Gn�.��r����m�Mޘ1勬1H�'�8xI@&�9C���������y;�9�!�K�Z����'(U?��n���)�0UmwG���p��P�ڤ�н��Dƶ5�L
�b�z(��7Ze@�Ci��O(�U�}"0C}b��b��g"��?hS��=�l�������x��<>̯�W��D�|�1O.��:�&R/zn��?@�A�,�[\W�V1�ͪ\��'B������e[�����Cr#1�m�O8pȁ0���_�7}�#��ˤ)J���w@�/����b��b+ajN�+�S	�{�:p�C���pzۋ�՟{|ۣ�?�S+`����QGӪUM7D��Q=����b��D+�Kd�3sD�= �"K��x�+Ųc9+�>�˸�!PRs��B�ezd�$āfd�r��Oh�)	�3�����iK�Hn�GD��ԙ����1v���#�-�<�9z�Ie����S�&���O
�L�PN8���'�6�
A`+���]&C2�4�	��9�2Ê�����
}~��p��	���=9�was;���C��A#%��܋td=���F�_���H }���x��1�$i+}m��	��	� �ca��r���������I^�� ���i������-�����-q�9\l����0�:4���c�D�_ K�5]b4:��|xu���N �I��n  ٗ�Xuʵд7�k��8��"�X��-���W�#'�G/�u�� ����gY<|_�t6nD���Z��F[[pS� @ZD{�"� ����n���ױ�S�a$����������L�����ݕ1���Y�ɭ�J2��^�<�L������H%1�i�I����3g��	p�m�	�
/�m�-��q�I�b�'ڰQjo���HIޖh��l�ARJ���O�)Q�l�k>��CK��ȶp��J:�!(͢��{�_��� �]u�e��F�����g
�i��=*S�~�!\����� ��86����^�]�V5m���u�t)���ӈ��񈩙�̊F1P���`nD��%��A�soLPx���1q�Rh={盫D5y�5x�kf�ր�X�^ٲ�HΧ?���<�FR�?cN�J�xo{0��t 'd�n��W�,B�ַp	R6b�'����J,�d"⾅�PōO�:��tM�NV�u��*c2���J<���NHm��i��Ch����������.���msv���AjUR%�Oe �LC~_���EE��Q&)���Z�?��:�� #w����T�R�=�O��2`�B��>χM�?:�����d�~(�qn>\��]�O�N����%��L_�D~RǸש�HS)Q9�7��OZ�
:&T�YӋW�ilW��>��ES,P��R�C���S.F��/	W~\ث9�D	�@0��7���ܡ����7I��aIF� ΋�	��>���5��_|� ������F�O7��R3�{��>�U�2��(�b9�iSe��g� �ꯎ���A��~��ptʉD����������A���r���S�6w�dJ{�d��?J�W�~^C�i4��)��8�VNX�\�qx�nuݓ*sv� �d�c~@'�r�
m"WU%f�����S8����V�Y�H���?�"H}_K@Y�����J�|�PL�7w[�u?fo^�B��/�Ƴ�a�X�]���TǷ��$b"r��E��:�"x�8hn��]��*J/}Ϡj�H<u�.��^��M�x���;���@}F@���y��)�A�h[�����P��:#z�PE>"�
�(��������q8U�F�%>��>�֩"V�o�)�� xpG��2�Ǘz�ߋ��s�W0ZB$x}@��$TBQ�ߨ^�҆,�!�,jI�8��́B	�M_��k�8T܉�	����q
�J�]�m���҉`H1�]b|��6�D��v�L��
�`HU������>)h|9jZy�J.6��32-@�C�8U
�p�	X��C�a�ⴉw��R�]������(.��1�q�"͋p��?�B�K��^w�,����R�A�n¬��_�E��F8�y�J�k�V�u�Guyד�Q�������6�L��k���:�q�P*>��$ :�(S俅_/N�����<�M�d1X9��K��8c�Nx�cQB��#J/�s�!�����Sc�O�i�g��cm�'4��x�)�e�P�\5�-3���7�`�}2����m�#�R����^����]zm�� �ھ<��/W�WI�;㑮�����Q�����Fz�`1���%�w;�#��·�v�ϥ,��I�A>�7��v�D2���*�vE��S�X��p�F��j�">.�eY���l�3�.�$#��BH�ޠa��,ɰ�-����>@��m�����Q_��d1Tc�C�}��>�vJ5�R�I�e_z��;&<l�Y�sԝ���+�|Ά���h����=��֐4�Z�Y���et�53�1�}�Ա�g���p���v3�f��xl2�N�ᅉ4�N���]r�P���{�j:Ź�ei�	x��~�A�m��c�4?����	��f�e�s���{}��Ԓv�k�$`J�����ߜ'_���ϸ},AX��p+��?�ex_\-$d䗱n>�v&@	U9Zt�ҵ���4�R1�Ҏ�u�G]��b�&A���o�lIb&s�HW3?�DV_@��b����Y�U��������A�.���@j\O/�{�{&V���tATr�>
�w���~�|�.o���M�X��S�SP��L
~�<�T�vKk8���ۗ[C�1�<�e=A4�BW]F~��vߨ{�[�=i{ܛ#cZ�_���ӧB rƞ<\��	���k��g�Z�By�3��St�)����#��E"���_�2��}�Rk�"p�O�I�'2��'i�.��&Lp}�5;�f����k�?����t������{ҍ�Z�������m�.�f�	� �Grk�w���B�s���Y߁i���	��|5�j�]C0y�(�:g�N�Z�)]z~�?��i�9�L�,U�Q���ڲ ��j�o�V���$�8d-���	�fR9P�cT�JG�uWF���C�vԉ��=
DI���Ȝ��4���Zx��bf�>ɸ�5Z���V��Ɗ� r7����eE�|j��O�mS�@���(Ł��N|m/؝�CR�����eGLe��P��4��{]41���3��(-�>}�Z���|����M��?�E��"�&Dt\?�HF;�g~~(�Wb4���t����u���6X]cy��������y?tZ�U�B@���!a��qR{-%_6�J��������j�|6�Y���8ă�C5���8���y�k��d=���4����ǿ��5|n.k��h; �H�B�/�4���&����L�{,��e��v�A��wJ�*S"8����5��Q�)�B!�� ��[��j������H|��>f����C���	뼂�f����Jyä\!w�6��M	��j�$�'+f��*�/�}���K̀np���O����V����!�BF�i�������ĳ6���n���u�����\7�r�$�w��~���,��Pz�(��)�ϊ�f�bX7+oG��8��\||u���p���B��x���="f��1��V���g� �Ӿ���Ic�4�����&A*H���b���W��Y�^l�z�^ت!�ퟩ�<�Jm��2��@a����I�E�v��j�� ��7B-4��NsN	K.�Y�Z�o��ϵ��gYq@�?���U�u���m�םS�I�Z�"!r�栕�.f3"~�6��D �{�����n�
��`�0.!�͓d�:�^G���Ј��>���K���?p���D��F�ϻ����<`=�rW�@ކpdxLK����AE/I"�m0�����<}7.$s��&�Gw��+>!�ck�ZGo�pt�zX�$�Kh1��?�8
+q���kc��=����;.���c�JI���nK:_����{�JR�^�<����3��C{�_��P'�M[��E���B��d��ҫ\��QE�R!��h�8c���t�$�F�-��7w��Ս2T�s�zL�X�OFA�Ο�H�"���~��.�����P��B�$bs�p[����d�C<����R�%���]�k�zy ����O�{Y@[��,YN���XTt��I�q��pᶑ��	U|�
��a�΁:U͛@�7!5�Kus�Kω庹��������f�W�t+����N��FO2�������x��itL�j0g�O��������1����ǁy�.o��pjA� P��a�8G�9xrZ�X�,��V��É���	n�Ū�v��w���@���h��H# g��(���6�6=1c������v��	w�}]y<��N�(�S-�a��h4R��k~��s��E<��������Q�	ky�]��� �C��|�����Lp�K�X��)�W�V�̗��H�>Ɍ����K(ʯW����	l���v��uPW��/���0�_� ���`�����q;�l@�̄�(��^���*�+�������2�X��Bn!�����0|=�9~XҜ[�Z���9̟ꁇg�U��*��j�}�Q�&���]1� �nn ���pt^۪o��L��+����6V��h��oe[Q��$l�Q$񥒃���4�?�k� �й�dJ�O��+��̀�D�U�\RM��U+K��J�ÉR���{���O���/�f�@��ƽ6@��yb��n�.����l�no�Hr0qR�Z����Z�qr�k{�^����B&
\1�t>8�(���?��W�&Q�MPt'�����f-�9N�#��a4��5ݺet����7�� ���7��S{�M]Q�f�>�w-�`�����X�k��jx��O@T3Ml:�܏}C�=ɍ�a��>�S�����H�T�KE���X|0�
=�"���3 �U�C����@["�ǯ8�mƗV�����š��g��.��:�L��H�B��L�F;H��k��$�; �4�b�s���r���[<V����Z�w�W��"�Bea{��@aײK�w� u��H�hGxQ�o��g̿%2߁�/"�r�����$F�Xw��yFX�^A�8��
/��7�#�0��g@�_[J�8N!w�o}�:Q#�g�>\��<��Qs�a���p�[���⻴�]ny�������Gn�㙭�oN~,�u�MK�)��qY�cx�����|N�9Ξ�߾�1h���!�&l��\C����ƕ��!�U�'�#�8:��W~���	�'���:�Vَ� ���E�SI2�������}�CH/���N,���@�%�H�S���D6�(�����0�d���38Ǻ�o��13��Ea��5�r:��h��H��7��Z�"�ʗ&d=��T�5~���R��>��A����N�gL���[\���,�9;`��b7��nƂ,��D����谫cy��(g����Fq����}��Տ��ゝm�4lObOʽ�f%Jk8Y�}*����I���GP'ch2(_��~F�T2��UP�zC'[[����x�m��c!aJ6-eju�NJ��SK�|�^�����R1Gr;+{�Ϩ��D�	.�|bZ����r��j��� 7i0A0��b}�����j.@}
�s#���N{_�E�*^�zL�U��'L�F �	����h��E	���c���`�G�O�)zu_������~����޾Xpg/�UK&� =�
�Q�(�	k����U��{��R�A��-r���J�\��vS��sJ)z�,�(�Ta��|8�Է4d��ďQ��S a��00����,,�x;�S�:����{���1�'����<D+��J 1��3��+��Nt=�q=}(����l/?���!5��渴E�2�E�K? �\����x�sCD�ye��9��?y�FYܶԛ ���� ��Y���;�9��E�Ig >/
�>���g>?0�/��{�?�P���tѹ�?�mnmB~�;b�X�Nf���٘���T��;?�1��(v�tD5���6���O�} ���	υ2�y$I,⇃D��P��\�$\�B�<��,BӋ��!{Bt]R������t{#У �*s��/��[	���̗:`iw�/X�T���UL��6{I&��|�M��b��	6��:y��g80)3� |ua����P�=�>ӑ��֣�fڮ�ST�D���cX����7G:2��#D�E�	�Ȭ��ɽ�1~=R�8G�\�6�6Zj���lO˫<V��JuUP��M�z܅m5!��M�� /W't_0�[��Kds�d&���E�8�L�#K�!��Yr�n��@=w�$8|���:sHmO�^#��R��\��lp�R^��M'u���u�
�C��v�a}��!?�v{
��yx�%݈<��(!������|�aka��X���s��R�5�OR��p�|g׍��k���.�OL��Z�7^��x y��4�#K�.ږ㰋�y�h(ѧ�g�����]�#�7ˮkJ���6�qO��l
���]��F��[K��5���V�����r,��R$^�*�<�w�R�>�-�G�����)���&K��!t��-N1���]��B0TJב���s�j�Xw�t�=��O����B�".���#㧤?6=L3�{^ ����$(ۥu9�w�Q�/a�tu������#��F�ňAw��,�hVs3��i2�Y(����i��P@&Q�JN��B�6@Y6Jn�P_���4�0B�_4���	��ފR,���A��r��҃�$F�$q�}il���ф)�A���؉�rP���X������[���R`�S���m�Y�6A´��Z;�樸�,�PI��G@2ں}������7�L��`PM�wysʇw����$m��$�x�\S��o��UGBP��yX1���t�x�&2�1C�8zQ��A����&�!(�Y%�Q�&����ό��
�Ԟ ��H��1	��aa���d��^�I�mzG�/ŧ�`]UO1��i�X�rP��6M!t�h?IZU�ׅ0�Y��kգ���9�3Vr�$*M6jE2�b�S�|Ha�?7WA`�\�oD��of*c������֥���l��D+6(���\���x��~�'.q���n��c̖w��2��:��f��^�ݱx�Ncqa"�g��_���-5��z�{�<�5��
�p�����/�~z��4;��އg�p�0�Tͷ�F�_`wh/SCxYSO9�I�T�ڥ�7�e����Ӎ��x�A�����-���!��\�b)�n�d�@L�a��ȉ��d,�8/�1��Pu�DSN��e2�s;o��g0����v�' ./`���w��G����r�_[1�N�qV�3ˤ_�1;��szC$c�._A�б*(?��[��0��Y$3�O�M��K��˧�☲�C�:1Z�8����s>ܯ�gI���/�����xϕ�V%��{�0ǀ=π��U�����5qV�X�<�c��o�xu-�_v���D�߃�ߑ�v����ٵ��	V� 8�\ú>F��uĖ�J��2��h�F�E�������r�.o���V�t�XP�i|����8,e������!�������wѩ�yuN8�;nmz��>J4���YS�v�B�ۚX#<9��*���Iau�,LW�ܱ_��n��
�׭�Ƴ�����P�0�>u?����N$�m�@�u4��y���WgH.H�(���d����lPA1k�nA�[�{,x�Kt/엥����0�|�I��Y�8���X��!�&�����6�bȵ����/k¿\��w�
�q�k�	�}�/�&�.2[X}���=���~��$<`����-@�^��$U 4a��< � ���'�����Ё�s�#[wp!�H^�
�,��A5��u��>;��q<�;�������^�IY�)X�Dg���3g��39�fT�����2��&��X�x��a�[��4#Ͳ|�W �i��w�7\��M�g��-�La��f��6������E��pݬ�J�,=����U&�-�|����*��OH�CF���iB�\���ac{pC��c���_6��q_'�E�����W�T��͂��
2.z�aȰw&e�ݒ�J��hZ"
kw��J�����Z������Go�E�����Ƭ V'���0֥��$!lHz�!��(VIBoP�+�6%L����U��d5��_���ĉ�e�����1HO�R���^nx����TM�3M<4�����=3��j��m,�S���}��
8G���#`<��ז<��p�=�+]�D��:ޚ�A�2��\q�e�BCN�DV�¿�����^�r���}�%Ih!X-?�F���@2�E���7K��Z2��\uO���Ym�;(�,L��ѕk���J���-[V�z#�[�kHKr���l��4�7O\��PP���c��qK�ھN�ְ��>�́/rß6wC��$m�8S���a,��LbUи*���)��ů-S��\��kvǿ���8�Y�i/gMg�>31~�b;η���H��埩���&+���MFҠ�#�r�(oX`>W�k�t�~hň�M�H�p�@��K���2ʭ�t�E^2�K*c� �����T��R=��BNe�>P�0�dHU�����<�>�e�wm	= 7n�-vQ
*�Υ��r0?�DE�-w��@D�}�Z׍��:�
aF�)-궱��*@y3�O��P��Ek�p:�
2uZ��m��p^�0��D�H�V�Xl�^�JWqO����Jԛ�>�՞�)���jo�^h�m_� �X������@�e�CI9��ݙ����~3�KG��G�?���]S�[��Z}�@��S(��GN�O�	�MI4J㨻,!%|������On�n4An �g��!᫑4���-ETEF��+�����L.ԁ£�G}��'�u<\�V�{�����(W��B?���y��%ǆ������j�	j�AUoZ���@�08i��b�W��74i���~@tc#�k��PǱ�E&0J��0������ES[�ǎ
��(���rK��`�cUk��3�V�e+.|�O�C����%��ށ�R���ax�/��nSf y9M/r��8�+��M3��ή�� �J������YS�3�{m��ë�.��sT����U��,DyG"����$��SEǼ��v�	���҉
�:���ീ�s"g�i�K<����pw����i����߂�=�q5��d_�N�l���%N���{Ϋ�X�YI��Nc�.:�i�� �t�^��5�Hδy��2�_��l7O�)�݀t�:�a!��eJ�d��T�I4�5uYO��(� }�ɻ[��0HAy�<����^"�^��0�:va-�|�/�Z̗�'6g��y̽���(�`��K��V������{H7�%ҟ��F��ch4�&Т�o��񮻡�V�=%w���{�e��yn�d�N�dy�5od�zH3@�E}Q�陻�E�s��er�@adqC��ҤN��P6�ʹ5#�#9��BD�c����+G�5�����;4�����lus*w�~��?
�Ŗ\�hS�V�x�܎��XYf�,�ί���E2#㟐�H7kY0%�+�(2���2K�ޑ������\����	#�nE�yz7�z4�=֢pg�j?�
���5��5��O���-�A3:į^ ܃ڢ��#QF�]�	1֖��N�iX��&������O�X���%C��|���m�l�����
��|�[ׄdkJ��oMFz����5��������]%��פ{>���Y<���]o��z��R��6z�g��Nr�ⶪ���,"&(��Z=�`'�m���FWP���>�h<�������~ȹ#ux����v4mUR����"wx�q�L�P��`8�ͬ�84������>*Kik�V¨�|U-4G(�-ߢ�R�7�� W.6/��g�CQ0��c�!0֎D1J�=]��_o��ّQ͢�o!���7��Y��G� 
JT2!���"~���^�]�6-��ѓت�6����k
�K�;U�g�(pUᓓ� ´c��?�8���&ώ߾Ԡ��AS)�� v�mF]���s,�I
�"��w�Ԑ�^��(��d{ ��?l�H����M4J:�l�2'������ w���$���K��Y^�J]�1��X� ڹ�������i�U-��8�1�4%H�+�E�}n�k�4~���_��`C���R���#����X�ZP�I]_�>p{�
U}��H�����N����@�EK�"���s��}Yڍ��H��p�横o[�9��~��[3%�u�M c3Y��f����AO*c��u����(����ެ�SM�����ԙ�A����qȝn�c���jxdO�V��VJ%��_D�}�6�T��������Ϳ�8�i �0w�tS��IZ����B�j�=���s$���
�6/(�PkJ�3B��iO�f'���z�~z\���]L���6Oђ��c�}��|�y;E^������*%���Vˑ�p�u>׀Ln �5�I9�֠Lc�B�Y�Ѹ����b{��fL�㬣���\%�r���{:�g0��"��L����Ѻ���,�9
ş��J��,���U� P�oM�[ ��z�z�p)�L�]��<\O�8s�N�%v#G����ϒ��g�������2�M>׾]���>Ѭ���x6L+U��-k�&ۼO�:���iHhPTU~TZZ��z-�	��j��b]���b�0�/�n�RP�eV�W*\���0V�n:�p,R��_�*�pv��h�N����uU�y�|��ߗ�y�=t@�&*T����V�'ݨ\ݢ+7C��v�~�����_,T�P2+�f ��|{{�mhfh[h.�̱z��P��O8׽��TT�g�Ft�af��*�s�AB����oSiJ��~�R�M�B�7�l|�x���%��l�"��h�����;l@���'&x��Z�;�3����t�}��b���L,�A��v3��q�e�F'�)h�="4�����u�*{P1ng2%'db��z�5�C���z��,b���y��\�%�VuwtEdh�� ��K����������t�-�������ró���'g�� �E�K=q�ɽ�������b��J��Va�D��40�:���O2^�[	��GͿ����ţ>-��A�N$nU���י�|��}�D�xe���Z��.7���t�]�Wsf����T��/�&�g��]c'����ci+�h_0���A�Fl��缼,FZ
R�,�WH"Jp ��J��]Of�rC2Q'ʇ\Ƀl��6��GE�-*1�������I��Y�<�$W�:���i�ҕ���*����wK��
�//�ݢ������:���Z�y��d'꧒,���r�x4K�<�۠�Ώ���<v9*O��D���>"��M���'f�����U��b����	��_���>�k���g�\O�@��c��[��\�9}[
@:4U�Ў�o�g����q3h�Q��ʟE�d�3���M�،�Y�9m�-��Y֤Ϊo�������wy�ڠz�U��}�E�n�s�Ga4�(����h=��sưZI�=�R��Y���>�1��P^�<Y�<.�ً�Yr�2��BJzLyf���EVڊ�\�>m��h^@�'\'� �S{n{-@22w����Rg��F*O�p,�?em��H�X7�e=rPA�=�n�	.6܋XLeq��i�b�+Q/�7^��3����7�~Y�����
)�[�5O���&'�iE�0��KbX#3����}�X�6��@��wē�jy��jʫ��X��&��������ʽ}�0e}mȖ�s��j1p�&|8��=l�q��Ł��NN]����Ӛ WT��_T5�t�����9�]�.|+fg�s$"|��qҴ;=��ڰ RL2Qw�k��8%��k�o<\D�����HM1G�̮c:��|W�2�f�$�b��0�����p3 ���kW�� X\R�&����k��ArŜ�5��-�P�AH������3�,��Td�V`r�{�Y|���ܓE ���*D��l�U�����7�܎{�HE���g���k�^A{����t���a�M�	2�8ǫ��')i7���E^hӟY�������f�glg�a�,�(��i'5c�Ѧ�?�Y+s�rd�L.>'�y@'��N��8e�-X�E7?�A���i��z,�		Z�4|��^��_H�Ǳ�`R�7$�#NH~�X��\I^:��#�CJ�6���k(�T�#��hO�*���;2P|���F�M���930pc����M�~t��I�.74o�"�w�a��Qi=gB��^|>'?�*�rC�\ǣ��
�Q���Ҩ h{�˘�^1w̞[���,��Ni��:�^�3
��2Ug_�E�������FANG���YY�:2�g�Љ[:K|���@��G"�� a=4p35`|\�ƵkRAv�3��l�ZE]�P4E;i��y��X��l�+s(��.&�����nO}�j&��f&i��ş�!��k�v�F9G<<�0�G�����K@Ug@yBPR�	�̨I��݀��Ѫ3hT��;em�7�GI{+��Hӎ!K�f����H6����$���V�@9��IR;�s{/ĕV\F��?�t��}w�,}�r�ƈ�ڕ8���X�M�ê<�p��ܱ��LCgr39�YX��˃ �4���e��_j�n<��;�8��)F*E���v��2$�cR���4nSj�Q&��{��h���
���G^Gzd�P����A��DS�4�E�FxL1�d��@��d��z*�z�0�L����M쭡/a��W�{���>1�������E��^�G�.D"�:���8����u,���G�����6J4�a���R��BH���l�����n/�n m��u�Aކ9>����'v��h��/�d I7�Jrx����!D�<e���,���؝�Ǵ�<!�:���Y���/�b�ҧ��#|!&"�$-�-i�L��y��EA�!8�c��ᙽ�>��X�X�]�jÌ"UHP���eri��߭�}:2hP#�#�@S,3�@�5n��V(�Ҥ$9z���姄��
�x�X�ݢeG{�^������O���@Ǖ�݄�� ��ӱ��~U�ZH��2�ܴI��Q��8����O��H3u�Ċ*��3�6�/����piE�n~���T����},cdCy�ZTz��;/Syxn+h�7I�D^��'�i��^�%�]���S��K��I��%�p��)F���D�Ś��7�}-85fﻌ��v�-_��;�K��HT7�-i��	����FC�����ldz� 6�d���.�P����N[��}�"9N��Ֆwt���0Z�}a�qa��[	���I`�L��Ae��W�yT!T�q�ˌ	r�H������������XGN��׋_�����v�Q59������in�]%��u&\�!2!LsIk���tjUJ;z}�CG��B�/Z�t�+��1��J)�%�q��#�o�/�jԻ���>�Ktj�A3��P�k�k}sR��/�!n�;�I��Ԉu�(�_�M&���=x���F��&����u��R��9*!��>�^��}']G6�U�o�ֆ�|C�ܻ�j�E��@8w����V����W�����{��9��,^����*/[+(�;PCF�=���8j�
�C�r2���~"�����K"�AGOw�/�]m�����q1�C TV���-��
�va`G'�+#��j�T0m��lh/�早ѫ��[�����k%`i�W��X:/���(��
�p���VT��@��4C�c�-�E-Ct\�=lh���I�� <��Rgf�*@?B6N�������G�D��0P�M�O�>�{u��梲����5��5C����ự't��������X8�|�pjs��׻L��u�A"�R��:2�4�58�?Ȧ�bU1 �V���,8�T!�5�Q�N5T���Bi�������C�U3����P���e�<� ��?|�[ i��حk^e�!��>c����=W͞�[�\h�T�[����DC{���>�����o�sc�� ,Sum%u����1m��;@��F�dBN�2��{E|��C]�-�{�zu���F���O���Ȍ.���?g�]cd�DS��3��h>���n��o�ZHb|�!�`��:�ި� �X���4��% e���֪طOcB{�Z�q�e{���h���Lnl�@yP4כU:��i;d����pwX��R0�c
�-���<7�e��ލ�{���VnF��ᄣE[)$LN�NK�/�ΐ-�k�y��=��ۑJ��6�0��Ck��$<aLѮR��n�Ӑ�j����!S�Z��1���~[J�3��Ջ\��0q'�6���XU���?_�.+EI�gN�G��-+�P%��(����N:�3%�J)�$�qz%��ϣ���m���ڋ�20����E~ZW�D��N�E|�7�)���c�u�k�1a���+��AW��aCB�t��!] 3�?+�m8[m��l��I��<��KX�%)�Yѥ�)���'ˢv�2�������IO�4Y�"2c�~�7����L��;�YX
2x�*��6��7v�4-N�S�?�I�f�;+#y�L��21����|���!�m���9,c�������ε���c6�.�.n����|m�9ɞ]3��-�;�8I��_b*��'Dh��y���g��� �1:��y��g�1�+�QSG�8�7��r��0 9�����O��W��
?��z�˝BW	�=){2f$G�"D'_��,ri��6�:~��Ҍv�!<>�Д8s��{aU�x7�"J/�b���� ����ì��i�
`�Y��н����Y�E�z�L)p(&����r�����X�Ҋ�P�m���GI��v��`��DnA��!I�7���_B`m*P����$L�5LLC�/���}lz\�(��V=��Ȅ�:wBL2�S�u}t��x�5�Oؗ��,��
KT !��>�T�C�/�e�)��=��X��!̏p�
��p�B}�x�i�&���Y�m��q8���s�>9��&�?�&�������Y}��^���݀�b�6���Q0������<�MUCZ��鰕��#(8Be<%�[f���)9���	J�aq���1ڰ'��ĺoY_#��Gy�0����+6C\�(\@�e�8B��uϹ�6��<�Y	�0��.���*��A=vc�ݥ�?�%2d"K�:ɮr� �	�b"k ��.U���v�~߃)�$�T�W\��H|�Q�����<�'/Y[fg1� ĺ{8�9+�\���^c20�|`��W�N~]��^��q�'<R�'9�C�Gt������k�}�4�pua�m������G =>�<\���T���-B\��yj��)�?&a^�Nil�a`�e7�J�T���(����wzLN�J�[�@�K*8G8�3�v,:s���>�[�0_��5��ش�f%z�9B�qr+�:6�ko�Y��еH����bg@��������.�ޅ�� ���z�|�M�G
�{�2ѧ��**�ׁ#��h��3� ���#ey*�����a��e�$	&�e����6!h�R�m�isX�ny��@97�XB�
@�s�|JlB���4 
��r;��ӡ5+T���ø/]�R���O)^���U�x'Ke�jc/��t��R��;�f�OD؞����ޟ���Җ��E��9�q�-F���X�����,t�vI;��>�78���~[�g�)���b����kQ#!��O�vS���/R˭bS�/K����yn#��S=}�4��m~��o�A�I��B/��k�6z��6 �A>�#y)�W�t��t��F�M���L1z�<�r]XS3{�0������#r|�'�/��G0ܺ��5P/�5X��Z�NL�1R�R�=%�zt�4�(܈�A���7�x��k2�UT�+rk0����`�Q�4p(/a�/H��u�p����&����!o�����+zz�Xr<��jm�t���G\g����dej,R��4+���G�	Y[���E?��E$)��7������������Q��ʀ�2*��~�Xf
 ,��M����`��Jg)��͉"u�%-�`�/��j>PN|���jl�N�ʲp�/R#�"N���0�{�H�Y����t�LT� �������Fu�~]�����^��K<pm&�Y�c�������o����Ř�1����#����`�\\qGn��p,YU��ȏa�/XZJi�U;"���9�$9�p���N4XaF5FWN��M�se$�����t������A��4���y�Ѧ��=�ݣڀq1�7V�T_e�w	m�z��6�s~%����"�L{�E?M(�$5Z�e7K�DP�C�U�l�@&������]b&��keHq"�!��V����:��a���O���l�V�c�U�U�;��Fp(X�EO���^���L��F�x�O9��G�?&�����Uq��s����9a!ԓ�`���Luȱ�pn�/�U.M���R��/�on��ʅj��f�,���x����Ӡ��fO+n��"��ő�k{lz�H��D��7��� ��q���T�� ��X�!���X\�Dh�l�B��iiD���'օL�ǽ�;��)���d�������EW���7�{���&*��P�%[�X��A$u@9ռ�N�a���D��O�\���
\����x��d�D�'�v;/.�K�a����[+�o��q*7�[�93��(���0���+�Q�Fa~���q��N��h~�!-	c�%�|�ܷC�d���=�>z�Ta�Q�9Ħ+SK�Nׁ��dl8?���h'�`�@��)&C�@��"W�� ���8ȝ6ޭ��"�H�n@v�kC��Ɲޔ�x����Lb,H4`��v�~��/0���Z�'����tr��ML�:\O V�ĝ2����*��Z>̆�!d�}�c�����c�o���o��m�iZ�ݶ�<=�A�=G�)h�#�p���G�&�F��z�/�X��IBY�����9RPz�h4�oNCd�W�E�8�=/�������P����V����ĕ�.�Ύ�E4ɣ�[D�}�]�k'(�Ӧ�u�zD9�{�:�(��z��>2P���*�����o��у���ʸ�����|쒰�l���_X�V�!�
;q�-B��I��)���4��%U��^*���=zխ5w��Z/�[��+ !���#e@�蟅�������ə���h.�����l^_�S�b�c=�k�&	�H��|��w��[w��ܫ[���YGv�r����VA{l���hxm?o�.��a�}��N�%Z|Ǧ��s��I#�y�����.�,
ެ�RF��y���!@25Y�AO(oSצr0NU�1g,^���UYAAaZT1%thH��(`3�-{��j���ʪO�e���j�]2��ʀc���=�2�[W����HLZ�FE|�q[$��o��K��G�a��(�Ľ�L`����Qe ���?���^�
�J�de�΋��3���H�wi%W�]���, _�*���⹦�6�(�T[s@��'��_h�ߟ^�6��rQ��l$��u�t��x���R���r���b�u��:V�JN�NQv��?�
[��wd����k_*����d���M����`��=��ˡ��{ζS�86���wK͗Ճ�S5���f�T�����I�>$w|h�*��K����7U���j	)�L/>M��c��������(΢Od����wc���j�B��;2p��gԂ���]�l^�SzVp
`����q��l�,�mokl!�y�!�����
Y��=��o�z�&�( d}��ࡐ�̦�	,����I�P6�u�F�-� ER.��x�i����y9�fc��h ��=&��D�^�B�ʯk�?��8T
��!�r��	���\o�3n`�&�k5Ď�%��~�<�G�Z=Y){��梇��Hp�=y�S6�/{�x�_���}~mlD��w��8�WFR@��:����r �29n4�ŨUc��®t��DPȯC!,vA��E:�����}���/!)����U)�bE���M������/ܭ�m�,~1�א޷9�&�9_�cn��Kx��=�\�v� ��ⱺ�0)#ˎ��2�,��pY �Zq�����R�]R�)�.�<�Q�䗼���SdŠ='Z??��Y��p3z�V����0�$�7h+q=��D�@Q��C������*	��2���b�3� *�&�}����U4,����	3
����{��q���lχ��"#��ޒ�Y�UmIZ��/�~��nS��O��
�7���{g�a�6��K�bլ ��i&ʮ]�A���ڃC�ڿXD�&?���}L C��+��H�l�*V�3�ʴ8 �b	_�	�M��u|;hW*�Pj�Ŝ�Xd��e��xL5[H4(�ܲt§�78'S���c�/�S�H�� H�+n����2y: 7�����O-��F�,vU�󁁲��")C�q}�0�M)P82"���	/"�k5�}/3s��$���UoRҫ|ۜ�kgQ;p��_�8}6"���u�fF�}��P�����@��H�O��W���>��ׯ�-ܡ;�ϻsJ��r�U��)�U�+w�>��b+\��R���^�s�z4t_@�@���[��1k��*IwW����N�����_���^xvU%�� Vx�^
�j ��$�P����6oa��R�B�3��;�^�V�7��i��蓐r�����P8�?_5�	��~��dH���p�G�q�q����8�[�Ė>�ZR��J�x��>���/��1�W	«��(n�~fJQܨ�pO(H ��(��~]�>�Ҿ���w��?��_�/�z�m�O��)l�K�\��t��$�T�A��}N�4l]h$�\v�j+]}�z�i1 *ZS$��%�SV���Kzۦ�/�(�����*RL�^���m�zd}��e��/^�"G���rLM�����Qb]�s^$7'�B떊��7x��i��Ǹn�V�DK�ح�TR��T�T�v��� ��4W���ęn�B�N{%��'$��F��0̃���7�.��K;rҖ�O�yt	�ҍ
�L�,i�2܁��%L��������"��k�'������y�haG>X���ϧ�*�a3ȳzn���ra�P������c�z��o�����=N;�r����CMg�fN�x���L�$yV��w�c�n/��vey=�}�e�gܵ�ȓ�)�6<���]�,���f#w���v���{z6hu����|^�@�l$�sA���8)��#�
r�M�f�N�f��Z�Mɤk}&O�,X��a�G�c�һ�����߿�'j)����w"��?��ɑXBܨ����O�~��b�pJ��(���44�#�5~�)HׯxA%�f7��xQ�ʺC\�:{���5*��(7c	uDv��r,�^�Eh:5c�4��=
C����|^a�����X*������\(��>�xVp�͡�㹟cWx��o�t>��녍6C�y����2z������`N%�;Q�mf�U�ПYĠ�Y!M��:�a>��@�IFC&��h ]G,�ąV,���0B��}���Y�]e�(�w�Mv�a�F����叴�~�k��@�Ǧ4ڤ��2,�.�Q �����!�
e��r��~�W	�����6Hh�"�)�qa�A��C1�	9[��'�и���֖��:��]�neWs�ߠӬ����tSq����m�}L�SV8�*�ZGJ%�z��q_ʕ7~.M�]Ͷz7��-n��l�c`K��V�i]�)]U�շ!��m�G���ZF�oq̥�R����t���\JNNq�A�/�(�\-3s�z�Ğ�C�X&��D8���"��n�xCc�S�>�V�����|_>X�iHQɩ�~o�T�\���G�_�r2
R~�P	H��I�Lug���	u�<C�Ev]�4�e�Y�LuѼ:�"��[wB��e�k皤�d�a�禑�9:$�k�!�!Ig>�g\�����YVy�ۓ�8�Pf�k	�Az���+�}�P{����qWʏ��j��p(w��'��rr����΄|��IR�Awr���>���p�#�9c۔��,r���Af�:�$1k:2�5RN+�H�n������'���C�˛IN2Z�i����A��*���4@�q�h%YLԥ�������@V�Z�y���I�!���^�����
�CSũ#�Y����6���F�e��ō�G���Qs���<%��ۦҾ� ��=@� �Pч��m��hBmH�+����vw�9B��([fb�S� ����/�F�84�]8��}"��Iȑ/�*9+'Ak^FB��/%N��j��WA��<,��^��Jo��:�G�a���3&��������^-���oR�	9S�e�u:!����*N���,��d@���V�7�2����]��V\�"�s!���~�C�wB'���N��F��?<��f�U�KZE��J�%�6d=2� �T�-D?��vV_{���#��X��[�=o?Y-������{$I��UZX�PF�&8��ܰ����G��b��� D�9��^Ҝ�O�i��PݲY]vKv/8�}����g ��q��Xߠȶ���[�|b���Wu
Wd�N�˞���]Y�jx��������
� �T��.N�{_>�˿q[��5߈S=���	�h�J��	z�N��LJF��H�z���i�)M��{7�7k� ��[on"@1Z�!���}n�V���ݪ�vﮭ��aE����K��.̺�ba�}q���d��,���|�G9�e�q�<��d�*����@KFS�p�{�e�%�d��6񟕯Bd�:����X�RJ;Q� ���8�g ��#W+(/�O���g�[��� �J�ү�OK3V����y�yBj�I/�������o�־����, ELL��,#z�5�[�5�������;�U���Ѥs��abB���ӷJ��Xi�ա$�لP
���b.����i�P�]xd�{j�0��R!��7��D���A"g=�P�c&�����WQ�&>vzDO�>��S��P�/�p)k��m힡L��_��̨��5*W����Fl��%3\��]���G��/��g�Z���������JC�fG]��)���!�F�r�+�T����gV{m�Y$B���C��
	�5>f'��.�݂���qq\=?$���E7���#�p#�mN&|rf9���X���]hv�u��@m�D��4� .��`c�U�]�u�q�W��i�$2n�&��r���h$S�6�s�C14N`nu%������貇"��=꽯�{x���=Gɬ���A6SGB������X�B*]�{E͛^6Ę�n�fUu��q���O��@�����>`?߸�1����d�����"Q��ק{�e�RCac�C1��VK�j�q��w�cU�����ۡO�6-#�:҆Xk&�������z:iL�3Qus�9�=G��h~��s�RLx@|a{�Q�7�����H��Ӄ�K��R�M���?�؃�\ f��<]J��Έ�f�>�c����I�-ý]�ώ����\K�BF��;�pǦ�병D��~W�y$k��d���aD�kUگ�0W��k_6 O�,�]ԕ���������b�DN����ָ]���
��Ů���^|��+k��&${�	�7�@�yJ��u�m�Z�=cQJ��W�7K�����4�/9)I:�#��$�g���O�������GJL][K6���n<�|*jkqk�%{l�ݿ��C��(ܠ�y5��л���jo�3���!�߉�п�j!0	+<1�	��Z���W޼��|���Yg�U�[�A��
���k���	A]�y^�C`o&����=_��}�� ?��f�.}	����Ke���&��@�� ���6��X[�i�
�]��5���u1]D�����y7y���eĂl؏�4cүYn����o�3��.��5�i��C$��h۸j J��9�m0������nW����q��X��Z�U2.�rĺ�~ލ�U[��P.��L ;K�x�t�ٓ�������� s��[��c��{��"x�+��Q� ��굦RT(T���v[�%qC�Q:|��u���>����5l	�ĒeQ�"�[�R��(�޿�+�V�_t�5|���Ax���4��pRe9���F��^��~4CfW��f�W1z(�4Nb$��(�*L*�Ჟ,���Z�X��ѯ��G���cU\�G/Y�E����0��)D34'&|��i3�:���jj�\������J������9�[�ۖ\�n�/$����4���=L�	G��������~����`1;sY\9GHr`7�J8�|wGU�2�zW��őe�nA�Aݍ."ܜ6Z%�V�G/YI�I���]Im�?����#;^jN�Y��i��4(iOх��B�R�K]Qf��x�78�
�����|�"���sʊ5�^�=�;Q0:�����\�-|s�i�-p���k��~S�X���Sc$��xD������h��T�2�g���@�?k��:�����,�͉̋���*-W��,��������,��y5���x?B/T��M��	�B��;$��D&���G���Q��5u��+ԑ #��*V�Vj�rp6���O��N|KV�����'$�ߧ �Hz}�m�2 ��%��� ��(��A*��g@�-m�`�?ҋ�q�I>���ٜ�F0g(w��:ǃNv��OQ��^>Zԭ_���۫��ݕ�a1�� `�ܜ�V�^�[���2�U��$Jׂ�M�6�aj@���b|໳���!��>m����s���D��%ܦ&�Q�]ۇV]�z�=���jt:0z�ϟT @�>S`��d�UP�D�6I�I SU��[K�ޜhQ ��������v�Ė�ÿ�{�NS�?�i�E�8�+� s��b�d��05��=�!g?�����$՛cS2;�3-�H��0qM��{�Yh��$���l�<ݔ�T��?s���Tf-'s�E��rp�ns_�u����:�[�:${�%kP[�ש6��/�NS\�LD.�ZUb�ŏ꠲���Gz�[��b{ĉ)P�!�BD�C{\J{���4��g7V�������r��*����5�N ���D�h��n�w��ӭ�D����u[�H���S�_�0>�tQ�i��,��Y4o`1����:����Bh�֖j��T4p{��C�t�a�/��Z��J.��\�i_�2B�\�7��)��g�Xv �.���
�]�����r�/(����Y���� �PWS��׃L����Z2r3�0`�~3�sl�6�2��q�F��18����L >���q�BT".����oF�*Lr��L��J_~5�a�8bv�Qj.��U�&�� !�P8ŜT����ڢ;ݹ��k˨'UY���M�}��b]����]�RfnBy0�ު� �m�1������c��[��w&}`{�c�#|�<8k'롔4�C��.�N-aA�/Q�{{�A�Cg@0$��`'������V�V��r���~r�����-�����Z`��\A� Ύe>�͔a�cٓ��R�l��5�.E�4s�>�baSa�E��9���@� !M�0�D��@���s�yz���m��I(����ڵ�S�>���8N࣑��Ƒ���ZO2��W���N>���.k���W��jd���犝���e�-=U? ���F�	��X�(M����P3v�ǻ<��\��{�\(���j ��a24���k��0�Dv�e8�h��])��m��~�&;Æw.���a�2�v��x��}
�ǿ��P�F��<��$�2�jbM4����NL!��*R	���|Y����"�q���ײ�=�O �3 ��6�uN���˗܊�����U�{������������:Q%ۤqU�N�
K�*����d��z�ꡥ��D։Ѥ���-<G�Ղ����]�}^.��0[wy��6Xi�%�Ю�t��!���}��p�F�<DN޻�I�����j9�dD�J�:h�pC8���X�#1� ����ghD�~�W�1䛏͛ӭ����`r�����3��D�� �o�F8]��q����\�>պ��N����]��EZ���	@FF�iTոlx6�������֣��������<WTؿ�4<b�x��I%L���Q|ƎX�hP��O�rY��tT��}E�ѧ���:ڒ��0�#����6/?�h��C�~Դ��P�{�=Pk.~1��aK�x���k�R�[�{(�{����e^��m���>54��]Z����k��iV�k�aý���T+Y�&�)�.��M�L�s�,��p��]��)q��*e=J���j��j�Չ�"�n(�p�������1�;T��L���vT�dBrJFƿع����H��v��;Uת��V��8;�:���� ��
{Fǋ�������9F�b�@�+b����m�Q�adT��ztr/��ܤ���^��'���=�4+�
�H_kYg{ΌC{�{��	�)#�M����!\!ݻ\�jhI���)7�
�W�U�m�г��KHS	H ��Iq\M�b�"7����bkz����;.F�Vx�%p��R��y��M�ٴHMf.�v�S`̭9����%*1��5���U�Hp��+b�>�j�qt
��!�&CuJ6�kg�O�����!1ѻ�/�e�Յ�^m�9K76H��Ʀ�A�3-ڜQ�g�>Jb�]��!1��Z΢�~��L�����j)쏚aiqd:��a2c(�8Coz��
���O���Et~U>[���2tW�)`����Գ鬌�+	��b�b�6�������V×C¢r�8�8���)�ۆ��X ��l��kȜFja�:��B�	X?�Dpۋ���u%�6>^Ҿ46O'X92��[d]�2r��f�6�Ҏ������>>a*�w����6)²'g��5�e]񪴛��dm�9��k�lODg�Ҭ�W4!R~�$R|�E+Dt�����XQ��5!W+���H�8�ɹ{�aTt3��&#O��8���q-F[�o��&�O���ڈ1����䫘S�̮hF���°d�L$Q\�3�E�P.Ϯ\x��#<�I0��oE�f.\����������p�;�ɟ��H� D3��T$��r����>(c��A���촆J\�.��!�a�ӫ��3Z��F���DP�*�>-�^0�5<���R�@ݏ�� }��x��wG!4�
��Bx�o�/w�Wş�Z;�i�����ӧt��4�hʍ�g>��Q��E�H=��E?��l�=m�581wG.z�D|J��0� 5HD:��Wt~�ՃO*Y>q[�u��=���]�'�P�s�������4]J)4�G��#��т@� �C'AAAN4�bg�� ������$��7�8��6�{��G�6�֦�F���p/Xuߥ�M�0�賯�EF����S8�A�(�c�F0@���}Iwm������oq�����ꉙo-5P�g�I)�2�N�b���]�6���̃�I�����d��9��<Ȓ�EҝAcj�K<6���Y1��ʮo�f"*�1tQX�I��H>W�Ox�γ(v^��ȃڄW�ܭ#�
A���KgA��חV��A	�` �lQ����h�u(uh�KI��	�[�z��d�eF����)8������N�֣wlvNbu��++�}٢�����%ظ��{�\�wH���Z��,�ǉX,]���/ӓ�s1
^���iH�| o�s�7�UWV,����31�`�܂_��>(9 l\����~y�;�yf�	�
؟�"x�7�zW�,�l�x~h'/;�O�)��f�J�F����_u[�´6�<}��sJ�u�k��$D�?����3���s?f�TlޭxD�J���h:㨣}��?Z����#��|�!]�M�[���ŏ�0��+L���K8�sߖ;CJ�P�olv'C�8T�2ο?�� w`��ήo�>���L��T�-�V̄�x�f�����^��&舨}�ߴ���aY�nfE��L3*K�B�Rud������|����	��'��Rs����Ŕ&
��i���m��&�������D�q��^�KX9�'Em�Fmf*S�5
	��|�-= Jlq0c;b�3������hPI�BP)O�E�_�AI��D�T>V%y;���g�L6MF����1QDX��:�`x(T��I�4kf�(�Vb^zQv��WڇM+� �|	7�i�B��7�Vjo�9����x�F�m�pOS��WSq�/�Op����Y�U��\�;�i�?s���י'��qD��l%"JeM�!7���Z�pBw��d��>�H)�"<�����/�@f+�M.'��0��D?ՑT� ��"����}�3��4ڃHr��I�.g��	 ZNK��q�jMX�i�RV3 ���`$��5L�"p�d������Ɓį.'K:�eY��;$�z
mk���0�U�۾s2@�쫖n^n�<��Vx��ٰ�G��)iX�=jui�^c���:�p����y���-�FH�)��g��-p��\�	�gm��(��d��t�1�]��JAv����u���:f|S�����T��<��G���P�c>�
a�5X{\oPޗ�T%jN�G�����u�좶��=+��yH�#�o_ıeQ��=F�%<0��r��2��e����V������w�?��O�V�խ�X�:�vJyfjuQQ���~�I����'5��p���2�i@rn|<��Q��Ӝ�K��#/�f&��^����3�9�34&r��[0{�w;��Ͳ�}��<8������|v-�پu��!�6�X�)Ll��<EQ ��c=�U���,7�p�![�����(ǳ�q���=�$n�2<��F.R��r,DA�2�I��f����.Y�[�90/mt��x�|���Y�RX'Q�J����`#L�z��Z�
����Տ��d��}���j޿ ����4��Lk+ �Bu{ae]L��0qUq7��7�?�mb���v��Ek�]S6�kt�~g�u�`s1̨�+�[T�_9����zEXW��c��>8�
;�R�W�'r��n�<Ĉ�].�ͯ�)X��?Lt������	�v�~��y �K����i������2��zw#�pb���1]�1\r�B���"�����JP_(�>v6�����HM��"�U/<�Zi ��Ʒُ��\q7	f7]�٦���Թ���{=4����_^}u�~��`�W��'�r�ap�H�,UU:�^��%r��j����ijc�^eT,Q���3����m�>ɻ}�)����7[o7�~��E� '{��<����C7�`��?8�H�G&#2[܋�Q/���[܆؜z94K�w>�dr.���aЉ�0)j�� �]1�u���ǰ @	���`�=�Q����UF�	y�sLE���MCu�bQڡ��y�y�y����7��`ɳ�Ρ^a���~W�Dv~�����t�o�A�3ܐ쐔F��G�Aؠ;��)���W���_mh��@���� 6\���%��|T��H�B�&ο	J����t�e$i�H]9X417�7�t�~ԑ���t� ��I8�J�^|�]����#�h�z[��<�����E��6��T�� �:b_D���*����+Kbɽ��bl����Pfi��"��_�"l;T�~FCB�"�b;�&�7��4^,���߳J���*���@F�!�w�9T�il�Ñ|����R|�̇E���'k��x�V�\|��>F��6�,> �ׅ 9QxѣQ�b�G>�ލ�;!P�b�:���/�D�����9j�����x�Q�km>6n!�>l����?��T]˥#�(�ӭk�E,H=\<&E"�i���6H��xB5����Pe���a�v�#��e�x�9O���lDE$��m�y�P�q9ʗ����Uk��J�KJ�ln[��,����|�m�@���CW���)�k���h�-$��~_Dp�w��F���ô�� �-�6#���	��Ŀ1E�$��(����r�}Ob����Vs��2X��"o#k=���R�Z}E��=��J������W�����Cd�蘰5n-��VIiR��[��-�����G揲�h�'*��]��"6�)��N�t��r�f����#�Z�)�o{K�������߅��e�	6���+<��j���{��h�/�1��;��z[X6�v����aq���W2��Q�.}�5{vdl؇�z�
*bs �4V�vYX��HC8��� SM�VV�:qM�gJ��3��=nq�!C��UL��� �""��s���x/�/Кg|6�>���aC���g��iD~+�"T���op`�%�m�RݰB�R/HV>�Ϝ��ڪ�vS��@��q��c,k4$����ۂ�Ra	zL�&���$��,/:.�9��!ぶ;4�s��r�z�̠K�9���Z̗<�s�}��ʇ>$�9�޳"��9�*��*�)�1{�1k~�+��]'�6�Yl�������l