��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i �ZҋY�i�y�l��ԕ;D�e&:����ɕ�ع���^X��e?�h�>h�Av�"(�ݐG!�^��b����l�W���;�yoZ�߅���̑)�P��g��%Ru�lI��x�	7����>O�;�؀X�D�խ�8��"�h�I邛���Za+lo�q1g,� 6}�k�%��Z�4^O�a`D�M!��VB�K\J=#�����H_�����'��1ET�O6�¥����[�y�E\7�����myIB���"i�E9DS��=&�r��ϓs�I��l��ۭf�*���w�����l����n&�k�e�J"�;l%NY��,�� ⊗]dCX���������k�;$-�%��au�Z��&X�*zh+З�8����o�gh�횶gE�"�f��ߌ�\��ں�Sr1�nG��MM*�QI,��I	���Ra���=���W4q�O���H�/]�:h�O:<�y;7P^.#g�?�us)D��&�(��,W�������=����וs��6�破��g�@�~%�h|�z���nJMI��h����5J�4:o$bh�����ʸ^S�������vߔn��Zj�P��M�^bdaT�����q��8�}�������������M��0��[o��r��KWP��d�逦U����s,�����J��e��7Ȑ���#�U�e�Ia��}DJ6�B)�\u��o�`��@TG:FB�s�lu~�����%��Z��\/خ���m��L�����]u�L���S\C�
bd���-�l���Jg���\�3��
.�Cbh���c���������]���1Z)\X�ACO�n\���X�&������\E��/.M������4` ^J�I��5�1����_t�1��,`�$e�J\��P�R��NQ�H����l�"U�I�3����(1�����^B���+Ҩ��X��!$9,r�i��|�[V7>�8���)h��f�ejo
 ���e�TO�si=4��/���_�4�ړ���U�|LZ��y-���`4+L���5�'�m�n2!�k=�:ę'�����$%�L�gI4[�1���(-vJ��!EM~�"D|��Į�q��$�z���:Z�i���䷳���`>����Ɉk�Uߓ�D[Ҷ,��Ê��;���#�rMw*ܪ|8)�5�0�K!�G,��4�Υ2\И|Y�Ⰼ�y������Є��y�[*D�N;�������d�u�}�����n19�k)0$u7l�0�+�홥��^���3�u��؀�dQqw����oI��z8BVh�#��<\}��R������,����!�q��_���ʩg�����N�������lɎW)�5PC3�ї/�������I%D���_����H��ڣ��.���V���#��m�h��-��?�>��i�q(/Y�+~Ѱ�܆<O��L/�h3d�B���ƴ&���^�������%?V����b@$QSH��n7�Ȗ��"��h�(�Ңd��^�:A���ci��D���K%W�x8S�]6o|�yԒ���g曈.�p�u	�O(ּ>7P|������=�i��*`�`�J�*5�<Y5/��%�K9X�_u�� 4E_���841��E�%����=u�ݙ��W��qދ��J��(�P��}���m����]�x�˭f>�����}�Gu!�Z|�U���#4"s�_��$���2���F�$c�x��gױ�l�L��*VN�q��)Y�I�c� �ۿ�{�I�`�=n.�a�}u�
�ߑ���Ʒ��ν-A4��p(Ov�6M�ʶ����O�-�NÕ��VZBGf��ܭc�?ZԵnn���g�������pK�-S!�G�h�(�$�ht��p�l_��٦ɮ��J1}�E*	2W���)iP�]��$�˽����a���ۨ��F��n
��g�N�-B��ED�R_��z�����:��9�v����"�Q#m)�h>��C_���X~�%��M�Z#��R��p�nZ"?�S�1���׵ik:��,Mb�F^��>�ք�F�/�u�o��U'��̲gR0�l˻t��.��]��Z� ,��uY+�
�m���#јuK�w���;�/䋛��k�a�*�����.��2�X�_,�K?�/�v:?�n��W;�ko���<A�����&5.̃ė��sԂ�����_*G��Z���13zGk �ٰ6?&��{w,���`Chp�4K�5�ȡ��s���R{U$��U5��ۢT\�Ԓ:��,?�V m��M���ʾ��vM�2akM\��he��T�� ��)�&��r�����V�`�廴����	�9��Ò�+�ݫlr��f������p�����.^�f�fG.����^�匆�g"|v(�<���e�?�`q�}�#
<|��"T�d����/�A�wI���W�\_n�dZl�g��k�RݍFby` =YĐe��
C$����2��1��/g^��WO��AW�>�*Y�Ys�6�=���
�jt���_�k��Dk+z��y���j��s���&f��NBپ<M�� �J'd�
��(iB����^��}>�!��	G�G�ɻUX��^ԩ�}�ƾ���S���C�����C�	x�

��Bu2�5��<'n��ax��,xxN~�5V@^x��F��Ui���{M���í�z+1*�����_��ȸ�ޢ���9+&�1���{ڏ��$P�2��J���Wӈ��Ez�&��#ey�)^r��SVqRql%�l`3o�a�� 83~�=B�E{)D�56�H�W�ӎ�X9��!�|�o4vc^�	�T�ÚU0�����]X�ۢ��֚R��E��|��Ɏ��N��&0�Z;�ⶒ�ue&Q~I�3�W�+T�P %Y�-�҆�ڤ���f�_����F�>�6n2�7R��IU�97��[勲ݳ�
��N*�~] �n�¥.�xr��������'��v#�p�tԿ���$�����b�L��~�:f�=M�r@��[�V�#ڻ04P��韱FB~�