��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�2&o�~xݰ�:�}�BUO�x�BʣA=�S�^<�໢��~��`��e��m��R��)���b�W!��~��_O\D)�M��#��验%�Ye��W)���>��<���m���dh�%�(�9�U�ܜ޷S'��w
�����A�X��jz�� �`w�sg]���Q�<�V�ɰ�����9U�gF�Ş��$�aH��JqW����{2e�P+���{u�D�^NO�:
�=���jڣ�)�:���YQ� J�|!�͐;G[JĠ�{�1��Eh$4����`�xp]�p*]���:�P�)��?֓m�q����HZ͔�=z�ֵSĤ� K�*��	�����Ҳ�:��t��c�zs���ܲX����2�-��q��|���������9�Q�W簡̟pK���WM�N�Nf�>� ��b���S��� �Tʽ2b��S�d����p��rp�r�Q�B��sx��'�������A&U7��2��(y�B<:��r�pfTOXw����.QC�AC]�`�\��A��r~�gc��)(�K���YdgJk8���M&]0��fߦ��f�)�[L:��[ƶ4����l��/b��x*b��yﾖtTq���
� W�D	iJ�L!��J���7�s�̠gfr���J3�ڮ���a2��{)F庺l`������������O�DT�'�	"�?89��)���t1��u��T�qw�>%�]"~`�M��ʜa�0 �0|��q�25}Y&���C���Ni��v�N�On�R�@�rkKgu %n!>m�2���"�g��ӹ�Z�Z���j��/☐� "�K���Ѥ{���`�ϙChGl���+ʨהY��$$���&�3}�ٱZ@�_�uM�y�h
ߝ�v����媄=}=�/Jx�˪��h�H��墢Jv�B3�)����^���\������*#k�.x�0_�k��pXwZ�[�����kQ�:���M��#� 5�������c��{!����zIg�L1� �w������ce�J
��^BJ���#�[����vᘀ~�N�dHfO����ڽh|퉔RnW^�A3�4K �0�^aNXt�
�]���y���[|��:"tyj�5��h���(M�փ�*a��5>��|!*�5����]+�'R�a�')���T)x�Qa�@b�D-EZ�����{f��E+����>���hp��\6�q\�Q����-�D�yr�+%�c1��v�OX��vbN1���Ы�ymߧ/W..��A�MQ�(�RF�͗K�%����|��⠵���r8�Y)�⠙�C��+��; sI�dl��#�|W^��f1πi�f���}��Rh��K��j�]�0����Q�$���g$��`U]�M<!Sܾ��'h� �qqPmA��&���<�}��z�m�x {Ŕ6 �r�ToOV��n���dfҺ�n�:��R��B�N��~(��^������i KM�����xT�C�X�@�d�!\� �`�`�Tp:w m���O��x�VPh,�-��ȺlR�}��-��޵#�� �"�����ъ�*9���T��-jĤ`��3i���__gNg�g��j�z6�#G�[��+���N��I��t��?��Y0Vu|�,Qi�);�Ul����ND+&h,F�B��Mܵ���2�H��A�.e
f��	ы�PxZhĥ&h��Y+X(�Е�U�W��ƿb+]v��vimӈ��3�*>�	O$9�,5��m�5�g���1��]ٟ�X20���f~T�%�H��⌠�Ѧx�.Z�M�/�)��Jj���wF��{�	)�-�G+��\=}��z_ ��(Y+{�4T���7.�!����:��r=�ۨ�YLP`>�DK�c�ǩ�/�т�`�e�IPxxrC�G�j�wIVe+�\L��c�<�;��b����aA.��)�{�C�㾚���;g���]% �M������E
�9,ץ9U��E2�v�5���_Ƌ>>���������Z�o�-�`���4N_�Q1����������z��D���� dWDG_�	;�%��G7�fT����|��H�__�Q�:�a˯�O>R-p����n����` BE�b��h��i�ǦGܔ��ڀa��P4�#�'�f��O�6"ye�s�Ҳ`>��������"�LҀ�
�)���#
ȭ���&��M8�ܠ�Ax|M����K��K�R@�z��/�!��GC�ĔX�AwPg�xw���oà!�<k�c�VG�e*<^������A�X<E�}���؞��^�3�7@`7R�F{޵ô��Ɖ+��2R��a/�kih���Ҥ�ԏX�0Έ�	!�[;���h��IVp5��������Uχ���w�J!����CD�L�n8=�����]~�N-d�ѷq]���Yp����>MZO	tp�8�g@����|vƜ����`f��eZ�Q��>��3*0�v�d�PD����}Ǐt,��� 2��H�����姤,U��S�ϿH�JO�.�k��a����ɉ��5�.�|?�2��FRK�A�.5W>i��y�J��Y��N�x�8�v�S�-�ޮ�U5��6��ZQ^0�à��X�ͺ����,vE��j�p8a'�d�D	BF��G��E��AA���\}D߾9�����q����������-�����!)�'��7�g��eמh*�,�T"�,ZR�|��E΅c�S ����W�RCG�>�~���aFÉ[��W�t$�z��.pe�Gr�2�~0�����]�ފ��JƆ�P��SJ�T��;e����W:,IM��!ʛ��o�.X Ȩ��P�{�W����L��������s+�7v�$�W؃��h��E�� (�Z,��U>��͹5Q&��+&g�w̦�NK���H���ށ�b��)�+ ���v���,Yb��B=\���J@´1��ժ�y��d�?��tԧ��l%{I򞃵_��%� �?*g<w��џ�B���}�Q����ʸ�����v��$*��5��<�]x��lN��H�=�Uʘ,�y��[�d)hB+��zf�R:�B]p��G]ǧ�!'�z�z�+�-�<wWt�Zw������K�綎�����	��k(�?@�Fzg����{.�+6�Aj��b��9�~�]z!(�\���vE��IZ����/s�5���ړ��)�H�����{;���Z��yl�� �̻voYBhڸ+��W�Nh懲��UF3DHWԑ�h��J_Ŏ1�ٍG�6��}�_&[�nz{d����{v�=���X����q�Cg-W� �� �����\���@"1���p���~�\����k�f��F���资%P�w?ٲ*��g��z��b��*y�0N]�(��ZhT>� ̼�Z�}�)NA-@v���E�}en����d5_,P B{]��<�_O|�S���h�!��"a83z�H����G���g��NIԕ6E}�x��[/��S�')|M������/���b�L8Jk��!9@��?�]O^�rVW��Xj�fA�l��t�BV��I�$ڏ)�-���VT�OV��Y4�Zi:�$���_�	�נ`L��v�䓩�+���R�6/>�<�&Ѻ��\.��ӧ��dH��")��Sצ�S� �A��b;�EN�%�P�^:Ht���8�i�1kО��rT�>�U�Go��q(5��ZC���з���������	y��V�1����(�6,�R�����{�*?������0�>AZ@V�d�\*N���`2BO���y��x�ͮ���=�$
[����8փa/�6��!	v�&�rVa��w�!4�F����;�d+']d�6�{_��	�%7�>���`��O_3�g,�<a��Y|�G�8����H�e�G������v��V��#�W�2F>W���T�4�����ɘf2xn�1ח~Ը�\��_�I��1���y�@��=�0�`��yy�J�ؽl�7#�&_/u�RA7岕mϛ���a�Ƶ�8Y���E��// ��X߷\�o�ح��''@nAEA��J���r�!l�HoԮ�1�CaQ�9�V�8%��+���<���ȘVL���<QX����q]�׿#,�OIe�h�e������!~h�|�ݯ7�׵g���U�?5����/u�x�j�`>��}+�1�����Ӷ5����[�ʡ�_n��(��C2g�|�MG��8�r�F{�LKD�(pp�����ps$�)�Q��".�1��1���v���B���RԦ������m�M	]-d\K=����
��k�4I��󽊴����%�Ry�7]��<s�o���B'�M�P{,�G�I=�q��ƍf��W�`{D�)ﳪI���<}ÁrJ����ęΒW
��3�U��E�H�a�4��T ��D즉��W�}m~7P���x�� :Ӥ��O���K�nJ�
�~s\+�(��X��YI��v��
�F)�P����PA@Q��A��~�����ҩ)��{�rr�
�.���I�!�ˉ�c�m���.��`���+�l�i����_@�X4�G
NK؉O9#���j���Gy/��zh�����`�S�l��<��O�^���\����N��C�r$����z��KT�Z�|}$���2�q��}����J��n��q��<"�Šr
��l?>�A�.�y���B�{4ç�m������0������P�d�A�Zm=��V �	Nt�z��N^ek�5�(H���b���źQh�)&{�w�aa�C[v�ث�O�͟ �q��*�����~���3�;1c1���D**���8�g����(+������=}P�L��=@s��R�E��^ꃯ�Rc5�ِ�<[o��ih�6Y�Oi7��>䶊� ��%�.�8���8����J�b�׹��/�m����d]�[<��Z=X�4$ZI��|�8�}��~i4�<a>B�j����}����̋M��4ێ�ݯ[�k5V�6���]��)) U�H�*D�F%������j!��P-l���H���d�{6�X�|����o����/3ʤ���Ö�+!Cp�m޸���ͣ�.�|���9/�v5�֛b���>t��ܔ9d}�h�P��G���G����I�J���>������]�d� ����=��}�d�۱�T ƿ�;ɠ�p�Ϳ���>gB;�!$.s\�8Ȕ���xh�aA��nЇ_ϜAڡ��](���6��W�QL�B�3��O�Z������Ct��݉���G���1w�4�F�d^>�]9��LN	H*B�~0� Y�,*�?�}P1��ώ�����{�ǺN�Eѵ� �{ ��(Oa.� �S�aY�|��l���bH�b^�,@�$�Cv4ݢ�xc9hd�Q$Y썣�|ؑ�Rݜ@��fd��+L�P,������~G���}�|^Qo��T�oK��?�14)�r�\Y9^Y�Aׂ�2t�CJ�>L2���F0'�wY��0/��X!Z#1�^x�'Np?�D��J��<lO����o6�i򝭊:����.�C�ZQ�<^��IH
�EꇝZ�Հxu� �籞Y����p�=�Da"�x�)'l`��)�&��01m$)�mw��~��?�%_��u�!ub�Ȕ�*�fq��uo2�|����y�Mfs��^�����U>�٠'g���h�O&���㼾���J���9[{�4��n-��}���2�	���a5�D�$2h����v��y5R!hX#'$�9N�P`
�6�'	(?�����[�h��$��]��Y��H0S|�9r7���� ��BD��-4���L�p(�XQ�:�� ���7�~���b&���46a�q���>�9�r�F�B0\�B@3Nz�e!��5��q��&~���z/��@/��и�%�)H�*$>Y8�Ҕm�q�RK��Yi�ٗ+���s����=�ov�����!2�̪^/��&��|m�����{lV���~�
i��Hi�-�ϖ�t�(�B�	;H�)�"��#L�n��۳�Kg��b5�u���KGu��S�d�#b�i$��E��c_�^�j�Rc���WS�1Pu��"<<��	�b��V�9��_=wm�Lޣ�:������O�V��8<x�%O&�̡(ʤ��POGS�y�rS]������੍�y�c<6Y�E�R��p����5{�y L�ǀ� �� u��Ͳ*@m��P�\᪓~� �㥿�������7��/
+�M8����w�x{�����®Ѩ��36=8ml�W�
jkC�%wx|����Y!�ȋC���|��=��-mO����R���=T{�pv�3u�r�8����}��#����^��n�e��Ə��wGl�ᎊ���#O���'�Ra4!
+d-��G���g�{	�gzk�v�B0Bl=]fhP�d(h�{:����P(�x���]խ���,m�臱��'��8�� b�#{8m�yo#E���QH�qv>df�B��8i���n�AS.1'�5�H2�l��2��W,'����jپ�U�BN��j�U�!��&��hd8�����D�X�S_պ�^�;��O4����n��v}EԃJ �ab���:��?�VdBl��x��G�N��k�����w�ǉN���C���f�l`��gY�RF����k�6:H�M��h��H-�6���9�a�T��)�0X�#	��&!�1���F?���}�O4y�Q.��J��IY��m�22m�}QZ.nP�**���C]C�Y	zE\��r���r�F���@�/n` �o���¦1���(�+����-3�n�� �;�Y�)~}�?�*����G@�g�*�7�d�	U��u�ӃW��ye��bOQN�<�ʏ~��X���GN%�'�\(�>�@�����D6x��Q�.��>ݶI���1{l?e���ƚ鐬q::����¸mGavF�F-��r�2z��G�tH՜���(E��fa�����	n�cr�i�,\!7.��"��9�(� �V�b�xҜ̶���щ�
N�1�0�(/ri�S:,�0��s�)DzKM��~0h�	��� ʧ#�W�f��&h&4���R$YU�!EI�jV_-��� �Sלk�P�~7 �̀�ĺ��w���FO��'��T^�u��
׊��g����K�I�ގj��&oނ��) ��)+$]�����*$�\�ڂh9�`��J��)�8�m��ЇFTU���hCK2�@	-��\��À�1Z��.X���@�RїX�r�~Þ�b*w
���^�.�逹t]=���q@1����l!��G���`}x�6k�')�I'm��������{3�D��;yY��G��V���<��4V��mf�T��_�H5�b*F2sz���:b�nj���q�mw�R��՜m��ھ�O��L����MH��H�.H�	x.�>���֋��"���*��k�n�0�1�)���`XW�T�S�[א`Y�;Y�;�yi�uo1�����7	�����,�-fu�L��Gٓ����	0�9r�H�'&�I����Rfd�G�G����L ���0���{�ѷt�P2d�\� �e����h
��L��{ʕ��u}+Ś��@>$�^��x,�Ir�ǿ��P+�,w�\}��=����wֈ=E.,�$��?v��l��l�}R�*�%=`Dd�*���=*��|��+��r�a_ͳ�k���F	ûؠ��3kt(=�d�X���E�|s��|�W$������^��zr��:��Y k[.e6�)o�Op`HfA8���߾)�s`I-m��o���ʹ�fp���Ź�`��y���ňs�-���C�����kz��(%���_�[���ȏ�f}ޏI��e��
`ZIsBJ���8m�0I*����2�j��gdk}=�Z �^9�~�4�T}���Qjߖ���-�~`�|�'V�p�AFOQ���ʶT���\�]>����;�ϤѮ��D��Y�!�Ϙ-��B�4�T�A?�F�p0��+"�D�y��:ٓL[b�*Mۆ���;�$�ΧX����5��#���q�c�%����+��o�.�`����ƒ1Wny��A� DT=�:F�Ø���b��v�" ��9�'{�B#��qh�I{�Z�s!��6��E�C�� ��(�jĪ�\U�����i3z+C� }�t�����7�����^����rGТϻ����n��j���L!��J�@�Al&�F��h�L��a��4����NNs.�s���b;k=W4�8��=��g�vVv���n}�lGةh�0�D�MH�2`1嵽%�C���䳤I>>pQ�_b�8x��ս���r�^Ou����C3��9���	&�i�Yތ���l�3�ꌧ`-�V�;xC��m�0NK���Ab�1�I�~J��|՗̒�p�d�i�;]�qI�@ńV֯�d8��rnN��͚|��~���Xg�FC��gvb�p)P��l�V�Tk9�5l��b��_ f� '	���������3�N���a�v��;c��A¾�m+��*>d�7Øm�a�$�����fo�����O4�{����q^�>��唿V�(|!��KG�����;��z��0*i���oM{M*�ugh%Lť�÷lJ���vV��I�<@����A�N�۠iN	�<�]B����dqq���i�/)��Z��R��4������-�6Jd����ߝPNy�˼�Gr(Nٌ	�8��+���i�ͮc�ݺG�/�7 �CpHe�e��kTS�Z��[M]Q�)�rL���/��7�4'�sl��i��ެ�8͙E���{<A�BW��`D��4}�4R��E�b0��5�5�e��K͇���F���a-��6��]c�VH��s�8V|) ʍ��t4gߠ虬>6�n����"���a��%��~dZ"|���աc���7 �t�9	ܝ{�������K�1P����kf�\���swɜ^Í��"Ǹ��>�	�nĠ�H���/��0^'e�e��ٿk���0��W��m�s�#�P��J�]�?� ��lBKeDN8�*c�:%��|vT6V��a���z��P�z`���a]�R�P�xӼ\E�-���YXd�!���Lؔ���T�lMy�ğuke;�C*D\��D�� �#�&F�Ir`_�k�f�Nx_�"����O�_�q���'��ĜN�^�q�P}a�D�dQ���sIA����'�h���O�V�Yө�	E�1M����@��Q-�>�����"�!Ý`KE��ֽ���>LU�4&�_`Â�	�yq�u���>���SCD�FEx&lhz���������� 1�i�V{�r��Q�GW�ف��B�x��|��َ�6��Œ.�'�[K]kC�{�4��b��@��uT��d	 4��Tl�=�:8��""*�����.J�99�pc�ad�GoՃ�MsqN��J�R��)�b�wϢ��?e���C�ˈB٣���ki!ev�c�$���^M�Ǣ���e�Y�w1¸#�g�7��~�qZ�
d�0��P�]�[GX���R��P��:1�z�j���d����
Q�A 6��g1����)�N����J)������Sߋp��<�gߚ�D4$Z��u�}&��ci��j�bl7/�Rl����7��GͲ��%+�=&-i˿"���J��U�h�t��y=�ũ�l�;�E�%���E��=�:�
�\�(�
�ڔL�
�w�ԑ�LFgw���q?���1�&�+��$�x')��N�R(,�'u�D־��=�\F�r|�E~��0��ƅ���U�4�HM?hG|���V�=3T1i��U5�,t=I�G��@GE?\�Wq!�K�s�,�Х�.m� ���P9�~��Eޒ�k���	��!�e��݇S��[��Nq�^(?�A�����F�HN ~��U?�$O)W[ޘ�:�/�1�a��,,�p���	Ml�maHL�zq-��+�� �� ������"�M�,wwU�዇�Z Qƽ%N�*������ɂ�L��j-��i*�62�E-�pħ7���49�x��.����I���e��Xu?ݓ���Bc��S=+������c�N*�>�-|����*ɫ\���2��G�����$�v�5o^��F� \΍o"�~hX
�Ze�k����`���ݹ�s9�6�":X,�W{�
� ��*žf��O�')ȒYu�tN�ϴ�3�&2	=�<��	�0���EŚ[Sf�6����s[����gX�.kC����Y=�8�I��K��o�ѓ���W�=�y�d�IyLQ���>�=�B��c�����0'��l��p���T%�w_q���c,+�����E���!fLo����*�K�D�ޢE�f{���-g�/�L�J�U:B��b��D�t�)= �\6�8`ۤHH�/��ڌ2�\�+��g}V�w�=��ݴ�7��mk�VX>�c�R�>�����n\#��`g2���E��s�Y���b��re���#�f�H�GK�l�7C�����@�T{���&���x���XB��SOc![J�a�Y��e�K���\%�3e6YE�&�z��!���?d�HU\�̊�J�`��s��+��"F��Sb~���Z�����������ʟ49�T����Ac��R��攪�5��yFҷ"4������{�@"h3:�c�aD��7EF�_�1����@B���_hZ� �q������*��ǵ"VV'�p���0�Ң�JWi��(��.GR� 9�O��I��!<�����)s_�_��L�2?��5��\�Q�K�,Mc=�۲7Px����t6E>����1�;�OW���#u,�o�	��!�������+�bc5f���k� C����%�_����UU%��@�@�����`�޺C��$�ӊ>Q1Z�O��\�-����ups�2��*o��7Z��* S�Rg���.����d2�2I}5�x��p8^�B�R��Ҥٝ�/l�t^�7�+����%���}� ���mu�ZQ�3��4�ߦ6{��d	J���y5��3�~O�(��A����|%Fޝ��>��YQ.��UF�i�va|WG���8����4��uI�7�0xq�v�
׋/�e�gߥ>e&#�j��J���f��Vr�,l5����	��3�y���������Q*�nwZ��I}
��܋�5��n0���l�ߴ�r���3����Vy(}H�n�rʸ����Ћb&���D@�r�衎&��O��E!I�_LrF��x~ũ��K��[Ⱦ�l4Ra��:���*k(�c�.wj�<q���5�ةv�P�$�l5�(����<�W��
m�z��Da�־���{0�5F�@r]j���6'1ۣ��)��_RIg�j�ݑѭ��[�s�?vh?Q	8ǢI�h>���tup �bwS����L��crw0��q�G�}qpq���_;7��]�&�wO�[m^�V��D�����+Bm|�}�@B���Q"��p��)����֞7�� 3WA���� N��"�QVCfs���`�AN1��8q���ge`��:�2K3f!!�xbr�i�0%��n��p ���j��y|LK<��>(�AoԨ�C�k
�Ybx��C��O�Z�T�Co��؂�Z�B/bbR�I�Np}O���PuG��0�~쿱�W�5��;���5­����WO�jkց��r���tt����c;~�&��X!y���!i�r��P���Nڽ�0с�l�@�1G�u����<��[d��px�x�����s����C��M�(�3������Ԉ4����;�e[*1�����>mƪȍ;Y(��R�":��-m�9���l��󸥂%�Ax�_�u��/܁��J����]rS�漵����ؚG����������=i�=�~1��	RN�\�e�G���	�0ԕ��Nv���*�����f�j.*����ܦ
]��ف?*7�F���Z���{��G�41�+���?�0���,>_�+���-
���r��zj
�BT��蘡T�'MP�^�}w�+�w��!�� Fm��C�ɭf�	��F,ً_�2
5(��3)��(��4�`����Td����h4o�O9fi��"ݘ��2�+l>�����[� �_��������*���3/c�sёEj�#��;���4���!4�Ge��:{��b�ݷ�MHm�U#K����K:����E��:��ƈ� �rL���w�+R�!*{���e���`�eT3���۰>ˆ<~҃�(<Z��J�2G�B��k�U��x�&ܮ�\����ߞ�5Ԁ��~�1�F�~+���}�G��d��X*�]�}i����{TgfC	�i�&�HՄ�V���^l{�xy+y��v���2D�Xe#W���ل�����v��ɸ0۪&���XG3���?�|{��b	��;܊"�y8ow�'�S���/p������-���~)���Ȅ�J�kB�
R�u�ʸfBc��R9BX���{�c}���Ɖ��L��c������P���>� SF���:�%n4�&��9�"D?�+�\+��(�"[]sI0����3���Ic�<x�Xb��K�u��>n��Bhi��]���IP.�e����!����"�c��\	�8�����t�ҷB�,0 ��/���fJ�ì����|���t]����Q�L��ĭ;A.G�~'5�Ǖ5*&����f�+��Q����\L�?��χp��p��Y�n�� �_c<$��:ސ��hM7��Q�!��ۙ�g ����C]6A��#ɫڊ{2h�
��s1ðC���k��A��S{Ԩ;`� �RwyJ�Wv��?�L␛;�N��#�[
�����T����J��[��<�S�̫4�I��;F�JS����g/�?�Q�P��ɍۮn^� �\rڠ����2�v��|�G�*�� ��V#7���TL�A^����H���P����"岅�$t}����p�����B��Ϭ��@���S'����Ө�r��w��(>��@]���hh寶Q.�/� &u��U.k�k��n/�cUX����w��Ȃ�eȪlݮ�x�w��������~�7p�W���P��FS3'����s=R���(\�]�X�K�Sݚ����e����U�-�H2D��d��e�(&&�x��W�}bJ	g�d�G���?��ؠ���8�s��6vJx��+���T��ty� ��y���TF�>�Ǿ�}�X�/���W.z��`����[y����^@x+g��-�<���MD)52���u����UYس�9d��(߆io@������&�I�z>�\f?tX��SI	��%� @�U����0�H��q����|�?T�-� Ԏ���۬{�Qd�a�w��G��C����@^��Z
�&�H�Ye��h����}�:"c�$�,	{##�$j�i��m❼�����u�S�{\`�|���������%�bR��87x'4�}�����U��ZAKU���s���H$�HNЧ�b���@ɢ�� "���<q���X���"-,�#�0��\��)�l ��w�wpf��.W:�_�|�$HYuש�j�<���M�� ��m�ʥ#s���K�V�ӡ�rkJm�+F��+|d�C��@�������@�LAp�T=F�R�B�K@Q[I���\��������!J�|?����5u=K�A��?NhK�K'm������B��v��ݡ(X��si�����Mņȁ4f`�a@ o��w�T�����I|�ka��6�a��_KG�eT�溪�i�9d#I�5R��P�}R�_���BI>d�����a���vT�j������ϋ�|؅��4���T��I;�R�Z4�Z�5���t��sΥ�i��2j� ��FW���$��S�(5�C"�Pbǃ%{4n�'�ޠ����h�}���-R���E�hd3���XjUU��Pq���#'����o���r�$|�Ulƶ9�6i�j]j�M@u��������b;xig�G��=�;��В����]�䏁�[m�u�!�-�z�/���_Ww*)����z^����ӷ���͊f�m��۩��ٵ�	s9���u9Mp���B�����L��sEzSf�m��T�H�d���K�u���4o�<y��j�K�t�4��.y�1�*�xmz'!��H?�eպ~$	i2�����KČTO�q Yq�	<C�`��Z��[�l����~�n��Ǩ�R6v		���agl�^	k0>8��`P�X�?:?�����`����zE�R�@���}����!;4� ��xke�W��'�k�5W>��D��D�;�h�ǃ%G<TUv����C�v���<����q�7�<<b܃����1Y�]F���&����t!VW�
zɇ&�|7@h�*���UG�7�0R�>%����(H�i�e>n�n����г[�P(�=^vP�����o�[LZ3�mA��C=U+�[�vҔ	�N�a7�Lh�o��8�,�4X��`ޅ�����.h8�+�
%}�6
��8�����O�����hAj��(�O_�3$�[�����f���R�A�R�\q�\���YXNW�a%Wu�O��cm{q��+o[�4��dw|f��� ~ ��<w��#_�¤<;�Y��Z�w�?�v:֥�˔sg:�jq=(�Mo�W����@dA�Lq��G)/y�V@�7n���e��4P���TVC[~��{��[L�c�=�@aN҄cnQJN�%��D��,+��!���ƺA}d�z����8E�!�r�<3�����F�E��x���&���u����DWG���mCvV.4�ΰr;p�4�r��IU�kBiiZr�a�%zG����j����t�ǉ0�'C5�z���J��#�	H�x��I���ܟ�
(�9s���>����)h`��X���~!�=Y����p/Q�..kM�*7s�rc�+>���Mu��b��F��D9������>i�������u��l�_5�n��嬿n C瘶ѱ`��(pn���18d������Q!��p��s�d�wN�*`FJ���vDr>�'��)��(y�?���S�÷P"o5� ?�Ż����y��½8��c��(9IR�l��������^x����xé�=r�F��q['���1ݚ� >O>��$�F������jD�X뀒=��R�ߑZ7ء���Xd�J�ެ B�j��3H~ˍy�$��"�zE�g�~�	��[��ڑ�ѝ�F~D�mv��1RlMƁM�Ց��u��]�6a��&���s����Ǥ��v���n�>�נ�}�_���s��uX"?�
���(��=^����N��hse�~�K#G�����z�NQ~��[3������f�_F��6�.��m���d��|1;�����I*��bS��Oz��(P�T���w�˔��u��m�ʡg}�'u�[΃C� zo�<����5c#
�$3)�hQPa���^��ףmm��>��׸�Ci�*\�'C��\�ҏۆc�����"���������%�n��p���7#���M��Z�@��<��3▪0nG����S�j�|�\ ���ϸ��2O�{�������kJ(���BZ�}����~+1�Jo��5G��%�1���i����G���{�5��f�;����\n���z9���4�p�t�k�ƾ�k�8X{�K_;�z*D}����=��~X��(Lqǖ�&q�Mϝ	
�����j���U�����ƌ��,4�'���S��
)�Gιn����qCD�����s��,c�J�ʑ���J�JXK��r5}��s�x�?�\^��t�"���{�K����2�l?���J�H�ӱH6�u-KM��PMfb;��d��\��ng�KDQ��
��c����Fc�{h��p�n��Tz��.4�/���+<r���|x˄ug)l�V#�*�O���f�c�k�^t|�((���Қ��V�[�l^��E������k����D����t�WG��Q�!f�n���C��:Q�$��ךR�~� *���6���96��ba4%v�F�+z�{���0ܼ9I�b��Z𖉉��,�� w��i	C/��?tj���X�h�8v�����8�V4X<[�m�q�+�b^$u����߼����y'y5wf��k}} �Q�������&��Z��rf^�7qMB�i�"ao����<Qk���O�%��;gXU��{��i�)~=�����`�K��S_(I��<����g��Iv�i&���(`�� �s�?�����'hF!L�/���"T��B�N�[�����}�k4_�9/\�b�4��	W3rCP�C��f�SN#�V�%%����Ԑ��k�7�2� �ʧ��5S�H̰\��Õ�9	��<W�7U|�!1P�^ȤO_d�)e��ɜ�-_m�p b@?��^�\�e{�?r�`������V��r9�	$�_R�=�n�A���1" ����yE�����{;ē(��~˰�N����=ZS�T�]-�!��rOA�/��̈́�eC0ב�l1ٌ0Č=6�p۴x!8\�F���v�'�YM^��V��c@����Ѷ��=�Z��v��Lw�EF8��n�j��l��Q)۠�US��8���͵�S��u0�Otj!��!+Y���K��
�dn��{\���:g�]$�n��+%{�u�oH��I7E���=+�Jˊْx��;~�d���u��YA9^�����b��<^���9�z���)`���7NB7����ĈS�}уW�2��� k;����û�c[��c�3*���`4!j�<�-�y��:�=��n��i�F�.����f,-��F	t@f/�yuJ�J�a�)>G��+[LB�TP��֋�n�LӐc�ZK���;�/�6:pz���/b<����g�]���?C����zz�/��������u�5\eYlimQ���R&E��uO�$Dl�h���Hoݸ�<�<Z03٪
z��8Dʊ����j��-���8�H_��jO'%[h�^��X۞Ox�I�N�jA�!{>�ئy�E���]	�eh�Մv��ěw[z��� �Ξl��-�uE�yb;�t}��o��#��U0�v��4�E3B(ո���Vf�5���h�|�I��JD�CA����v*��d���y�L׍t���t��$7��k<R�,ԝ��f�1�,���R<$��pP�I��ܨ�?�ȱ˒����	1y�!<���߰��l��c�@ܟ� �di`�m�u ��a.�0O�-Z��/#���� ��l
��d�����5�$�M��/p�0W"Q��\�$\�w�b�v ��+1��g�����:L���H��DQ->�ָ��ç���֜�@=)�)K�r�8�%tW1������P$M�KR�+�4L��!۵B���״.�i([����s�>-��ls��F������5�5m�;�Q�9�P◘��e���+3�K�)���]<g^�F_MY�{�Ne�� PK�-$�k/�M��+�;��̙4��w�%���N�6�"`lAk�?��D�?bXB��d%���EI����j��qEs|z$��aj8M��%�(�M����%�2p25��S.1&�=���u%����JGߗ�}�c�}�R~�������ɱ����� ���_�,���n�ǲì\�ˆj�������������y���ۍ���D�QoK;�Bd�ك�������I4�P�^�Q�����KK٠qN��#t�Ԫ����8�H�>RA�Wr�h��/���a��=Z�'MG��B�!����r�eA��"'`���~��r�e�b���ᆄdx~��麉.mG�[�	���-r��<�ӟ��Nr׸:�������<XO���[}C
C1�kI7FXV�����d�+'С(h�hA$����k����>S���J���ԁ�؄�|���\ǣ����Ɋ��HO`��k�a�u�0�S���N�#?�+-c�F����� ��%F��<G�AL�/�$hnR��a��z�豅��gORQ��v�O������֭���"�|j>��͐������4Pƀ	_��,ߠ�Ȇ��v"a�D<1�^&��?��L�G N�\JNj$�����j��i��}�%�	3[[��z�&%_�5��.���h��l}ɇ�v�]���Hbh�,�A�.�m����ђ���}��t!��P4ǅo%�X�s�+���7���^�bWBe�3��|��QT��.W����3�a���ft�$��y��*Yz�c��c5hW|p�ғ�0���u	}@,��/�$������.?���2���~���:��yY�
���
�2�ejކ�օc"�9�e����!�6<�<o�AU%�/�ic_OM����Uv�LR	&��w3�#�����أ�,^�?�B0�b���� �t?�ʟ��E�5`*�S��B;+�M����4s���`�LA�����{#����j�=1q�5P��5X�kY��o��^U��1i{�.���zh������E}n��|\�&%1w��65ew���������d\�8�ߜn��e�z���vLv�&�����'�r�� =	�O|��{Z!]����2��q��L@����Oi�zv�@�%ص~,�C��ўY�J��`;��d9�}�KWk������`R�gl���zn��P�/���ax@Ȋ���
��h���Ʌ0 _/r9����T�q�ZC���YyN�,? ��S\�L�XR{N�j�8�W��� gh�()��,Z��Z��p2�R��������hv����EWa3J5��"�^ߚm�}=x[3�t��'�#�5���m�����O��Jِ�>�#�&��뙘�/��4��W��bٟxq�ԣ���J)���LeS�Rs��F���a�����������j��XA�Q�)T�Z��c�<�XHܙ͕������ �_se�a�
����X��m���kѐ)� Q��5k��$��禒�yo!g��ŭ�w�H��X�A��iڜ�R�X'��ʌԋ|T���-��`���s��AґN]��S[�PU�+�!Z�#����<Ʌ�k�a�_U��FL�t��j��� ��f_	if��Q�
< �U*ؿM�u���;�V�����#�3Tr��WV�7x�}����Y���.���P>n1H��6eek#��Ԝe�^/{6�6����~^M������j�Ы�
���BǕ&�,����zi��c�����u�Q헒�<��'��L���R����M;��Zd`<��Y��X�	�N۴����j���vڥ�a;~-���f�U�,�?�8{ ���V¯���U5o]C��X /�qA[2R^�����8���j!~&�����w|H����<Tx�aL����0Fwc9�wmP)���&�6�\(����[�l���+Zuv�	g�ۤ��U�Q
d�^�.BR���I6�QK�׎F�^�ˊq���-���B�~n�v����"���Y_ׯ�Od� ��w%2t��{g�*ua�P�=i{�������CƯ�ݜ4�7ҊX#F�t���[��M@�hxU��@���]RH���3	&Ѧ��5�+�0��-�U�
~f)�`_�6h�1�?kB����
���X��{_;f���e��w�Ï�\�������s�\����,��%y���n�b�҄���&��)F�/�DРC��V]DC��y�c�Z���>g����W),6����U<FF��2�#��p��CwF���P��k�U��{�o����y��:�� �,�����HBxLϽ�L9(��,��Q�i���+�{ņe �ԳdMB$ւ%n7�D�r
�{���"c�b��{�Uվp�����Ớ~��8�W(a~�Ƃ�"�G@v��dj�>I�l�n{l�ߏq���T0iP��$�%-��A��/��37=^���(�ì�#l��mY������P5���-����rȅ��/�m�]]�A��������:0㲺��^6(�A����B��LRc�e��0d�j��nq�6��p���f��ggQtY��DJ�kKj�\���l�����M3��$,Z��A�_Rd��@�������,/$%,���Du@�ȱ�|�,z�-x����v�HlW����as�J����ݮl��<��x�L��,&�e���8L_T#S����c�h��������(�=���R���JB��)�	+_�$�W2��9y��Ws�O�e�(^��a��?��bK�1v��K$�n�(p#�POF��Q)I-�Q<g�u�-���6�,eQ=��K/�����}��"�.�ә��n�MR��%N���%	m�L��[�������bg�e���6|`�Q
��5�Y�2,M�	�� ם��@L�Q0�Uk�O���cw@Bz$���7�l!��r4o�Et��M�"�����FK��7T���٠�>.��b[��M�YO�rQ��&4����lN�Ů��҂#;���u���֯37���f��鮦Mǯ���v�g��̿��V�@TM�7���.���)3T�1Y�ƣ�f�0�:ʯ<�`���OLF����Ε��g�#�����o*�4z�q2ފuKn����c�[�,���xC�T1���"}��B4���s��f5�Q��� �-�N��;�F��5nWN��g��+m�M�:�_���/�@�����!~�&*ѩ���<o�x����|��6�<b��:�j%*"����Bz��ӂ ���a��-U�`�G��T�K���ou�,h�g�q�۱�ٍYV�2-%nwWěܭ{$z�.i�(�<�8�ܤ�ް��n��+���	�
�j(p�_�)k[��3�c�֚+	����~���䘢��kc�l_�P=*�	_�o��w���P�Ю>g'�5;P�F܎�Ʌ3�|�&�L���uW*H���ٍ����j����R3�md�r}h��Q\rh{�z-��M�б�A.���n�2`�7��&�,C�׺�W"�

�\8J�%}`rtu���� �գ�����(���0n���ŏ�J� �#���/U�+���O����殨�b$���	�Zq;]�������� ���_�k!S͍TQ��BN����޵�xNQ�<�yoA)�����[��H�Dڦz�cFH 
I����*��w���P�Sm+/�]���1�W�5;覆����P�=r��#����7�M>�b+��T�#�ո��΍l�%B���pz��\)H��gŁG��V�fu��8��2� ]��w�&���h���4�~�?�h�n՗5�ŐC���fڱj Nd�I�.!k�X��]Jcsh}�7�\@٬q������Ť�I4T���X�uXƣI!>N%��#��w��������p�������{HQ�p���I�y������-qa�/�oUo�{�HMS�g�x>�H���c�3�bv,sM�����nb�EX�uP}�e��m0��%S?}a���6�ε[̫l,����?�v��$#�68�`,8gY�:���+�����]�_7�2��T��%��<Ʉ��U.��4t�4��e�#!�����q���˖?��i �(ı�m�"�D���u��>O�܊�a�[�h�na���PW�i
�w{����H�ģ~��^Ou�Ц8���~s���5����0w1�H�
� ⃧�i�!�|��'vXq�����q�m��˧�W���3|�r�9v�1�I�����yN,_v��a�vÉ�PtD{��:�Y����R-�؄���E'�=.�p��qRm)�[�e2'��+v%h�[}���6������`�*��
`�S	�ZyH
�۵%��0���jZR��r�qX���R�5&����F�`h!#'�s�����n.��ׅlb��O�͝�V4�S���t����V�	x�Ysx��hIjWʻLA_̸z���\�� T#�eY�J��n��Jmo�Es��κ���CE��}	0�c�^����Uk���������[m+���o�zF�?4�w�;��n�`�>2J���M���Tv�nM�5r2�8�<&��`>p��������xF%#a��B需 ���jKWa]�{���ي�?�Ds������ib4ȢA�����]?m��L+@� ��f�(���å�$E�5�UQIrO�eq"OY���g��(��>ci24����������)�m�<�]�tr:*[z�Ax~ ����*f_!ǁH�]�7�w����8$a�+�f�^q{��Z�q/{��j\bq�.�Y��?��1yB�`�AjF����I��hv�k����"�df�jJ�_������ݘq_���)�"a�:�&�ˀ���P	�GO"��^)��&���b�V���hPQ:x�����r�5�Ur0Ȭa��r#�r/�&�ì����wi�g�b�X]{G7���0:��Y7��_�Q
��TL~,�OH�xH�$�e�;��S,�|��M��E)LWB_#��.B>���4?a�L��S�X�:9L@���ܿ��ʤ}K���[���/���뷓֥SG�c	Y���7`��㾿O��<�Ы)�p�˴�˞U�Dy'm+f�k�9󳝣䪣�j�m��eE�xJ�W����@&F� n�!��o���$|r�4�2���Ei䏑_��G�[�!�6C�(a��
��ZoX�٢(A��T�B��QN��Dr1"����*��׎^t�c����Y������7���T�?�I7�Ո~����.�����F�b�����QWd��ł��U4t �`�~����P� ��@�eX
�
й�&ҡ>�T`F7em2��&j\�����Um����Ͷ_.xv|n�7-���w�p��9$� �?�2{�,�Ѭ�����MV M����-�J��MB$q�]�Q���:ˠڄ��?Q������5���#�	l��%[�Ǎ\�� �%7��-��ن�0}������(c�����
8C�	ή�aR�?�N��M�I=3���Y��,~�Y���ʓXF�Q�+6����V7L�����wiEh3
�r�S_���ˊ
Z��E�Kz�C"���xK̰�5��~
Nl]�����Z���zC�?�%1�Վ��c�4}���6wUA���H!?�^�$ ��G��s�R{N.���Tڵ�u��!�b|�1��T)�v�5�P�o[s����7�^��H��>+u��c����]y�
��6��o�zST�ZK�CiCqm#�U��Uȗ��D�Rw�"����B\����W�e��|��ͥ�֭���/����<�i�W��
�S��!m�d,@��SJF�6�8c�%*�yU}�?�IR�E�/�9�j��S����O�7�`E~삑x;�D���n����bL�R���'`�ֹ����E4���"�z��4}~܀i��?�C��5y쾦9�T���iH����������r����)����{�7��v��9����������	�	�;�/����/��v?"Cu���fw�lu}I !@#t�A�팴�FO{�1�&�M��T� ɸ-������H��1�`���H����v��v�Z;m����Uy���+>�Kk0��5���ū2�[���/�D_}!V��{v�� �B�E�rNo��Cc'y�G ���?��^2�=�m3s	2%R+����AB�!�6sO�0Gh�+���E��#�^�4��|�Z��!�P��.<?z	��6JNtBn��N�|ݽOo{�1\.,� ��	�(a5էIX���5�^ȭ���`��L���4lBL"^W�f���������.SR�nI媚��Os���,g��л��Η��Uz�J�H�ae~9�؂�-��i��&|�^��0�e:��#C�E��Rl�Y�Խ� ��c�Hiך\F+
�q�X�],�/!��,�A�A���_?�g�C�ut6bu�-Z|f�ɓ��̊E�_q��\����I��^�H1�ψ�J�V�����<jh�A�L���;�����;}�L�
�Ih��]]m�Ԩ-8�VQf�}���4��5�9B=s7�n��0O�صB7#�7jm�%���&�<݇Ȏ�}����8V..%�� d�"�ԏ �"�L�r���R��(�*��T!B� "!T3����8O&^m�Nʤƴ'&���z
{���V(�D�H-������C:ag����ۓ������S��YV��+D���<�s�g���p�BI�;�E�g2گBӃ-γ�.S}H��㩾4��ף���� ��ɯ�)j*�f�s��Z'i�T$6±�+3��7\�Vt�O�8;jq�]�Z�p��u��k�9�XX��P��&�l�g;�_+\�.�sŢU�p�2Rhu\� �i�71K�.c�w��
�6q,��A��F��+�:�'��/��b�	�K��Mj�*= *df:��L�C��Iݓ�@���_�Kp�{|vѭ�*����S�>��#;u�e�D���Yi�dd܁�M��L�*{1X��/+�$8��3idm$���%:���B�c�*Y7B��~��d�͓'�1�\HM�q�{.��t�|����8��o�dd��r��4�4Ʀ�Mg�Wo!�O��S�E  #�Ӡ��v�l�o���|k����:ة<�҈C70���J<�I��љ/�7�x6�C��A֟�ϡm`�]��j z�qDŲ�u�L������52RƁ��bHs���\�J����@!*0��D��;B���ơ��S�+�8*9���hAO$��u�����j�|'0�=�=w+������j+u���D��\���������5׃����^
we���p���:�H :�is����o'm��~o]�����q���p@g|JvpE�R���� '�|k7k�W���60�?u�w��e��%����
�����<6aSU���5��+=���V�r�̃�|S��(}*���]�xˑyX�Z����O�"a��-�BN;��{�m�f05Hk���h�i�x��a�?��{�e��8����i񀎵���!�|s~	�]s���Pf���2lٚPIA��7�C���ްˡM�
���6��q�*�/����������'��0>���B	�����q�5��6{Ѹ�Bᕋɮ 4�j��=d�
��;ϳ����x�z� �pK�!�'�Oj��6����-/�$�+�	3x��I��6"'7�IX �f� LQZ�E�|�_�/���D墍c>!�#���1�s1}[!Y�%�\�\F��:cp�Uvĉ?����]S�Xt��e1���j�l�0l�({\k�"�!aW�0Q~o&К��~i���	xH�j9mjd�n���h�^���2�˚�o��0�Y�A+��5>u�K���F������Gy�(H�q���E�ʬ�2����.t���nI�6����4�t�[`Z�*zj�����p@,�)t|�m
��dGW�t3�k2�(o�}@b�E��6��]�_ѯ�9�,w4�V����K��u�/q�'��[�ek'G�YR	����љ�>x�� 0��<����V��T���&���n��%���0M���QZ��BH1��PEo��v��snt�r�쿨��lJ�����9�D&S$�n���)J�-ݛ>|�h�\�#aRt��Φ�)K3�OR居i(�c�R ߤ�=��4۵,����Oy]��~	�.����jƋ�FF,��i�ܮ��u�)��J�᧘^�r���/��}��%O����t5(�
�� !jhE!���W��$�.ݑ04Bg��p8z��I���23bA���`:�O�Ӱ�*!b�t�|D��ע�>���]�\�!�+��}6�'�����J�9n�b��a�����m�Š/m[Bd$w�6,�-Y����Vf5�|��M1��}g�Dy;�n�����T��;y8��e��=F���IB�;T��u���R��HF݄%�m�G��!���iV�=ˀ<�U�)U�K6����[v =�OF?�N�����?*8��P	(�η%d75Wx�N��mI%[��5��C
�Ƣ�/h|�q�e�
�T	� �]�*�"t��;=�F�)p��u�/6=��D}j�V�ZN�}S��O���i�ˑ s�������6X�����_o�9Z���V1n;�[�MrS���?�_m}�	�<��e���=I�i��F��?�;|�Hp�Sj������C�M��9�R�*ė	��q��.�8�Q�S9�k�=�+6]y�Y��Bﺱ�Z�c��Ǿx
�d�IM�:����Xoޟ�v����ʿ�8;���gN
��!���#�X[Y���u]��,�����`���U�5�7s3i9��Ǒ V�������|�����۽=��sF�e��zO���4&.?��9ͼ�G�ƀ�L�\rWh��~��Ă�/� �>���C�S����]�4j��K#�o�u~/�$�|��0px���0��i�Q#�.1yM�\Z�q��yݡ��$''���܁�wm��|e]�y,���l����e9$Q^"	{qМ[�GOW��-W3��hG�sZ�*��Z�so&PV�A�-��+��B�}��Fm��'��M!u�_��UST`��hxlG��"y_�מ�?�>�+���S�d��'N{S
�ľ�u��;d$F}a�F؉��=����A2�3�����D�ql�M��B87������]A��9S�aQ� ����]v��<D����cY篪��mG��2��X=ڰ(䈱ܖX��D��tEL?�e��������	4r��|8d���y�0&��Qz�� ^����Y��Q�~f�X��%�Ԏ�5%>|7�O�ݮ�Â���;az����7�b������3�j-c�\��G�H:�i����<0�x��b�Jz0�K���j;���K%������pI<P\����>6���lc?�G΁t�����+4���r�@[�./�=0���}#�"�^Y�ީA�C��|���L���I���)������H�v�-4�y�z�y"���CnW|�eQ��-�r}v���Z��:pc����b��cB�Z����}7TfU?t�Ș���Q��ݲ*��q_O>gh]���y�����׳�3Y"s;yM���jrӁH�9?����0���_g�&�9n�aaX�Vw(��J,r2��_��I���Ԓ����UC��+N��ΰZ%��S_ߢ�OmTW���Y"d��q�جD|���f�:w��[��ޝ��OJ^0�ʄ�^�4QF����o�d�m8��V��2��c06� ��&o(��X5`��P��X8u�F�Z�<!���%�YSh��Rg�a_g��jj)��1~����H���w�^@OP,�GBc��f�
:���Zq�b@hI*��Q�aR�<@�L���a�zko�� ?/�}�F7Z�*IߒzoЎ�
�ӪvJ��L�;�.	8%6.Șo�;�Ɋx[�����&��O�I�A���)Z�� ��_f��,���`lb�L7o�c�Ѯ�Q��c��,n�`M��$����XOc�J
���i�I�o�QC�$����o.�9�G�NW� `�c���y�N��pD�m@U� ����q��?\����C%?5$�>�7�z�ʝf>��8���bc>��
Z�l2q&v�":e��e�6f�����zv�}�h�|�����d��y�8�q�A'&y|��:5Ȅ�[�K���t�9y�@s&����J�w�o�k��A]`�]�3�!����淭tx�0��6°�˳�eh}�vh�X���g42��LT�(�nV�j?�f��#~�c0@��.�J�$�ָt}��j,>��A��Y_�N��D��־N�M��r�1S7��2�n�S�,aw��Bvk@u	��¤�.�2�q�oN���x��U�X�,a�&sGI���%�C� ��w�u�@W	�(9e�!�=�`�~��p��r�c_��>�k���{:M��Ƥ`W*r�d+�2����}����7����Z%��XT�H���x�3�B��{�~hB��j��/2�y��'~��*Kua|��ށ��2����fto�DxF�U��%��Vƣ��k�sc�ط���Dq�ڸ`���H�"�*ݨ3mPO5?�V����3���I*7%^�Kۈ��r�b������(:���#��@1���$�3՛�x��zO��� ��s9�=��=�>)�_@א����+��3�q�:�{|��(��[y����K�z��Z�}&���$wcO�s�>5n����|7d�T�s�`�R��7�h�ԅ�0cND�!���d�IY��$*<�u�f�㠬���W;�+�.$���m��p�h�MS� �f�dj�C�մ���mi`K��[�j|D[������8@(T��'���6���;�p��S��x�(Zhk<����z�.�'�=TQ�,{��"��_�AMWG�a?�z M��������R_h���껈6{Ҁ���'0_��Uw�VW��ض���(C����G����6���)��od�����
n���{5���|�{��
��r�2��7����������/����
S�R��P���f`�$�HW���`���=3Mo�?�5=q���a��ϵ/O�F�4�6"F̝"�����e]6�9�$IV���DG����*c��}K`�jG�J{�E�[��EN�a�H5)����/����L�zUz0�������(�YК�~��D崱6�`�����p*Tڵn �(��7�1˼mF�M�����������9�ɡ[~���@�y��3�&�Ј��[���ß٥�<&��<A����WmMf-��;�toy� ����oZt�.��5
xL�'�{Ҥ�X�gZ�)�dA�lC��l�)�N�,�e{&W?���#7��V���>��Ю�9�,ci�騠A����"��z\��Xf6"����BJ<��/��uwY�H���M��iq�=�[3p�+ ��� R2M}Z��/� �w`�Y�M6IOr��Q���A�{C3���(��b5Ҷݕ�UO�-�B,VDc�R�T���K�<q�(�E0{-�����2tu���8��c�ߣ"<�P���r�P��-.Cl���-x4�U�,ƍ��s�����`ռ7I.%"���/�Ee��,��,���v�0��k�RF�&��w,������D��A��� o��R=:����0�H�!?�S�v6�y��fE'�BMF�=i(TH,�(���/X����0^�������9>;���
U-KT��t�)��K������s�ʈ EǇf��ԙP[���Puu,W�W0KN ���G���_�VT1f���d�k_�v�I��6�M�����eRN�C�+$B�p��&-Z��k#�$�^�if��i��~.�53����ɎA�@�ēS�m���/�:�}O����\�4�&�b�`�bɗ��+��	���é�Jʁ��AC��x��B�3�Ӏ����\��<�*xO37^w(��0o�B:��0�#��_��q���ª� k$�^+�H}�������n��wحi1=�@3���mz<�^	Ej��]EÃD��v>C�bi�
mnD�F�fܲ��^IM3n�w'��|dr��l7������c�\)������ܧ<����׿���#2�J�{g�;[��@�@��Lţ?{H���~����[50@q�(�	*#4 ���-ų��o��VS���^^K�I��y�B֘�Ի�Ek�z�A{��GK�k�K`(�F�)�~�h�q`���
#EP����O1o'���_! 6#a��{����
����$@ܸ?�S �ih�U�"Nw�+6ϵ1g���k����Yz�M�������5*c^�bw����	��-F4s�:M��c��a�&�Hc�F����6F ��e��
��]��E����%�#���g���J:@*�.����0��%�X��d)�̜�tM+:l]00 :�)%����S���,)�Œ��ov��)rM�Q���(����%Z-l�b�i�E�p.��5��8q�!�q��2@�K,��26G���U���*6�MQG�i>�6-]3M��	�p�Up	-P8��gsƢѰ�.�?�[E�cJ���[�Vn��xA4|��iz�V%L!{�����
���G�w�ٹ W@��n$�'����e݈y��mF�		R0f�(�n������f������GY�C�8����m#k�fL�wfЊ9�!Y��!Y�/3���l��n�Ǆ�$�,I�%4�$�Dp[�/[yI��{��^�j��kV���j��d�#�BQ��m���� ��|���ŐB\8�3$�3'0�')4��}�Ku����OT=P��l��kW�ϫ���ǔ�����E��Ъ7*����2�ou}�JO.��kɴ����|����X���F��ϰջ��4�LY����19���@=�zG9 n��x�9\��݃���ö?�)�)t�;���A��C>�,�"�(��*Ut��A������gy3��ի�����B�e6'2��9�|����,?��u�s1�K�k�w�\�cɾ9pm��-��C����#_K��K��9����]?�J���ͫ���	�U�̆���b�xƌd��0Y��'� r�,��� ���Xi����O�!�bY�Jї��	�y?�X%7�9��UƌCEv&��w+Cz#��_O�0�բ(�p<ewHR�]�)�6vt5���_{��G��5�M3�%�+Tٛ�7���y��_�����G��蠳�/sٰWS��C��k�xZ�ቄ=�pY�u��
�b�`�@���
�^� rq#��'؟G\��90��j�s�)��I�Ĭ�����ܒ*B�d�i4P�І��$�[ٛ���O����P��(�&;�Awv��i:9�ǋ�Y�1��=!�2Jw��[�>�1��G��s����K��T����jۖ�aj����?�Y0��p�{���f�j��[�`E!5;[}��(;/+�d��Ao�b���148�>j��lsb�^��I�qa��U֩�i�)~bc�j����Ki�o�U�7ʮ��
��R�d�9�H4X�<����쿅��F�������Ė}�@v!D����%�Fs��;6����x��4��oW۝`PJ|� �uU�n�),}����J� ��=/��G|Ѱ�?^%��b����m mYՈ	��u�Fk� ��t��[j����F��IP����I�r<�7!~u����i|����L���h��XnA�G��\�)Ί:�r3n@l�&��ڴ��D��j~�t<N�f�#���(����r������ ��=E�����"ml�?rt�����5�_��!Xa����xϤ�/f��]�M��r��"EySf�����ʃ�ƍƳ>��A��F*�s�{�H�57�D�C{�W��9���zi�~  �N4A���;�f�N���-�dFq�o��C;ޜ��u�������m-2K���$��1�~awө������b�t�]73Q��IaN��$�u�M�DUDK����G�o�Pz��Ћ������,��N��6���Jm@;���+X��P٫�X&������7 �Iؒ�o�Q7�1~���T��>��[��A�s�b"�5�W�R�T�t�nC_���D���oζ�O!VM|���H���./�6D�Tv�B�}ӣ)�"�%L-E-IZ0�;̙�dl����%	��ɱH���6�
0���#�H��ݨ�.���h�nopFj�nF�E�Pp���>���e7w����1G�����3�&-���̳߰F�����QtM/��
|�c*���C�m�@x�Z�;P� $�=���sq+��M��z}���1s�(����%آ�~�{�G���ݖ��PnU���z#��1S��;/��Yι4h�8����� >wI9�W}.̾4���0��^�8�ZRH��ٰ�V�|Ǵ��Ƕ�-R��Em-���L�E�.	��&R(Mx�8��)Ua2�P��Q�V��u���h��؝RT��TN㢝�0�Q<e���d8q1�Xn����D��q�����3�E�X��V�M˴2FU�/OF �Xd��$��[Pl���LS�	S�����G��uAx䥠UM<�vk��9Y��6�$���o�:���$��8$�;B�@�V���Z�����:��C��TL'ti�J��(��Ex+�L�d�M�bFU���LFߓGQ��$hl���#V�츚�/����i��Z�����Ћ������e�9h>���?��9k˵#-����q@W��Ց���/�	A;/����h##n��`ߖ�F�L�?��Fì$��\G/Ҥ�;;2���!L}Q'&��'����ٮ�N5�\��re�:���e-�,�q��-�φ*LH��jke�=ª�_R}~��E� [��C�#(#�ve!꩕�疒�6@�MM�Q"!�w���Y2�V� ��.p��,�w�����d"�򘡋$I~�T,��V�9���x�*Q��"�4tG-�f,���`Ę�of�k�cO�.��L��m���l^��M�z�<��\�;-FJ����#a��V��2 ��AB�C�C��JI%`/���r��i��n���kD0�Z�"Z��c�@��,����Q�lq���w���ˇ�=���E�����/<�	|Z �l�&����{[�^%v��]����J��Q�k�5�d��i��/�Ϯg�������px�*UB'�̚6�*�Wm����8�5��c�?S;k���[�����z�fָE1�ʭ���:�.gr}d�S�)(i?��
o�K_�#1�k�x��h-1/�.�� ��*)MJo����[�.��:F.��m�o�r'��n�-%I�u
���5�"�`���	X�F�JG�#�a�n�L۰��0�I�W�~/%x�2c��΃�6���\.}���'�K���9��hm{����D~�'��.B����駢���&�Q���K�d2q����Ә�����苖���c��9��&`�Ǌ�l����ryE���*�~ȕB�"�w�@�0���`����X��4	���i޸yf�%Y�d5&�����������U$�PK����b��ɞ���ʹ��)2g�;dR���\1s̱TP�����x��p�4D������-��o8=�4?l�^`]����F:8�H49[�Q�+��!��i]ާ�

O�MT�|t6�sqc���Ό�U��V>���WY��S|��͓ް ��=�;и��|*?9��
>�Q>� 8��`z_S�����N<�d����mG�7ϳ1����w*�*�V`v3t�!Z�Q�^!3�@�;��*�堁hWb�Bx�e�4�"�t6e������&JxGꨌ������Ra?�^'���.���G��~)���#K��wwF�����uy)8sk&+$�uJ��ò��'��U��
�b&W'�}�:5w���!��k}�O�y3��k�-�ݭ`ӧ����u��F����x��L���I��] ��B**��`� �oIXD�Lvc�Y��S��-�@�vI�O\�|� -!N1����4�&l�L=>��kn�$G*Ğ�un�w��`����݉���3�����=Iǖ�������	�aU�Ɖ�RC�]���g/�΃��K\�ͺBa�Y����bA� +�R��CCm�^ɧSKR;I"9?��F����6Ɍ�t<F���u����ZMA��maY$��HmO!Sz����ӑ��j�$���1pɂ��]t�粐�W�.Z�W�0��uq��9{���9�����|"q�ǉ韵�:��:vb�/*��K���mr�銋�0�Vʗ(p�o)=�g��\�g��\�	YQ�(��q�"3��U��i�O޿}*���,rޏ��B|H��*�R{2hmm� �YF�~?�ѵ�(=P�f_�W(��cg
P��aQ�3XΝ 9TjD-�1��-؁��ըkj�]�Z�� U�5s��2\6�}��W(:M�""��%�-�w�������"3�\e��m)v5�5g�y����4�)L�P����w#�pN���:�])��8����/��{�[jg��z�� �@�BÈ���`VP����8�_ì�ϡ$=K�T�`� u �k#��L�q��소u���J���{����.��Plc�ڧ8lW鬤��x'�'��\{5��qJeNkR������7Z�x�t��Ķ42��3��5��G��u'I�,�Vbr3K��˞b׿�b���{���6zNMsr�!�B �V�V���~7�[�r����zm�	&���q��D�����H����Q��}����#芋���*T�����T�H-����J�O��1��Z��9�۵��t.S����ɨi�
���OVh���XA���S���kW
���ψ�����.�N˩��
�7�iP���I�7����
��FL�_$�g5ə�����&�%R��B	�M}�`�\ǐ�bVN�q�<��LJ��Y��o�q^U�i���/!t����&H}`^o�`�q��}Q^I>6������rj�*��{��k|m��B�.h�����������ؼW�z(_y��lRTn8D3uU��F�OMRn���J�?�%ӥ�*L�H���a��MK��G�w�
�e���+�����q[��2�l�7û�����Ҭ�!��Q/͉������{��X1�Јg20]6��m�t�z�ڛ��h�b�䓜�����R��J�DE� �����tMQ�!!ԅ�JkKpvLpk=�Ԋ��?�	T���0h���;���p�'p`:)��~���w�����O{�:��ln5I��N��4[�>O���r'*;�{r�_?m��մ��Y�q@���?��fP���E�E?>&7R��oO�Դ�;��!�š���br˃��	�i��D����@<q�������rs��v��4W:mo��Uk%K<��\���p{�*}�z]�M��]P��ua��D#����Cǀ�5:��.o���_��,u�]K�{�;�c��=2��ᛦ2�ELQYxB���}Q�N�3_�� �-`�M�����tদÅ��`�f��P��'�3�!�������<����F���	�g���g����W��k����d4����b=�CS.
~i���xe-�܋��NMÍ��K�ߣ��,�C�f1����U�|�s$���3�u�[-�w�(���̱���g�QaM��6$�\��7 �D ���>�)Zmܯ�#��"�<<�Z�R���� 	g�b:l���	6�|XM���m4Gz�������
.�/^hVA��e�O�2�'d�+��lW)ûu��ى���[$]��� p�K_�Ac*�f���?%< � U��t�5��!�E�?I���s�^\�l��L�1�=��񤢖��� ����T!n�e��]Y�^D}Zv�b���?r��e�@i�Nȅ������2|�9�x�g�.� ����/Pp`ġ�6�t!�S�\�drX_��Tn���T]�rv����vH$�!�.���OI#>[�8LH��A��{~i��b��
�4>)o���!͑�핦�ߦ;�UG�VJ�1(S�7zH*
|7Z� �(����ٰ��Z�v2d��#��Æ�U}��l�c��_�h�����D���*R�C[���Լ��'�=���[��fu\6���l��2���h�G���E�#
6ٷ,�6Qkw�Ίˍ�%�"	5�o8�ҏ0����ۏQ��+W���@�ΐ~�����lI1	{+u��YP|,D�wC��"[" ����C/�9�UQ.V���}�׊"�{��/��|*v�T�WP��,��������tl�W,��~g��O6:EPɡ���-�6�WS��Q.u���*ܞ���<yp_:jc��hs[�����a48�k`F�������G�cYd� /z�
��D��.,�W� 
�� W-l� Uϱw�^�)�jBC�<'r8`"B��ƞ��Qy=>c�}Y/��S*�Q�!�ŌE{����|��"#!����[�q�ig��$�� ݇p7`%P]���
�!@�2���>O��v�����i]�1�O��64=����(ڄ_Y���u�I��M_��"V�=9k�9��e3_�(a>7g���0SW�w�t����0������$��9{�Sy
p���||����7���OY\��J��q�Yڋ�̤�������q��h_h�S��J�Ǎ��q# HRk�Z� F_�I���#�U��w���!�DQL���K"�ϒh�f���,G�C�h/�x�Hq��y�w����}Sm�h�-�j�h���Dm��FJj?i4�y�Гo"�)H.P߹����Q����HO�c>���#�k9O�~�sӋj�M&�_p>@ �)T1b#� :�^=C�/r�/��@�&]|����j\՟m�B7���=���h]�ܖS�mߝ)z��ۧ�T��e45� ɍ
 ��@��T��W��)�X9��lP�|��XeX��x��_&�㌳�q�]�Li;o�㞱�(2B�ԫ��-�m��G�0���>�����@�Ѕ)1��;k��!�Y�"%�iTJ��Έjm����M�+e6�8.��B�ӳl)g����y����J�S�%m��K�IMu։��#������*���:� �rs�%���46�.)�xKrl �lH�p���h�����@�Z���	��o�Vt|4�U�(U
�N/%�;��MVc�gd82��-5��䙛��]��A��Y��刈�`���c�t9��"�J�����'������k�+�֯��[y< ��߂�����o����9����5>Pc�q�51��ŧ��YwUj�L`l��B��Ղ�;�;���i�32+5����e`�#j���'�b�ȷ=���Y>e����q`a�It#�vrj�2�7sm���+����j��[BBFu`�Yn��-Q�5�O��JN����2��w�Z�o-o �r���*+W��]�ϑ5��z �W�ܽ}F#�5�m�� ���\lG�Z�'���:����D4�v�8����p�bmv�:9�`�~P�}��5MR~���ÛBi�pՋ:���˦�9��͙��=@�D�`��tM4��j�م
`�Ҽ��}�}��[��}��~����	�ǑH;+1� ��`n����v6���o��?����N�wP.��\5-�ܸ����U0�$��m�{����R�n�_l9ZҴV�u��O�N�ߵ>���#n����rkV{�Z�I���_�^�P��Y$�D�F��hg0�3j�n��>^A@�߈�*�}L?f.���Z��|8��9�	V��`i3�nӸ���Q�X�w5A T��1�b�®�.��i���O^$
����G"��Pj%�?ƌ])Z�YO٘�Ø��ʳk_\	�Et�s������>-�X�����(�=l��	��s�����\Æ�Q}�8��Q@b�G�y�0�^,3�unԕ�ѽ�,�F+t�+I2�!���;N���s����7�V�Dsw��Y�s����S�}��S
�m�0�XkK�:N�b��%.;@���M����x��UԔh�FKۂ����ۖ����>����ߴg�>j*7�t�l��������r��W��f핒Ň��i�U?��r�d~�V�&Rm��~���c^"Q�k'��G�0�� b?����,�ViVHdI�	=�Zt���Y�D���q
�Y�[_��XeG�<Jy?D�3�z�b,U w��,kF��m����
<Ը��j���J�ӰM���7�f��8��E���QB_oW#+R�\��|=�C���<���0�����}��b�c��9�ȻJGN��#��Ҙ`�`����C<���&.�,�dڶ�?����rG^�vAGIqi+CK�H�俽}hd����x�{Է;��T�ݏ62�,���}gm���(�ַF�6sp���"�=�<�M��(䧎HK٭p֌x���<8��u�4׆�I���l�ُ$$�#j{��P9GOHMk��	e��$� nX�e����F7h�����*��m:-��&�[oV�2ҟ��>�՚��T1A/����ܽ^�zXJ6�A�����<�Y*?�K�VU��p��mQ��	`(cZo�f���s|��䶦\�Q�j�y�jaܥ��c����Һ3��*G�<����Cӯ*�7�iB�/F8A'�^�! /2�;�^¿B���:���;�*�	l5��iu�5q ���������1�4��|�J��� ���y�	����=��/;� �J�?�U��?���M��}T=T�u����gI�Pl�[=��;��&�M���jG�׎^��4���8v�(�D����+����/S?x��Y^6t��~$nXoѩ�|��L�sdz�O�������y��$>=U��O؏i���{���فe ���M��l��`p����~��5
��븁��D#��2�Pz���P��;G:C��fم/r���Z�2 ���(-�ư/�X87'*`���⃰?�D�,x��*K�S=�&h�J����*xN�Ss�B����EAb�eqP�1CϿ1�w {o��Rf��8}#zV���k�*���\��o��l|��$��4+t�~�D�����GӪ&���X�%�JL4h���8
��N�d�g����V��;Fi;���S�^zJ(���e�95.�v �
5�<�y��`G�nd���SK�a>����
�����Z��W:�?�\&<խJ���r�����B借�~[u�mW���&8�Y�S*�j��pVv��P�t��oB<�%M���R���%��#xT���j�K�u'TJ+8f1/$����=��IS@pg�/Ձ\��o�kW�R���Bٟ s��ẀM��|O�%���k�6�f���ite��e��VH��ӃI�)�<���k8?,@�&�T�4q�Z�\]�@�&�n<8Fz%�����;���m�o;���"�g���d�,E2ր�=�0�CeUZz�!v�����A�fA�x��Z��}=B�E X~ �Y�t]	8`�Z��%Љy�&3����I�Mb,��p�ӆ�;J6y� ���.2�ڷ��s���9D�`�bW2����%��}�ݎ���a[@���,8_^[��M<��s;��#�2$6��[�Mav�8=��ޞ!� �axԇ��Jg�&�3�a�m(+��� \�������P�-�?pI�ٵ����M�'�*c�v�?�I���Yk)�?R�R���Ox��DF�����4:i+{ʕx�Q����ԒQM?�F�)m�۪�@,����D�&p�<��>61N�q0+���52�{���e0��� ��y37�%;��[��3"h�GzY���oPOC=O�$���zq��T�������ܸ�Dp�i��pN�y�*x��"����b8�B�ŏn,EyՒ�E� ����x�v[�a�����zK Ë	�;J���@���EՀ�U�ӬįL&�4�DU���-p*5�uo%Z'���|����:$� H5;�N��e��F��Dn��Q�K���0��.vPA��)�L��-y��S>� ��"aë<ǺFIs���QUo�}�݆ȸ<E"� �?W��I�t�><���ڂ���C�ܬ�`'�gd�'p;�w�%�o��#�uNg�&���W���I������hb_�QmN(�&�H�60��|`��Hw�SΠ��r�&��y�Z⑺��������eֻ�~�h���������|���l���9$A6a���Y1Ē.�:��R��&�Ia��b�"J7'���%���ҩ�#	�M�|��JO����\�t�!	p xf�_A���|�F���[w�,��Y�;Tm���d
�dE@;q���������>����h�M���5�e�h<����
��|1@D�N�N���tӟ��G�?�_B����������n+�X�}��O���-^$f��o�5��*G=�O����:��i��4�7lR#��T�0�f["����� �������(�Q�A[�abM�w��'9�VR\�/!	§�{��p�^9���l�����p�e�"���ÿ�֬����f�͏-�դU����N9��V�y��h�Y/���׶L�j���)��у�l@���a�Vę�b��Eo��Hm0�~�M7��Oч��H!��`N�Tᗇ6ѻ�:��7���1�|�l��}�*d��3w:�[6���~�_=)�a����.s����%���K�	vB(�zv�oxE�N����S.ǅyƈ�h�kA���}���2�߂k�è��ٚ&����a��4_�W�LLtM�8R�TV+�'b���L&_9�)k���Ͱ�f .E;ע���Z�7�z���>.���g� q
�"5�wH?�����: ��a]���@z�1��8@Je�_y�����7��t^*��J�==�����R/�q!|�������Dqϟ�R��;� #1�Jm����iğ�+��cَ�8H$�r[E8A=�'�J���W�i��	�p%8��M�"p�шS�\u�ٍΊ��|k^H�[��V8��ۃ�o(�9D��|>�-Գ=_�Z��G��:}*���#�Y�K%����; �!����
煙������0�b��k\e��8#�=��]I�[E�(�&`j`�c��ĥ-�܁�]�,|F5�0�DE����(��c��3b��ET���Y=��Wx�stm�T-��̡���ba#@8�1o�qd��]��?9*�[>�U��y(L�����X֗��V*�ݲ5qS��/ ��0 �SW�*�,>�Q���,�ٳ��j་�o|�E�6���4�1���hDk�!?����5�.�-�N�J����M�e ���Z��t�LK7P�C�����vc�����lI���)4]g���%��"�j�x?>$1�B��~�N筒+�	��D��\��v��vmU@���zS��Σ��[��u	���v�ϒq���jM���9F�������b7�5
3Dny���2vΚ��kȅ��^�'���<9�l�C��86�ձ\j��2>r{<�e�!�~��txT}��F�Q�Y�ێ��h��úq�Z�f��r�w�<���$�&bL4�o׶@�r��[h*�*�&
0a���^��[�a�_������i���m���$������d�	���7Bs��igN��,&��6����W�J�$�dzTcˑla|]�F���&���0�d����F��d� �����r�J�����Wϊ�	|8�7�Q]��a̫����ʶ���\�9<��o�R����g��H1��_�1��I��Qa�����y���|7tZ�υ+ˉP���֚�����ӞU{�@[������x�R�����CK}�+��W��_\7�.1W����p��\P�
� �e�^;B���1�K�`�����^�G���V"ĿD5�F䏝L����,���h�܀r�~��[�\�4��!�`�x�c���q/q��8=������8����W���i�z��Qqg(
��^5�Bm�ܲ��͠6���I�ӹn���N�쥒�з���'��K�����"�[7��i��J Sg�=x���su~?w�+|dYT�/� ������DBZ{�3�Je~t������@
<?��K�;��b�E��ݭ�V���&'1eP�Ww�ҵZ�k����U?��x�������Ķ���w��M�vl�1`����H���f���ǭ�#���a���m��
x���F>�*LQ����ۼ5n,g��*�&r{KW�md�@�J���'!(2A�ޖ���ѡ*�Y�)�ݤ�J�$�\��hJ٧�P���9Р���dX��&I;�]�:�)XP�q"�i�rS���g��1�� f��OA&O�'�6(��>�Q� 4D�~����i.W*ĩQUh�<>���F�=ok�������9�Z�v����e��=��� ���Wb���s<Y̊�����hS�'�+P�d��B_��l�?��� ���.���	J�c�6$��`���E�]GL�ͿX���#�%�3;X�ABw����C��l�����4}�[�ļ��H�`a���7N	.̐��V���}��kV���LJ�k�`+��oq��Q��u�3�}a�ק�;���I@��(��E*IEj�U��N�{� �q�6��A��X�&�3Q6��4�S�P��Ź'�����r	��c͹so���U�}����WoEY�"'^�۹��`Ҏ�x�����h�k���B_V�r��mFKz� �����lUT#2ױ�6�X�AU�oF�!B���^뀾P�m�7H6�Vi�G��ʳ��m�]i���&?ي��>qp���M��\$�hR�v~C5�?�=C����RD2r�	�]�6�� o�\�+�$[���A���s":��+���.�}���Y,��t?����6l	�P�O�j��t~E`�~�=�i4�P3��`E� 7P8�$�3	g�n�@���(:�K8�v6����)|�0*wb�; �]��^Pir[Y���� ]+��<y��!m�A��\t����;�#ZN��,�w$��<ob�?i,tĿ9���p�v+�i�ЍBկ�:?��CPF`i$m�M|F��}|������A��gT�hS(�qYZ�pB�CL㊫�ex�_c��71�c����
�swE�I�+��L�mS݌'���c�1�I��ĸ$�J1�B�<޴r�}��}���(	5�;�[`9djª�]2�.����`�bG��#�����K�47�K4#C�-|��^b�~�h�pL�qkZV�8c�*~� q-��$M�^�"�F��2�9��1�Զ�����~�Q� d��aD�&�Ie�7=�F��H�Qn���5���3�a�����n�n�l�V3��T��Q�L¿s�|���:����"T�o�*u6��'���vu��+D��:�e�3�X2��(H�nZ�ODɀ� ���@����=�8�X���ڞ�i����
���V�?�_K����nEل
�1Լ�Δ4=�q{�XR�:�^�{Pz�F�}�X����r���0b�����9����}+b�Z��.>�랪�	�4HK��c�i����h���jj���J��*P�a�.�wV�|�_�<���RC�����!��l(����@�1¦�т���xy?�������#0\��HM�Բ��j���٬��!Ѓ�r�	L��mB�M�i�
Ԉ(�����w0�X��>��(]���' ��o��G��>�"/y�Љ����<�;��/P�Dfpó���|���w�y`+b���b�v9��i���I
��ִ�z��|rn�Ws_�A��#pJ�F�|*p�T@[_7��gNӒI�����1��%D]�,�����z�4�n	ƛ)f�@FO�	�M��]���%�R퓿���ܶ���C�u��tY ?_R~��<�0z�M�װ��38�a�Q8�3�(>�rO"9j�y�쒘��z����j�Jc���}q���C�d�RC��G��7��u���j��RL?'I�dS���ݭ���h�NJ�d��'��r�����W=M8EHfʫ�Jk��D�, Ԑ���:��mg���/�Ɔ#�����V���!]B���PJHks��^�5�3��m��~��\ �H	l���5+��q��4��G�����ь0�c������P���i2�E���;	}��gN����uGQ��(�^�;4�iA�P�P|o���޺�����ά:�z~؀�i��cf�&aAʥf���b]>��aX����{�~O��nF"4��9Z)x�s�U}Hu<����૟�00�3ʳ�d6S�'-T5������w��T�̀~�lP�y*]K$W����O�b��*۾׍B�3ڇ���t�ǽJ=!���y��%	 [G�c�4��	�%�P�Ɵf�v����ã�.ì�f��D?��e�>,gÂ�d�	��;���f$������A�]Ҥ�NR� KIw��Yڄ���$ϯ͋m�0�t����#����6�Q��J���I �	���1t�x8�m��\�{�>�xk��Ր{��NpS�M�=�i������^��2̼�U�X>k�#������$r�V�M<� ͅ(�-�}�H[/���5����<S�(<9\��W�9@Ơ�Y���^�}��ROěEP�u�H>�8�/	<��zߥ�ڂ���|
<Une�b�ԗ�r>���i�����D�ݷoӎ-P[t��"��;��ʻ�ef�j�L�����#[6O0�mb륅��U�{��V&<�_��)�G[�Uu+�����V2*t�|k��a�o����!;@w������0�

��@746���zr���f7[��GMZׄ�S�3��"�S��z����bӬ>�z�&�i��͢� EC2��w�j\ZhD����MmT8�Xа7���Ц9����K�*�1�x�+-�E��$����=`��ey܊p�ӎO{PA�o5�L�[���;yN��'ů��$�ÈҫW����Թ���w%nŇe(��Ug�s�����M�}�"������͡���!��c�%#}' �I�N��_��'��M����nh� ���#;@0����Ľ�HFh���o�B��:aŀX�L:��hx����4-�oe�n��U�]tZ%f@����B��^+�I�jm �5�*`m�R����3w���6'5DG��vU�%w�	��Q���-}��"��e���*5��`��A*�h�~/�[I
a�<j��!u��{po��F?z���֡�g;a�[�Л�ߘYy�?�ؚ�zg�_Q�16$!���^s��x�9I��&�������!�P��DE�:��1q���0��\m����7%�eUB[vɖo��W��u�/�+��q�Y"�Y���7+;�מihA�J�[�n�V�i�XqF��W3�U�O�qI\�7K�js���T|^צ���ڻ�-ӘN�/�3�����[
���N�`�`s���j�~l���Qvm���*'BC$�n�#����fg#�n�����Y��:TJs�*J;�'���@��]>�g�2�_I���O����itGډ;G7I��^	���V)ĕ��X�Gt�Ocm����Ɏ�A��5�|������?Q���U�1�I��Ń1��c��g�m�w�x�R�Ӽ_bX�з�<$ ��(����l��GJ���C�R.aKɤ�e��{����� ��nζ;j�q3POz���z �H�J�7A���z|h�D9��,Sΐ6�2%���}�r���޻c>~�0��2�e{�s}kd��A�$�-h����[[�����6��T��]1[�Q�o�Z	����ո\���	��h�-[�)K��F
�X]�����UxJ`k�`k�+�M���f`�$H9�X��Y?E�Ib��,�5��6"]����p�`hD%j�3۳�Ӹ��&���0�{Q�q��NK���W��:�X>��⮸���A��	L3V���7�ȑ2De�$�9K�K>��b�̕�j��٤.�)����fX�϶�4�<=*m�&��o�؃�����&����o��nN�q5aW�H]�I5=�`Nn��d��6vLwz
8� ���𱄪߈�m�g��q�}���_��}�vb�8Ϳ�3�:���:��A�	-�MM>�@�dZ�q?V�
����D��+��,�~��~�gQ�v�%uel Q�"f����6���' Dڥ>�P ���>��~���@�5�Q��%rސe��.;�	�7Rͯ(=�	�ĝV����Cű�\�`+�4���EAiZ����,�pc�sk�]�9UJH�m�y�����8��A��tmn`	���c��C��67�[���YeJU�C��/��b�)���7��q<t�^T] 3L����H�K�f��vz�Hp�/��&��i:q��%�K+������%�)-�<��9g+d���B����S�1��"�i��K<�!p�6#�[���p��gl��ô�q=�������Re�{?h|����eܢ�����������3WǍVx&�� �!�t ��2��|�k��d��N):���H 5����>a���8���\��%+7u�N�%��9�+�.�ݣ��j{$�J 1բ�>�_��*���w�Ai�HJ����p&7g�1���-��>�r'�j*R1s�.�d�'1��m}�KY�I����0K��!Z_ E�Č�f�%�ߔ���W�U>�_4�EK��i�.������m� ���౔<ⷌ�ު0lxV^:��V�����(�L�f�`'S��7ɖd�@\��T5�c�� ����:�"��}~�¸r��$��'��ʪAad��'pU�ܰ.��C�!��^�7tnxB�16k�p�X����FD�F<���U=��.ȓ{9�G{"�Ln�3��d<Z. ZG,J�R���hX�������/�N=��I�'O�ݞz'��t60U���H̜� Qm�Gޤ�mg�-��&j1��m��gk�>�~4���i����e�]H Qc#��\�A�;��Ց��-z�폄�se��^'�i�IdG		�}�O�Ǝ N/��/�K�8HI��di����g���c�.���!>�E0Ӊ�Κ��+�*��D��SW����u�_νq�E c��"߁B�Dt�UP�v&�����X����/|�Q�&5��+���|�-hD �����'}D܌Lb��ˈ�%��@l�/�͈�@��ş�ɦ�T�Ļ�1N�.^���Oa��K59�Sr�6���W�Q�+)�a���^�d-Hw�a�a�ڍ ����4P���$=��9�!�q:��x_��o�vS�K�.q�1E�ȁ��O�@�Q�:�x�i�j?r���.d�+v�?)�o�k�?51��5Mn�庯�ՙ�����۶����k,�V
�	u�M:ù�ɋ@Y۶r���6�s��T��I����Et����z�1�m=؊��EU�-��ߐ4t��� �k�fB���Ǩ�=������1�=�mzx����§�('�v3g8�X٭0��C�r�|�E��hյ����� �t��o�D�\K75H��B���Fӑ��s�LD�������������AhN�T{bS�E�̳m*S�4%(;�����o��*�eR�P3U��F*�`�y�������z�������ѵl?�g|ֈ96��I�}E}4C��y:���ʪ�m$��ѭ����!s?MXĹ�J���4�u��*5$�л���Ĳ�)?'	���ò�3�\�Q�.g�Y���ić=����b4V�p�D����m��q�å���u��b�ƣ}�.�8�w��;��Er���C��R�X�����3�\Do�)��T�e�w�Lp���:w�`3p�v4��`�x�6ف��x:�����}��@�?g~�]�]6�V��!dH��:8��'��Zh���%O��G^U�[��R���:����>q�(^�`t����S�.y�j���S!.�:F����m��0���Z��,��4���R6��6 /��s2n@���J`H@ ������Z��<RR�RC7�l���vu����Y���c�%�#<H�)V��y:5[�>u���0擉�)�SΘ;��F�m.�[V���qr4���/3�oqA�'����2�TP�]�Q��oq�h���(pj��e��;�@TTvr�L�hy����01$]�4cu�sl�t+�����"J��߷�=h�c�̒|�I�6;��%ؘ(���2�i���hKt�kyr���.<���#��7(��A�Yݨ��)f��;��)CzKhÚ�8�!Y��܇,�YwF�s�E�Ҿ��5�.P����5�,C<9Z���U� �^W�c3R�F�Y�Y��J~nq.�=�k-�¨>q�{��Bc3�������,��%��.��?&Ts�$��o<zFzb10�![]bG)����F|���C!���[�3ܹ�V��n�L�m�D���{jcKH���s;Sն�F�֢�L����38�V�"ǾF��8�c�IcC��9��%n�b�+	P����c1
�I!��:B�F:dk
7���(�w8�6Q�-�i�=�ڂ�}}f�`�����l:<XȌ��MdT��Cպ�XD�o��}�w,��Z-�`���L�]���A��g���r[�����"���i���M� ���'����"uu�vqg���Y�hSǖu��ݱ�eԗM[6ئ�ǟ� ��J��厎C?��s��@ٝ��xa���HwW�y>.��m2��;�W��+,�;.�Z�����X�-�[	|�)�S��Y�9����7���<V��`�?hB�0Ʃ�ٵ�ПO�+,��o�������N�A�(_�M�ڦFT�K0z�"��V@3�(0*���w�DOR�ש���"�:�?�?ּ�a�Q�)�/�v�sO3�F��jS�XSy���v�3u2$�'�s�w�-�_�cN�Z�g}cLl�G:B�HA.N�aj��E9�g|N)�P�$�F��*�_�V�n�� 	�uf�v��t3�,��*��+^�3�hAh6��{��c� W?��h���(����%�������4�߃���$���H�x��3�R߼y�i`L��:��k����mx)j�+�zK�R!Sį��g���w�{�:��ă�S�W'h
��EV4jM�yخV�ۺ�Jnk�����7(�t^՞�e���?��%�-�ń���l%��o�R�@���uy��DC��S���	�JţU��(�u��*ϴ��I|��LQ��� lhе���L����,Px �DY�.�Q;:�o�]�YzU��A�Y}���[��b�>$^���v�b->�,,.͞����ϒ�/�������ۅ5Fa�I����f%e���gU�ӟ��(�H�8m^�tN�������� &�W��k7��W�+3��c���#�ke��~���^�2��k-�?��1�������{�ܰ�F�.嶐،�Xx���S�[<�|�g�l���J�3Pm?ٯ������flۜkF-ե�;:��J�5����vCx�/�X���;D�Ysg6}�#�~Fk�r����X�jε2Pt?�?bp�oFբ=s��3b�O����\�T��A�%�KX���-�9���5���b�>Y����&���H(Jh#D�D �2:����Rk���JL�D�=��j��|�������$���Dz���?F~7�o��ٿ��mg���p>␆bJ}PL�A�����������ꖼ��+I^��	d�� F�]�m���x�J��);��<�z��!�P��u�	Y�s�?3�����?I�c`q^͕c15��Q���vx${R�O7ܡ���-*=?�L���QB����Q��+�5�2	���,^���\�:V''���������{�k�s	m��@�ܢO�^m5�(����
4�w��J ��Liʜ�_�kuI�[�W�D]*�ڿ�d��.�Fqnߘ[��㨪�{���)���J�X�-":/!R&I}4��ނ���ގN;z�jnApm+x�@��7�T��K�a�jң�sj� ����`E���p������/����b-�kT㷟�KcDdB�����]/�4�:�I���*�G&��v�pO0��b�I�a�lL�ØtM�-���$��Po���Z	]|
d�i�F'�-$8�������=Ѭ� �yť;_pוV�{z��q9���r|�S%:�SI��4�s��o hh�;���r �0���x��1�Mf�D3z��t��+�d�B�U0Wo�,�}��J��ٍ��@
<N������z�p�]�|SѾ� �>hm��p
G�ܙ��d��E�{�0�?c�n"� `��	�-f���u0�(p�0���s&�g�S�&���Tb Gx�c|ZLz��є��!�/&�R��y��V�5d�G��N�C�z��<�����?��� �����������P���.L�L�������'lZVpLf})
��JR	->�b��%v���(�d��,���Q�eD���pLHq�q�M���\[�w{ݏ+�;`��:0�{���X��yF��E��[͔��/��f�����?nd���d0�"��)�-���#�UqQ}����K�ص
�IWd��į�F;��g��b��� ��J���Io��ݯ���^k�6rۄ#�.g�����*`���C6������^^�� ϢOq�V��g���|;=.-�zʙƒ	�i8�u�αDp)�0�F%2�ԩ 5 <�XH�rm`g�|af�vb�f�g��hZJ�{%�0��J�{&��TN�&+cQ�*����z��m��u���sw��W��-�]e�pӖ;��\\Q7掆��|[���a:	��'[
���;l���Ն�m��^�m$�d[t�3����R;b��;�(����G����A.~�*[�RC��P<ND�#�G�;ޒÑ��MgB>v.y��dқ����Y�j��M$K�t*)����l�;ob��m�t�=_���.��!�)���BB4���-�]��V�B�U��(����\��q��4�T+�N!�Q���=k�2�[��l,C�D*�<}��L�K����_ȒKS�6�V�����J��ch��ЭM��~��ȹaT�ho�n�ս>7����N�����oI�"Ζ)��Mi"���`��n���I�!�]K[�qz��r��QV�#��3g��+t����(����a�xk�p�^����v�c��.��'���6�V���e9�n��+��j��7��5��]��g��Rcr�B�s@|Iw�yJĀ��}ot��<ꃶ �w�d�d�.ݾȠ���}+����v-g�XAi.^�������+b�B�1N|�Rp���h�v���KR��V���qL�n|�;]�^��%)QD�6����O�~X��X�E0L��L�d3?e��`�y#Z)`��!!~vL�+����)�e�v��[�����x����O0�U�q���*���ҁ��8��'�4ۼ���I��`�[�e��(�� ��O	�r��R�EP+���,~𩉬��%���O8/�jt�✆x��s���5d�',��O���"�HT�����F:@^,QڣG�s?;�H�V�(A�8�B"�m�v0&��gB�����-!l V�|�hZQ%�3�����tM7�i�-�csu���
b�:��+���w�),^w�I�&qI�^����_�W�έsǂ����x4� ��ꬾp�����wB-_A�-u�5�^��)���k��c&�k�M��ӨJ?vOi�3fR�����8�����0����]3��Oګ��
���&�n��@L����fD
���S�Ԫ�$��.M����b��5�+���縟�H�Yy	�f��k`b��i�O5��'�K�������I�R���WHX6��� ��8��Ň��Q�3�.#=ɾ�T΅^����u���O�Ӹm�;.�d�1�����;�=��ɴ����$���W��jT�o�ݾ�h"d���xmD�-ң����[�u��6�Qz,�,�5ř��Dnb�)B}I0�'�T���׹�M��5X� I1��P����sSd��(��B����9�{r!��h�u}qh�FiW����.ʋ"-��'�%Շ�yc��	}�T?��7��� �/����3�}��<�^�	��_d��B;-�Yn��;# ����+�����`)�ԣV��صP4��0��[-n		��{ז���n�E�M�H<F?��g��h���|K�qS��zI��s���=���+&�g��v�p�#�z�8?'�͸�� 4���0	�����;��FA��	�c^08�՛'0B���,��8�>xc�B2�Ӷx�ho�������xS�sB{Ɋ��>P\x���P�i��0����_'���G��h��QK�$�R�Ӏú��y�{G�ԙ�qchF�jsz�7v!hES�:�Fzl�K��"I��VH�ɸ5����9BJT������Q6�H��YK�B�q���Ry��B�2�uK�h�4��m�{��<��І�8���0ll(�F����zTe���O���ӝh�"�r����[N��]�h�@QOh��Am��u��W�ʒ���T�~9!T!�I�O�E�s���L�@(�R;p��7]R�)����O0�%�{:�Or=����mz@^��m|����rY�F���7�);?u��O��{�M9����^U���%��f�~8�z�����A$�W�h�nT���`!K����-�`^i�<�GuM�p�y���r��Ă���1.��#�j�r�r0ӣ	��a�q1L��I���-���'�-j�-�k�2���#�����Ǯ�".��iv��_�K��O�PPɌY� �} k��  1�9������F�7W��	Rߛ��9c�h�E4J6L�1�
�DQR�6į!Pפ�J̽�O4k��@+�W����h(|��4�V��P:e��Jм���%rPv4�>؎���njz�^���G�Dʑ�t=1�t��i8��$q���Me�L�7	5n �ﭐw��m��lM�;(ƒ���Sؙ>�Q�d���D�"�5��˱��q�#���T L
�MZ��+j^o0a�<.p�������ײ�x���1�e���C��~���h�)׋	4\�����R�C��Og������|/~��_��T�
:��#�/�@�Vq�L>�-6����B!��YkB-�����(�-��_�QK���"G!@X�i4�B�(�:u}�J񭡑Γ�h�h�2��H�/����@af��d5
�+"�qmƷ,�Ĵ��mv���}~_�%�ki�OL2[�D��N�%	�9
���JK2Ɛᜏv��<!PiM,�>zL�¼Ci:�;�~��z��ޫV2>�&��͊��� �j6"7}�G��3�/K���;�[����a�0��Ϣ?R�(z��YE���Ğ!G<������^�����0�U�y���s�֙�!���N�6]��# ��+��S�&��7^����tڨ� �htB�w�� '���F2XA���>k�;�����լ]�¾�Csd8�e��?�S�3Tw��Ǹ�P�"�����à���2��az/W��B�b�ʖ	P���d����9��z_[)�j���gU������E�V�zK�=V�@�I��k��A��[?�C���Ѐ3�^�!��.?��:@[�|o*�'��yecb&"s��/��S̜_����;]�a�U��B��;���a)8�a��(	�-�bss`��;�Q��ojb�C�&h�6�۴��y ��SG���a�9ֻ	@�i.�(��)�+�ՃH.3AXg4�'��k�&sk����Q�׭P&*�v�*�;(?Y��Y��b0��G�0���q�d�z�V?om#'Ô0Ω�H�oxQ[p�q���.�cp��C�FɆ����T\Bu�������u�no[ej���iO_��&����%g.1w�t����
x�]��  Jt�^�Q��!H�k��M��P�5�p:a�H=M�ۤB@��c$E)~�-]��Xr���ƾ-�l�Kģ�?�!Dh�g}c��n1��QU�t��01��;��B�
�{��f��U:�-E����:�����r��۳���-�?�b�E���07�;����Jjuq竔ثJͲ�Mh��F�RkC&�b+��'"}����0?�m���K�dx��?������.l�����7�i��fs�E^^6�=���ٓ�/���?�T��m����<vhz��B[G�r����s]8�q c�1�x@<`�)wن8�;�]kO@���x��<X(�Q�m��ri�|���r�Ė�Wj�:ߘ[��<�rT9ˁ�QR�_�� �F�Z���}~Yr���"�=+�m�����kpT���H�Gw2Ds����i�R�G|�n�R����vv2�3{m���T+��W�)ϐ\�| �Lܟ�bȑ���_����o+����rA�ǵ�X�F�,u���S?|?���퓹ha$^tA#���7��ꈠޗha˦���h��.>��<�*�>h���,��n/�%�k�qi|z�Ϟ�FV�~:� �l!�1�@�o{v:�a��%�F?�!��ly~��88+�6��yXE��v�pR~9׃Dr���w���Z�[2$Qm��
)��l���n�Ox�K��\�Õ����;�8خջ	o�Lʄ�}�4ޅ���I^yu�-k6�	"�D�hC_���R�#:��X�1�dR�e���P��������2��m>˹�]�"��zNҜ���mEE�����f^�PݳT�[���\C~�/�/���	�]!�.��
��_���U�������~����]��Ӛ:�����(��֗"�T��8�����m>���?��_?=1$����
��3M���ݲ+���+.8~�.Ɯ��!����\s�(��c��Ζ��`J!$9��œ��8D��r��=���|�!s��x����`�UV�AA���'�EW~[���SV����[}�=�Cl�If?)N�Ӹ5��� �7+���ߢ EB&S[��M�,�ɽ>WgR+]4aw����r���J��Ԣ�"̗{|"�-�'������<kXj�:	�e֓��7N�W�vjI��D�
3hi�3��U��,��a"�	��,𼾹�����$��WcnK�p>3�N|���ǋ�Gc?�l�$�X��j �dZ�fxZ4��¬a��V��M�Q)'ᘊ<�,sθx=��c?f#H�4;�z�x���-��k$j�%w��x���\�*PM���H�?���3wkG�w$��r?KnF���z��9Fӈ��khO�y����tȫ7�L�9��-+1p��8��$�xDl[yغ���P��,N�2w�R{QO�FZ�8x���5
������8��[*�[S�ۿg@�����u�h�B~��&���H�+�u80`�M�#��j�����-@m�s$���� 8pΚ̓�3������T5�	m 8j�_��A�T�=��b,rm�;L=�[�:\�l8��q�.|�?J>y�U9y���NH�idـ�Խ��c`vuT��H��h!���čߝ�{)o���\��wR��)x3rXH<���˓�����T�f,!X���+滥ȭ^!�[T�&{k�fR�>r�j��D����}Eܼ�>S+ h��e�y1(��<dyO$G��u�n5���!N <��Ui��|�b��Lb��'%#��I��l�����p�A�aU�Z_�r��m��rxnj��HU}ێ�r!g���bx����B��Љ)Jf�eb7����it���^=�YC�7�4_D:^�5���T�'"`(O�2	X�NX(�r͚���ʹ����۟b���ȼ� |�R�}�P�M��rQ��Z�9Va�@Ȯ�ġ��y��yh�ꗌ�Z0�"1���&h�8(V5��e�u�<`�eU���	�h!�+���	�-K㔆�nr�i�~��;Һ�
���Vj�a�^�j�b����\�A���F�N�T.:4_y(Vߛ��ʎ�>H�[aqk�v���K}Vk7��z�{^���jW�'6^[q�&gA�J��"dF���*p"G�d�X�����/cuYeT�X��B99"2����>Q�D��]]�pZ�<��n���'����b��Zf��?9uQì��@>S�!ɂ�G��(;�\e9����cj��:a
"F855�Z ]O�3�raaP�����tǸ��{�6￲4h?��o�Џg=l���[�p42��Q��En��LB=��j"[�#�Ф���F��(]������r�K'��'j#�|IT��փ���H��A�L�����Q~I�,��=����0��5����f:>La�	�Q�¯�HQf=��=� jZ1��<Ks��;���s�<����F�k=-����2J����+�L����[����u�Q�XM]GJ�B�H��4 ��m�;k���8;[������\-���Odf[_��uI�2B���P�]?	�p:�o���*��q�SqZF"+���=�
Ru�z�s.7ҹpZ����Y1�B���N�v͓˚�X����@�58�k� ���\�+�U�v]����&_�O����`���Wsbs2�KŰJ��I��m�QQ�(K��ۤT��%qC�$�`��Ar�Ü�xF{.�i� ���KI䗳�b����
�NY���.r�n����8��d����F�j=�Q�y�h��[f���CR#��t[�j�r e��|F�G0'=a	o~�W/< �=���}8(E�8�� ��u���ܤ����i
�D#Gd�~s~��0�2���=��X�C����_(���ܸ~+�Po�*|M0k�և�V��n�!�������`�� ��K����F�u$E�t��(�����|��e�S�L@�G�wF��oV9�r�*�<�m�1�[�V�=f�ū���C��A^q�t�{ ^^���9� � A%�d.�]x��k�tI��� ��v�����|E.}w;�x���Hh���B<�+�R��{��;��zđ�72����W,������+P�K����(?�����5M=�S�yGX�Ãڬ��i�e��(b7c�T�=W%*�ɒ׈�S��
�e�[
����a2�]�@.�(�<">�f;I��*��bs{ot�3[.-c��	 OQ&�)Cfدڬ��^5!un�>���j�]C���M�AC(��̐��{�Άh�+2*o�X�
�����P�zteO,gfc{� &hP�����=RX~���j>��6j���ʬ���ޕ0ľ��p�kpw6�e����+�<�c��o��!R!H�`^ٮ�8�P��i�=@,*AK'�v�.�Z;�?�0�$�0Ha���!=dXN�a������T�'h����J��G}w����}�c��k:�vt�@����a!=A�gP�Xg�����s�گ�> :J�UM K��*V^t��0z���;}��r)%�Kt|C��1�u��I����k�.����&44��bJ;R�\�.�O0Rٽݺ���B����o���eG��w(���{"k�E%Ǫ��A��~�ת��w>�q���D)����<k ŕ��[F�'3�GqЎ�@��rǛ((�۵� @�)�����wb�'�_U��$��$і��pLn=��c��g����^�j`+Y}ԇm�#|�#X�5s�-�e�@�𓄉�oD�����Mأ��|N� �$m9�kp�����(;L�aP��"�	�L�(#x9�R��H�|�ǜߨ�DD�c��w�Cl!�?��yn��AB����W���� 0�d i��I�׌��*G��(\<�17�?$��{P�� �]Ǹe��Jk��DE�y1�����޵H��9�i���.}'WxA�Y���a#�bc
����T�O?@$�$SH[�Y���x�{V,�Q����d>n��~yJ "\F�AÆ��j��<fr��;��2�V�u���w�x��_�}�Mn&�����v�6̠������d-홯�g����!��vP�[ISBKВ@
���"Ke��Ë;$��Q���i���9�ޙ�D5���;���R�Ci阙���mz��Ce���s~��Ɛ��$�����O�$�t�� ,H#ϳ%�'��?��`�M�#$lw�;$��
� x��r�wx�(�v�ۥ�K����(݆�C0#�x�7$XT��I ��/�O�D���g8����f�2��Ǣt\n?�Y�슘�-�5r'�p@��sJz�@E�=��v5�8I�&�. ��[>��3�IM?��0�<p#�L+���j�����N_f�m����x�ÊX��#�����`_�vGi�xC��(�ʒ��e���?q\�&�󐘨t	.�/9­؝���1LV��z�C��7�_X"D�F�m��J7�b_�*N�zl�ד)�M��M�й�8�^��>�DDۛ�;ce�`���33_w6̛?&�h}Dt:��\�7�Mn�;����:�2��M~Ku��'nHY�Z9�7�]�\�!�<:!�<;��!� ��ö�Ǭ?ac�&�2G�8i���Ro۩Cߑn�Q�4�G-�j�g�V��S+ۓA��,��6�� )�C>$��=Χ���Xݨg)���,'�z�,��	Z&?V(`� g߽�CW�`��\�˴�6�J�O�V"Ӎ`;�*��[14v�S)�D=Y�>��ӻ�c�(��4"���M� f[?�bǘ���N�c�XvK*�ӎ�H��4�0����0TO��c�)����6n��-�}��!�ً�^�8��#Q) �f6��Xv�ё\#�aW?�� �>.N��Hhr� �����f�CJI.|7�An��EN�-�C�N!�g��\��0��Y;�D�t��t7�Uakr
g��# ����������0�!����0�gz쏴3�8{�����VG�Go���a|��i���=˦�W`��w9` ��9m>O��y�c��%�ڐ�q ���*�Ɔ<�����[�hf�w��$i��2�B��Tt�����L1�ri��JD��GvD��OY��T�]����Zp�:�T#�N1�4���Cw�]#�\�K����2�s�4 �������~Ï[a)��k{u(�E3}[{5�q���W�Ѝ��?�B��?a�+�Y�����؟�9[*z�k�%c��$��޺�� uC
2V��A���E��-�Ɂ�Ջ���?�u�j.��,h��
�2}�%2jM�7�a2�N�H:�Z��ӊ��D���3�������]F���oJ�b�2T3P�������<c`ܦ0:Z}*�$vn����C��2FH�\�ʎ�}�c��&�̧�#��I1�N��)��XBp�ga<���c�$�8��}�
2P_����-�(e���|��CF�BV�G���.�ZrI�U_��v���ҩ��H�)�NT�J��3�B���p��*�u:�ߦ�y�"�׮ӕ���%�g�"��3���Xn�=�x&�ט߄����������4��O�#*; �9N�z��
�{��˙ݑU�Y�̩og�������h�j�Ħ�(�Q<�U�gY�B���l����:~�&}H<o�5;[��@̷逪� �=:�����ӕӹ���(��t���rǩ���D]�p
�#l�H�4��isڴd%p��ĺ���D�-A��Y�o�@��k�e�BW�귡2�Pm?'Л`���f�Ş9͂ؕ�2�Ks���C�JBP�9��vـ����J�A�o�} �o9�项��!�w4(�0��Y�0�xY�۲�K	h}ȁ���U��>�K5�A^:�Z�u��*\9
���Z�u-U��y����I	��	��Fo?�Z�ʜh�dQ�&���|�`�Wn@�yk?-�eM/�-���w����b�Y���u�|�.���"9*���r�i˜�X`Up��կR:.���$�״ ��~gP ��ޘQa����nr>	��~m���)�	��0�E�1�EI _�ɷoA<�i���&Q�:�`�")��]�9��A&J��Cwb9��.|�C+�h��G� ����(�3�:9�=&�:~��/���g�%�6���Ë�q���f��"?⿂F�%EjRJ6b�Aݠ��(@���l�l$��'3�Ď]���M�lT�HسF?��A���?/�"�~�?HF���?=��A��J�f�S��%ҨX��:�� JG��&J�ۿZkjܙ|�?٤�s֚�j�����*���ړ��:|��7�J�8;q�r�̟"u����Y���1��D�Y�;`E0rZd�"BBY��M��q۬���
�0�*nH��pZ�N�#=��A��|p��g��'��\���~.�ޛ �*S�V9���LB���	�C��/e��o�'��(m*B{n>�"V`	h�G��}/f6v������{ \C#��6k����[D���}�c݊=X#L�e��hNʅ	-���ST>�|�$�����9��>_^��~+m�\���Y�M���G~W��T�9�3	u5�OR.��o�y�u���u���
��Lih�Ch�����ˤ��&ܽ�Fc�K�>/@ˊ�A6��*&	uA0��V�Q���4s'B'�`������"Tl";U�7��P0�B��r��|��u����9V��K����2L���������5��̱͠�g�7'�C�z*������iӟ,�N���T��f2�t���Ig�Z�}�Q�i�e�$�=,t �K�"���)�&ķ�;\��܍ h�I�9�,m���{�S�ȚhՂ�fH�@�h��Cqr���q��-�y;�ӧ��kDV��tY�a�ۄ�]<=B�Y��6�K��h2ɂ�p���k8 y������8�`�Н�Y��)
�g��n��S���*%��bMX�Ā�X��W��ئ�%����@{��P��a#π�>M��z��B^��N���Wx#!5
�z���ﲆq|�i���e��ZCnj��v�����Ƥ��n���S���]�w��E�]��V��6ܯ���W�pR��s`]z,]��f��>YM�a�c3t��a�}'�����t��A׉O���}���@5��n����`��;���^D����~hE@�áP_�sDԢϊ6�$����|Ї/z0R��TQFk65�6f�/�LNK�@�?S_��o�����O�,8鬶s�4<�)yB`������2Z�������ު�@�*��Iaɇo#�aw���f-�k�,K��{�L�{�k�q��N?��{e,�Ɂ����5�K8�{��p��Ih�X�9=�񷯵�2w�(zs�^��>Xç�צ�)�B����t=�z�v�j�3}�mӠ��~�/��@��ĸ�G�蔘�ķ(s�;�n���;ɬ�,�q�d����`�<!}0� �y��\�����mzL�B�^����lp�b�����Es�yBK���o�7�kۑEj���IJUpiD���v��
1[]�q=��o����Ք�t��*<�.�^s#_n�T�z���0����GFÌ�����{D��K ��ގ���k!�PeG�N=�u��ĕ����H��������D:5�O��ZP��e�hKNH��ߋ��K�f�`�Z\W4�_U0ULv�;�̨`7@@�����c�,N�qޖmy�|�K�6e ���E4����ML�|y��2D�4��8��	޶�����a�/�ט��˜O�d��/�讓���D�]�]EE�gh�T$��������6����H�$c���2v(��"��oL��K
!�lk�S.�O!B��'t1�I��:�����_�s-$G��d�3M��8�LB.&EAk��-
y�ܟ]�h1��P9P_=G:���TV�����ej�D�Ϸ�g�W���kFD��2��w�9r3������s�%�6�K��I8�i�ʕR��J2��5vvdk��s��Sz�e��X�i�u�ʯ2��HU�E`Ӕ�-���i9��+"�#	��e��ȷU5slq\�|1���)Sk�}P��f�/�w���P�PD�_	E�a���GfZ� ~8��,ܺsn�o;��%��O�ǳa��y�(��4�B�|٫����/���47X�t>�S-AzQWԉs���8�<hz܎�j��<���N2#z6b���e��P�s�#�c�Yk�F����b�d���d6G�B��a��� �;Go|�P�d��6Z���YT����Q齚Z��E��("��YI��1֤es�`9�"K#��[P����W�O}��)��YQ*��A����}��$� ��Z�SS�����Ӎ��(�J�����D|�_���E����M}��f��Ǽ;Q�Z��8��#E4lٍ���/ �/��~�#��-کg�׳.����|�8��IHpSBr���H�Y���_��tlPD�
��:9�����g�+��wg�iE�8dFn%�@`��eG@w�((��	k��!"-�S����7�2'���e�߭���Ԓ ���L%�BԌ��B�F'��o_��Y�4U
􃾾M�I���X)C��᰾8�3���̾��Vr[O` c4�8 ^�R���m���(zG��(;��`GK���5�D]	�0����h��k���zz��x�T� �=UDzz����!"cB	�Oӊί��.�B�-.���H��xi[�e8�!�'a��]T5�Z�����	��AP��7�*��7�CV�C1t�<%�,�@��3�<���ٶ�碪q
*l�i�/�%-q]�$���cѐ9(����%���O�Cyu,�5|v(��C�t2�$f��.p�oh����"Q�8r��J��j3����˯�4��F�O'�H
��P����38����I�
D�k\NQv���x[ �ѱ!�=9��=��4?�K�����;��R8�ބ�S�w.��M�ͤB�����0�J��:Ϻ]c�.�9J�����^�{��3��E��"��� Dɹ�n4($�r�Tma��u���V�y�<z�,]{uI��,�m9J￨B1�w���)F�vxt����n4����3��*�4X��t0������X�u+��};
��7`py�`�<G^��Oի��3�2C��"vf�au��	[F��ӋeX�}> ���y���sx�� |�L��gC+�Y4g�X.�g�ט�6D6	^��V���>;�P��WK^��,'W�q�1{�`����ЬNB`��K�zh8C���o�hl2 ��������)��C��q�[G�=Q�����C����}f��,@�r-�:������4z��:�/55�R=3C�&:F"�('N�2��>��c��t�7��t� ��$�RC����]����@�&%m[Oɾ"�/��#sJ5O[�_Z:���W��W�cy"��e��/��$)|垞WY]�8��e�u��m��B`4:LK�P��F
� +���C6��k��ٻ�|yÏ�f{aTw��+颅�|�Ze���}N=jw4'��<�!]�`D�:��ɸQ���$�W�k����:����঻���+H7&�(��� }r]M��dk�®a.��/)�}*�d'�f��5�������?KSx.ߙ����Xw=u5�0�����s�'�	Im8��t�E�i
�r[ozj���ܡ��:)�!*�t��5����/��qƹ�H������L�� .��)���v{��;�/�'"]�F��L���L}`�O?��ʣw	�4�x}��%� ���P]p��2�"��]�SG7~��ťt
yk@�wV����X��ap�5s��o
�vxӪ��(z�1;�7�Л⌷���FtRu\Sw�m�ۑ�B#A�_�\=�q���C�-��F���Ts��X�!�7��d04"ʁ�3-�ΖǩaՇ]4v�VK����q=����a�4�@���_��t��:��M_��a���x,��T@i u:�܂ʍ�Z>Z��(p�־�_4�v�9/��ˀfm�~r$�u�3P�8�����cיX�=;;-��˖6Ѿ(m�IރF	.t��������'o5c�hr��x�>ʲ��{��*�`"���N^��0K?e�p�i;��+?s��R� M��{�����Bt �m�"8J/D��%T� z�#7m��<O���7%@=�E�XF���s��+�O
Mbg�h�O��j��&H��TsVcU9�y$&mrQXm�:"b���]'hm��zlSQ���W�K�+A�'K�	m����v�����]�������z~Cy��ੌĽ~��'��C������������,�� --��h	�H{,L��|��K�)�l-,}�Nw��=���mgt����/�%�����4�=<����� �/1�~�=���4��."��C+�����; �"�n��ـu�"gdb,ゐh���pU���z��@�P�=f�M0+5����{�|f
��RR6�qp�X�MA��
v�@����:H���a���3g��i0.<�U���#���b����%��n�j`;.��9NK��kf�v*�?�|ȟ�;���;5aÈD��\�@��+�q �/i�5��@���'�/���[�z�huI��x�C���x��f��e�Q������ǭWw+�a.��"�����I7�����[�E�g�1��G�؏�h���J����d��EA2���+@�����<�s��lg6�g@\aU-�����VOf���ԕ�Y��q�-�rxU[D	Ϯ �8�o-��ꊏ����$����Զ|���^'�]0�/���qs�`���A��
��?�M�y'��3��)�M<N��ëո��8�m�I����K}�'�6�$�q�W��9 �8.�7�+Ȭ5�0�}���9����qNq������b�i�x���J�r]���/Ν�N�HT�����E�!��6�? �>����"xS�8q���ʓ��GB=1H[_g�#?����������;��JSǜ񿥀X���D�ߕƆ'���Zk�ؿN�G���]Fm������N�Y�X/� \��2VH�:�7=ń�rD9�u� �ERFw���U���yJw��D��@sB5��y��l�'��bka$ai`�ch�ƪ�e�֗��E7�� �b��48��c�+�Ō0hu�ĵ�6���@�ҷ�0�x�L��K!��%������|[���B�*]Nr�d0���_P��՘=����J�����1_m<������a�b� ;T�:���₶0�rw$�mX��y�:\�Gp�B5[�0��R�n*m�9䋜��<�Nd���)HU�7[߇]��i^�C��&֏��yѽ��P�~Mua�i��Z�Z�fFN�.�+��n��I�샗��ZO�˩B.�č����^v㶠i�/�V�s
��X��%����؇[,��@�a�K�,�]�Y9�_��'[��:D�]���>|כ�gE;Il~+&0�: k�i,�?�ȾO�a�t������X+M��W��U���{�3����z�����B���{@X0� ���D*�D*'ra�����ҙ��ĲK�<b�ș���Q�j`������\m4�^��~������16����=��B&�Mhq�#��%@�(����V��ܖ3���-�G�cyS��)[���ݛ�c���ۗQJ�����zi�c��kO��=�X�[�m��|/(���}U��=��3O���IK��|���/�\$v�sF�@�����YL�@�4�a�-�o���+F��2�׵�*EN�T��0���>����.�� pP�â��)���z�;7섟sJ\�5k�W��t����pz�Ñ���5��l�P_�C⽦�7eI#�/=3�nqC@������������ʋ������AY�j�mƌ��������c�iԬ�q�x ��{-"c���\g���3� f����}=	��nc��?m�V}�!�ᑨ���[�.�<�d��i�# Q@w������gb�\�[�op�����OE�y]�6$i�q�;���[��t�$x��+b��Y��ѽ �m�G�D�C�p��%��A�+T��֏����O"V�Fx%|�!kG}#�!�#dR�
�ܱ���1Q[�\�^fǪ��uM�?���T�H
G��?/#�v=��(E)��x��h��NqT�"����	�\=(e��2W��Y��u��V|O��9-�����GSk>^��+pRU�ȽS�
E�y�QJ�l��sf�)�g�z��W�O�J80��yM���_+7�m(������b�Ͳ�+� \�'�r*`�c��@0�����Ew߼�o����<�Ȧ�Y2���F��*"���p�,��j&0x�#�� ��-�*aІ�z���� �s�f�N��G/�wy$��q�'�(e��o����#z)��B�N5 �[��/�� AqS� -y�d�����K�����x�?t6'��złd�N��������V�Ji�مU��s�q�o�W���!b�b+W�ꬠ���O�pI8��.���lvR�-Ja3.R��`u@;(��FM���Z"�Y'���"�D���"����\cQh��="0��ö�f6��k���ʝu�84� �~�r������X}!7T9��ګn��g"���ˈ���\m(��+���i8��16�����Rު?���*ZQ�D�u�7�����x�ؤ�8o�C�,�g�"��?���r���ڣ��f�d*�u�8z	-����lc��~�xFz.A1�$�|��g����-�&'+@�Y�T�D[�
"fMk�)��n�x���{J�	+�j0O���>�k"`"r%w J*�`uC�Kbv��nS���Bw���Ż�~t����u�,�	�Լb�8�[��o�>[*�os���f�~�)��ku�߀8��\���֓�C��ݮ�H�.�aH/���R��M�����Y٠�9dL�7�%솗�����+ ��,v�&�s�*(q�Ð5�& w�6|v[h������;��W�|�G]�M٧ (����f+ �5��1�mA��IG��B
/�xR>��g�bt��5A��p��"tЂ�h��$��8�XUy��BgW�uh�p|.����,�[bq����4���S��W�on�0�t�j���!8�2P:S�sm"��HQ�0����Y�rӛ�9n����/��)kiA����C�J�����?��]tI2�$��m�Ja
c�����qE�N�F�NB����iu����)�Ӻd)��mR���`ɣ�r�^��.�����P>*׵?3���)�9�;iU�$SFK�̝ɧ���5�<��S9 ��82���R�'���&�{���7޼��(ޒ5G�y�~��ϑ&�o^�׍��u�w�Ӽ-�"(�S���*��c�� Q��rH�K����2��r�9B�;�\��y�Uޭ=��l�x�f+5�X6`���)�ItQ��%��{�O�t��0�Z�/��krB�7~�3�`�͟�h��2=�b������qʶ�P�wP!e� pA��q�� ��,'���w�#wl1U� N�&���V�~��kU��3�zM��ʐ*�-��Ro-��DΩ���+�uM�+�̆b �6�4���e.;ߌ�j(��B���T%'K�e��*��'<_�.�VK � �6��N��KG��&�n���	^���G��M������]�Y�~Z�,ˣDn@Մ�3( 
�
���X?��*��zX�7�I�%C���:�,��_��zWr�0<Dt�i���g
�
2��7iE��g`(�N����3]$�67e�%3)<Cx�B�)nqk�\���ۜJ-؅d�?��*H6�*m����o=�Z����,F����N�l3=�S1	��b���&S�/(���o8�@b~U������O�� ;#�xG#�A�$g����o���]��Zz[(�m���g߁�0-rO�)�`O�s�y.4�Wts��n����O6���B�А�Y��x`aJ?A�:e���F�>�K�,g�F ��3ڇ��x��9��/y���zl��W�`�:���U}��%�h�Q?�� �d}�
�y���K��d�@�a"���Ψ[�'XN��.r{���KL%?�-C�`����R}/]��G;��i�i�CҺz�
��T�hk���0����t<�����z�5;J�7�RG� ����z8 5؋�	ʞe�E#���W����Ʌx�X����H��
lt��V.O�P��;r��Q�!�3 n�&J���a]�=v�Kq��mJ��yf��P+���Hgη�e^n�[����$jtm�c>���ς�XpC}R�=�0����;0L�5a��v�� �L-W�]ʎl7����NB��|�=d����2�~B3珅��^k�O�p�i��@�
<>L��dt�~*ò'@Q���V��÷L�D���<t�
�
Wש�ݯFFg����\��ȗTϙ�tu��3��l(f_����&�@���]F���9M��h�g���\�O�[�9g��>X�oOTȓ�FDp�1��3D�f�؟���ު�a�Q�a&r<�A��2�+LX>i��8���+�B��w���2�;C�)2F�2U<���ڣ����Jc�nUl�vj��(��I���&U
ן'90�:~ѥ+�y@F�ѝ�+��L��mH^��-�L4�}�ejEB�U�<�e5�ɽ�ܧK#���г;*��#H��W>��a���tM�$B)e�
��NQčn�Ӊs
�Q��R�D5H�VG^}۹h�hT�V	�U�6�ӒT(���	q9-ai4��/��r���\p�ٴ_,E��_)
K"�������ޝ����V�+f�T�r�F���m�6'�W��=K�D�YE��d�j@ D�{h���Em����Vl[Ol@����	c���R��	��h�M[�ư�
Z��� 