��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd0�0m���x,� �m�ѽuw�y�,`庎��|#�)��]cBt�z�'�f�Z��!�k��\O:���F��\OB�(i��-�"�jGJ�[#5aD)��KX�S��ǻ�)��~0f +�Y�3�yJ��&
���X\U�]�����*���&��8��b\I$pb��H�!��I���������,lgK����Sѡ��N����°�0�Q�`ؖ/8�(X1������ަ�4�
� ��]�W�oP�����ńʆ4�B�����ج��Q���;C�$�	�0'.��Hv[��>"�3Ȼ������¬Ʋ�����?��;A�w)aѐ?��Zx��Fή���^p+��	��K��]��s�dՋ_?��&EBF����Z�o=���8so��1Db�3Dem�i(���0����"
���!n��PO�
�� fB���IQ�ƪ��ͳ��Z�J���4M(M���|�6r��Mx��3�ɍy�m��g�.�]<�<X�tڃd/;�SJn��qS��#�Y�d����g��z
�OR��i��M�#� ��r|L���O��+@VK��y���^Y13�ӭ�7ۛa��b<ݬ�^p�8�{��� !�/綁hZ�Ǘ�揔��%���m`',ۑ�%2�چ|x���Q0�AWz�@�ƀ;hv�nI��:x"�9���-� tx��� �r��xZ�:r"�p"o-Y���-���CR��JҨ�e���m�5	��5w:��۱�x);�������Ո<��3*��u������G���gx��`��ۤ[,�+.O���H�DE�e���Re#6���T6"���mwX�XV��&`�4 ���2j���Z</�(�"˚���i1�ia��}�_4X]Z���Pˋz�\���wɐ
�,
����{�	d5��`|F�5��Q�������v�J���(� oU���J�]�\�AnM�e\��)�����z3�K�h=�?Z1l�P�����.�Hq��MX�V�T��1����Y�fe=���GH�2�ٮ�(��`yt�e
#�x򫭙������>D��P{m���H"bsݲi�溅 <$��;�.��O�G=GD/�s��q?̻[0���2y������tz�?֌qf���&~���9G�#u�vE�*ǆYv�}�j�.�9U�Tq�b AI*9�$�d�R�
1�=�,ᩜCF�Ҿ���x�����":y�e`�K��j-.�*E��[�r��R��Q�k�Ӵ���iw�G��T�c�6���[X\uJP�E�(J|����mV���~l�6�vr��P6<��Ү��x��g�u�����EC�aO!�i8h	T,-��\%8/=� C�d�[Bp.שi�	$���FR���j(.�	U^o���τ �U�����˞[��(/:Z�߹F�G��T(uw}j,�( 
�������D��ZN�)��L�?Ϲr3t��ǫL:���i��0*��~�m0�q�_�ΒFy;K�[٠:����)�a?RV'��馾5+����8����F��t:��_c6�Ĉ"MF����̹u!yϠ�3��c��{ca��ڹ�c��A�^JZ�5F$�&�w�B�?`bH���u�δ���lz�O;���� iL�x?|�ެt��\V�������>�P��o9�E�aw	{/
������By�qÐ�e�>�3��0�qom��ܫ��9N�� c�S!+Xc�<�^��#h���z/����Y4�������"i�k�A~z�b�-��|rL"��5;Q(�;�/��񍍦O�M����*V���;3��e�W�]6�ٔC��	�Bd!�d�.ᮝ7��㗉 ;�c&�$�����穝��?��>f�O��g�3�L��z8 �d�`+� �J�,<V�D��A8��<�!䨗��n{��r346��\�HL| Aoa��F�7�4��k�p�J1)�T)���5����ѫ	$W���_�=�G������,v�"<X�j��m�����.��=��J�Ξ�]U7]� ��	ษUI�d>]���Lma�g�Ky]^�����Q^�?�\C����<7$���_8��/���AU�����i5e�&�o�}E��-��������#o��������3��FO��R��ꋛ�p �T�H��<�ϔ|���M+t�3�	��33�v�>\<�Nx�m��G��bX���kI�����U�vg/���І-h�]���ϺVTk���k�co� X/r�������+�gXyG���7X�7����7[Je���P�������7KQ�m�q���^;����U��Iֺb�ܨ��&;�*-����k�oͻ�Nz~Ts	X�q���t�� ��,�H�j���M�a'�Ȇ��[�	��U@�|������@���ʹho/:F���&U��۩����{�T4�����[
����ap�dB�.�"���r�1��P�bC�ޏ@����~<�[T;N��%�B��ī�~�%=�D'���uS �9���T!~���4����s��G@��{�2���w���u|˪�0�s+/�ө6��F������
h��Vg�^6�/�95�i���G3.F���R�3�	�ǽ� ���^A����ے\5��2d����J0��(L]M���c�b�?�KG3��(�P+d��d#ax����`6��F.�Yԋ�z��u}%�|s��02D�2���bϬ�k���!vv��d8#��v<�_��Tw���Ϧܟ��8b"�����-ؑ�J:�NL8�uk؉Oaa|8�*�[p,TUs,�ci��I:*N�&_��4��TC��%9���v�8Kacv�~Nry�Ò���Ym;��܅��hKdU�Zm�8�$+΀��6�>�F���i(Ļ�B�}�h��[�	���Eg��|���~��x��_GJ�=B����!x�m[R���i���S���R�?����?��V Bfr���p�qGjP�ۊ	2gIn�>�@a �����Y��w��f �y���/��l��Z5,�Y҂� S}2.�#�VNb��Sڪ��T�w��wl95[���%�p��n��࿵�{E1�r��l;� ���m�5C�
8�������������-���g��wқ�%T3��@j����:9YB���C�~.h�C���fd�s|=$�0�f�{��{$7`��!C�] �rIO�fp�go��K:��u��h\�lT���ZOF�19^ �E���n���O�n�_3°~Դ�p5��gaf�"dW!=���F|�*��~59�"�=����K��
�����'�ҿ�\�2d��-����9�Cw;�.v�t�����-s(�g���ԣ��t������_L	!	@��G�2��t��8����
\���M/]ף��{��C��Ƥ��0X}!9tQ}6pF��Y��AP�����l��Ԩ��D^
��Zq��=���k�3������c<��nz5%}���#&�����B�*sѾ����ՠ��4�,]z2��?w�[�n���{��-�1�!��C~�5p�o�Ʉ_T�"e���Ů���Q-h�>�bd�s��h�M��D70�8�bR�Ɗ)���g�&8Hy�Ď�d��fc�.��`�*�'Oi����V2���:����E���{h"�����<dt϶+����0<[�)� j�VF��[���Wu�#7*ȅ��TT�f��S2����bL��5��T~Kܙ��p��:���b�n���I�h��Y�~v4I�I%K��`���$�ޜ
%5��_$0�B<(W�p�~��3�\�^���eR��zE��i�a���,)�[8ޖ���Kz∃���΀�V��sRb$C�a8�/9�fP��n�_�bv��f���O!+0�Q"��C	c��Xu��H�A>��?�R���Ah��YUTG���
�ڃ3dk5/2K��!���O�Jx6����W_�r��jAT���p<���V��(i���NC�7�f�')~U���FŇ����$���;��5�rf����r$~�0qVj���%�/$�ɮ���@�"����ۺS$���A*��(�b��7�c�����z�5�;�M�M�=XLS����鄊A�(te����n�i�xŚ�E�I�%���@����O> �
�x�3s�.Vc*_:�Pt��&Q�3�l��tr��7[
�Tw�=f:����V&U~��N��*)򍑣g:��ʃ�Z�微�s�ވ�1�7[�B��0Ѿ��Ui~�萭��l�־���$T���B�򡳂��):�O�\U:�VA�t�%5bI	2�L^]�D��r�#��X�U��Il�G�|�!�N�f7�z,3=�8����#�̺�.��DZ��!���K�x�#{c:o[|jx1�Ō�i�k�I���g9�ۢ�Q
���� �Gb;.8_$)�������	T�z�8T����w�OwV�O�W5��v������b�L|��񶃖!����Ͼ��Q�ѩ��-K�aMv�������zCQ����ΰg8�`��LAH��8�Bh�[ZUY^=��D����Z:*�%��z;�F��O���	L���F7uXa��,�?+^����*5�8J[zH�2k����NJ��s=�Ԇ�b�" ]���)�҄�4�=�n��MF�	���<�@P�ͭ��������rP��d�LH���㕬���ՕbT9�9��0aV;��y\�K\��#�뼜s����/J� ��Lg�X|��E�z��������lۋ��"/Hr'�R��q�/����E�&~���ʛTw}'�eMw%�>����*TL�Y���v�@��)baL�kl�BW ���#�i�̬۞5�4���QE��*�b䰥^Ҩa��7��+2�h#ax%�j+5��TS]Q�A�	&��+���lRZ9�fc����2�~8�)~��Y$$�����c݁>�����L�J ���IW�>������{�]st� -_Q��*��w��L���ŚD�u�E����8�)�j���.t,sމ�@�W΀
��uP� ~���Z���q�Э��Z�?�ڝ"�W?cl}�D�5�������Z��vѠ򫦉���j���q�R�C���>\�M�<*����a:��ZEM�1o���qeVH�Z�2�Y��}�3��b��;���Ol��5�d���z�ֺ_xE;�Ua�]�#��Q�\���%+Bǣs@YW�R����5chM�L[���� k@�<��]�q�S��˓��������t��1�11����ΰ/�Q�>HDq���IC9&�ssծ��6{�?4ǿ�����ϸW�ea�&���\���Ƞ�S���v���X��! �7�e��D`���Yqp�Ocz�m�&Ōǂ��xT��/k�� NM�7�	J��"�MF�,-n�4\�?cp���mZѓ���F����hʼ�x*��:������qJF� kAf��>+�A��8[rP�w�QRD��ݐ>�s#�}��q}<�iz籛Xm/�K�u>Y�a��~�6�X���20K6f��mqu�(��դ[1���6�"[��x���O82�΅�H���vUk�m�~s��$!c�^W�&��W��t}'�Y��P�ȜV�B5���7vW��8
Y<�
��FG��]�gyв�M�Hr�����1 ��G�?�]d$�\A�%j߭��TM�6X�N���W���P��!/w�Hk�Q\x�!Qs8�mG��~ơoaA'-!�zM0�ϜIb_���ֹs�u2l���&1%�d-c��#�k#�/H�s]�r������܍T2��h��J��� 
AC���m�P�¼�P2��0�_>w����x��W.:U!t'�5.=��&���:��҅�4ҿɕ�ܨ�Lq�e����P�iR��(�+�j���W��~U�� +��9O�?6�6�:������.���^�r�v�E=�ٔ"�h�Xw�y2:����(��/LJ�C� �Kc�:��/u���5MI���OB�S#:G���[Y~o�=2�M���j/�/Hѹ�ɻ�k��"�j"破��%�a[<-ۙ�@m��>�]�4����N���Cr����Kz��_j�q��H�=��@n�"���b���O��ވf�I(��gcMT��6����r���5��GXŐ�HCt��$�zH�Q)oVLz]�&cZn�p�y|�g��bp�(�_�Q�`[�	W>_���<���cX���znMpԉ�iLЖ��Lj�
�@3���_���{��"qTw!E	�#+�a��(Od?�r�`?u�����|XN#�N�M��^��|�̵�u�Y��5��kcy�AZ�6�X��083sƘ�H<;=#�(?�:;jz��w�e���$���Z.�����
U�r�2+��k���k��Mba�cgn�HV�L#>h&a�8�4@��[��fzk�\���"[Y�uUJ�v�h�QD��<X2�Gf�U���*Zʱ�����q~p������ҁ���78�IZ2=�fy��-�V�B�U�f��(, 7�]'��Ak!�VH��ݩ�ċ���C=�c,N�]��*�?]ǝ�$<{������e<��˱"T-��-I,�E~uZP�:�h��r,�Og�6�Tz��N� ,�d� ՟.!y��4<��^8/�j��V��� &���S
��!lRC��Y'j�*��_I�\�ˤ�hY�p�z�d)^c��ګ�җ��'�ui�n>�Q%�(9�5�2'$�ҷ����,��4@���>*:%�2,w���j��t�����r���lY��$�5-�=�`��ݥ��~+���Mi�+��研�*�Y�2lQ���Iڊ����JC�V��[sΈ�ϓp��%U��;I3����To���4ġgu��q:[�x�a���¤<�>Dr ��NĒ��j��S&w�O=BC���B�W
Y<%]%���m�w�;~��bg��ź���{@�yg��-Y� ����0�}�Ml�)��#�����1��1Y��vJ�wA
��q-���S%�����Z���=/�=q�l�P@��l)w£�B���	I��HO.Ef�tU�7g�!�h'G%hXq�*#g���L���FH���P��y�+�<6��L}C�d
ɵ��PEcRj�P��D����jj�:;ą���5�'2\��0�K�1���G��C�/��T�їI�= �SY&���(�$h�@Iť����I���:!"1�J*I,a��!}�n�	\�W1Raь]IV~��� �k&�=�y�b�,���.�8� ��/f%M�$ffL���f��Aw>qղ8λ3A����=Ʈ���E�?ň`-v�Ȕ��Q�P��h�c�s�v��fhl9��lw2m$|��;(=a�������,�f�&��C��U�'I�uOf�����ƃ�T�⭎�,J��':�5��Pp�:��7���ߩ���E���4�=����$gv�Mq��ZB�{K���H��7���������g�#�T�iw �*�7�'w�W	y_Bm��5�Oޣ[�*��pb[���c��+u��I͸�5�Y�RPK����������,��y�5��;��Ew��V�[0�_9��]��rj�8�i�R����^�b�&M%J�k�t!�|+j�apі�$q!��X�Q��LR���OR�Y����0��(��Z:��]Ti��-�<le%$�W��B]*fI�-���P����I�`�p����7�E�@��%|v37T�!�FE&�̠d|�7w�t�!R��㽿^n�p^�9}��fvg]jO�)4:�d��]�����w��	э�&@l��aV���ܿ�����1j�E
�2(�&�a!�4����
�z��5��{��o�L���L��i����#T
���{���6Pl��_�+�1�}�:����L� t%�?�P� X#zv�@N�iК��e� bzi��rR��1v+C�%���h!׶����ZM��/S3�����Q�lt,��u����"��!�K~�����d;|d�%��(�KrD�\��_�˭���=sR��(Hjξ���$i�i�f93K�������!O�
)����%iT�L�V_��*B��^�?1�?Jx����tP:�c�����+ ȴ��.i�i�3�����_!�~:���,�D��{�BJ,���w���'l�������򹭋�!Iɪ�aW�g)PFT��=Ip.$�))
�e�f��S4K#��x�]/;e;���@U{�$])��<�*�lW��}a�\���,5�|����W����5N��#�݇�W��J�h�S�:P�h�5#�K	�c�tJ����I$�KGr?��|C"嫤�jV��Kf��� -���g�v�k�	��|�.�����5�O7��[0Ez�H{��a/�5��E���S�k*�R�͹[�R~��J�k��j�i<��$��e��~��g���m&�B���ߒ��~�� oK��0�{����8In����{�6%��3-�1f���%'	��<1)Ft�	#Ug3�ꗒ^�:�w?.��Չ�T�	�#�V��O�|�!��[� �>��>�AلM)���H������c`�۪h%�\�!� �[3v�ď�L(������U�aec�ٙ��U�m�J�9S_V�L
������(��[�]rհ%D�,a�<$q��=����u���Jb)f|�]��j�c�]�t�#�q��Pv?!r���<�C���Xٺb�f���� >���An�`�M�b�Q&WK�FC%Rh���vr�Gz��ŵ��㨒����B��T_���(}��;� ��+RַG��po�d�z4�a����쭇Q�`!D[J�r̓}Y�v%]��`��4D�L`��k=�RѮA�(���܆��7������m�o6��w�>ե��|�X"�|����/�ν����*ǚ�%�H��ü��E�o���Xn��J2H1V�q_��|)��';�'L�>�T�G�#+F�����U�`U=`kJV�(P����{��B������P4�$��z:2z��<���I
bC�i�4�1[���1
*W]�7x[4$ �4���c�[�˃�/�~]eN�YO�2�v؎�i�5�H$q<s�O��uy^42�p�*�O恐g�½�m׀���Z�22q4Y�A��@#�J^�^a�/Y�";�<������#��y#'�B�-������	�٫i87yįDx�X��QC襪e`��p�Rd�������ˬ���K�_�}9 ]O)�Fy��K���n�%}��`��D�B$���U�Vw�I��_�w5�|���Ķ�Tl�&I���)�b�.U�a=�mV}�(�U�E��B�7����"�;5�J`��ז�&��cGى������O���4�Lr#��
78�r�1l�J�k�;�x5!��U�����@-�k	5���/д}s�r�:a�k7����b5ϙA�U���R���K�6�W�ppmBP�nK@�;�����ݪ�`ι��u�&P�������_�C*�@�1q��_o�G��[��ӑ��,��\�xe'	��[!0SO47"a�`����1f`	ªg��ߝG����������w�&,EOF+���#&��EB5�D�܇m��H4~T17�득�*E��;aT|��c��ҒG��sޞ�5�J%�.܈߁����-7���#۶��f��"�ra�Wh��od�׿|HŰk�x�d �A�UȻ�'�ڂw�޿�?�͘Q$� �W��(Ӂ2��	�w�e�'H.߿�MS9S���µ��P'
F��O0ss�gKlL�NB� ~nd��0��kQWzM��HC�fC�T�Z7����?�5���GQ>�)��j��lȘ��x�MS1-u/�LXٮCk�_�Z�@�m��D}��J��۝�ʡ��I�E�<�7�A2���j�����X����ȏ���Kxjl�n�(�L<��p��!��S,s���u�*̿��� ��
������!�8�	8�;l���	�_��?t�,�Ab�,a@�O~�fA�؋Q^�:w�ܛ7߽<	�T��>�Y������<"���s>Z�7d��������
�|`��KU��&��5����}�3��t�T��f',�3���b��y��i7{qB��@��`n���>�o�ƈg�f\�� ��<���0�x��>MX�2��m��Br������Ԏ`Z��[��a������}�#𒟻��1d��)o>)=�{w�guh^������ǖ�������m�{P�Տ��25�/�*9��@sC�j��{T�K�Y<$�)|�a7*9ˀ�������}�_x��6�+ţ�<�,�u�GŖrj�۴��k ����0H��9̭�zQ��%�����M�`�����(9*Δ�V��p�,B޹;�_�a��8��!h��qȧ��@xg�7	��7Y��B�:K�]�I�0O�����޹g����C�P���Ù1$_��]�)^�	���z���w(��CSn��
����n�6����{���֛>J~&YB ��L�6��bL�k�Y�;�_����b������[[���*h�ݓ���_� ��c{ʼ5B��@��{į3�h	W�bm�$jG�gX5@^u�tLS���)��?R/�Z��*.t~X|p���H�CԜܩîc`=�,���(�A4^ KR/��ɫ�gL�1|cq> ���hb6�(Ө��л?}nj���i�_u����kDQ�҃eq�O7��Ty���F�a���%�&�ˇ�U�/!�p��^���夙�{iЅ ���Ϟ��`�z�
�?R�(�����X܈^�.���
��φ�,%X�;9<� S�q�nR�Ĵ��{��:f�h� �9�d_02�\���}��5��NE�[��D�|��r�}�{�N��6���+iPMĕ�Op�專a��<C�}�ù��2�N�����G�N"�ԀI,ߵr���T�B@�̃���U(,}^msA���Y���;^�t���x�m(�D�G��T�嗘��њ��q��֎�캌<���C�4���=!��F��n�ikݴw2[�36���J��;����x�;��!3���m�݂�lρ��NoL�>�u����Q���`�����K�����!V���RGz��7�n����-����������MR �ء�fw�i������P<�T�ʯ���a��V���7���)��F� ,����{K
�ιش��<��td��a�M1ǫ/�-b�sy��f~�︹/JO�/n{H�D!��<{������yQ�J��?���D��lG{���U�� 'rtO���wK�@��'Z����.� N�V���t:�Z@ǽO���'^M�)W9�G��#��!�ص��^[c9�d����]��eG�Н���J�����I�^|w����&G��ژs;�:�S!D(�#p���*�*��rč>U^1������ǗZ ���b��1����
�	l.F���z{���n�q���Ne-�VK^I�m�@���p���F'� )PC�h^n��cc��{��`����j����,Z��PB�,0%���W��U���x�˲ře�H�D�Sŷ�T�k2Ղ�A��C9ʖ��U��d]�iI<PT疢+��h���%��oI��J����wm�;$9�ľL-�%</����A�l4�,4�/ur��
7�r	�,��p"�8�H����S��17�ِ�֘���e �Be�#�荱d� "�Bz��.��m�
�����%����_��V A�r��V��˽1��'LRU'X�b�휵�����<��R�?ў�� E���r��N};���~��"�;&�}Ո9����33��Q��И`�F�+�m�(+�8����D����fM��� d�~�Vp�z�5Q�;]do�q���jNv3b8`.�W����ɽv3_�����[
@����S*m�ڎ��4W�\�}v�f(�[\B�<����͞���#�'#9��7�!��~�wF\]/�f���ԭSI�|��b�:��{G`�ͺ���I�/�����-m�{sg��B>�U\�[S���o��uK��@�H�(�㯘)����*���6��S6�j59G�~H���Pw6�ȼ��B<OV�'�r_�_Qz$�y��j���c4�!���=��U�g^�|�S<�/�9��ϩ��� �B�)�c��<�?��р�m��7��gG~�P��<	߁�-�H�Ԣ
[�EK�/<��w9��N��ቜDֽ�!:��[��:|ܦ�߈ �U�k�rA��*4!={x�ʙ�d��ڙ����O�a*�-?�R֧$��1&�d�E��А�����ts���?���8�|J�OF��<	�sh�n>�eZ�>�1�;5�&�Q`�%�库��i9W����������o~
�J�������<i�xA|g�v,7�9˃�:)pL�~X4eĽI�KG8)�����ӝ^|�ﰹ�@�]w��Kjq�G���{���C�(Z[I���i3��i�Q�����5,h���I���Y�!� �2ۚ;K�S�h�'�ϊ97�� m��V�*ܧl���A�� �ѹ�헻p�%m��h��Y'P�)�+n�L9\֨�\ϒM��J�9�m2�p%y��(~}?AlQ͐t�3��#z��@��)���+�Ap�1��3dt!g�Q&�I��og�ÿ4�I���ӳEQ��V���ˇs����@��6��S�]hr	����
C������)V�Y0��@w�O�`���!5�K[t��+����0��,�� L	���u	/�r����v�IӨv�)��ى̋ԅ�<�ĭ����έXZa�IP#�[R9�t�K E"hd�5X	����:��#p��� ���C(��N%�[eM�uƯ�>
	�������t0�T���` Yn3�'}�e� �������� �jBT�Ӕ�I'��*���cR��c�����LU�5$���8ҩa��'��*$�RB&�J����e���g=�K�|��[0�~�є=���vTJy�x�����	tĭ����EE�V"�_��s-B�",����B"V�\�g4.C韆9>��iHF��\�A����1��Q6s"Vlm;hxCD��Эf�QT�GP��X�����Eh���y��^�n}�9�7I�A�j�:Q,ӧ��5�1���o�5f�u�P8���5���Ux��؀�6���ÉRF���:��5%,��]>�� ��Y�ue��Sei��������i �N�6�+7G��Ɔ�j��
C�Ǵ��N��Ĵ8�d5A0�f�w��SE��H�ؒ�
������˺|�������?#��_�F���t��]�{��2�� m(Wr;��	�0��� C�r�>XATSw�zV�^9o~v��í\%�I�T:��7�z�7^�s���e�C�r8Wz��z���W�&���?El�^�9�{ֱ~kK	ǧ���**ot"��	:\�|�P�,6��N�Q��y S"4���r7���68�L;�5x^j�z�@h�)�� ��JOj}KV4��%����e� �hd�n�l�բk��S�$G_²��I���ΈR��Y�!���kR=R��d��M�ڍZ�&m�^#P_ۅ���hP5^q�7`���N�S�c�����ͦi�@Ԗ����{��5g��/l����4�lA~)ݰX@�w�T���S ��a�-���L���3�@�9&q�;;��܅�g�O�*x@���(Ӊט��>\��U1��ә�ր�Qb٪���CJ�JH�0�hE�7�W֛����F�KՀh��+�O�BPB�R�+
D�EG�Vç�dހZ�5�J�W�gE�V�%��uOWC�m�I���"o��W���]�7���"m�y5�����c[�d�]������~�� O@���-�ΐ���YsA�L�w�����g����(�@y<�p:�Ԏ+��bͥq��mb�,��`F ��{j�&�em���w�]��=�O�<d�
����V�Z:�N�W��jӏ����	r���V��` �+��S�z���W��cId)c�_y���:�16p<@���3M��is7J���\�U&<���|�e�\?���V��%$�z��^��ڡ�y4Z9�����h3r��KXlc2�"��w%��(��	ة,j���.�S;��09q~,|���|T��z��q0ܻ�x�ҥ��(�i�o�HH�c8{���p{!�"�Eb��E!�1x�-�V��b��ꡔ�v�=(��g�֦ï�|l�U����}���M��7�ǥ�3���N&�b��R���?�c�L�\*��g�l���	O(Rɜ6�J�тVmcݨ��ia2������4� �Iug�`߿k���,9�ͅ�c9�}�<���FX�7���9v��4=��+����M��������H�8�D��e���l�}�����2V�!X99_;�5���N��9#x�+m��m�6@UR'����)��z|���B�7�#����e��H������I�\�#�Ԅ�$NhEm2�e2[>;����9�d�>�|%���j/1U98��\�� ��Io�ag�a��ѥ��UV��E	+1@=���O:kՇ�$d�w�џ1C^���˱D�o�~̝|�%`P�hm'4ע����Zo�I��F�dݫ��(���wr��GqFJ��vʆ�Z/�8��m��B��ʘw���rDÞǳe}S���c��{�X�oF�rj�~����T��i���p�Pͭ�_�p��kҗ�Ϗ�^C��#^��Q�}�;Yb�eF7d�+y�Gg��F
E^I��-y��B�S��6ZE����>�y2~�`�f��ϧ��˳���O�H�V <;�;I����0����[����X9��t�����Ȑ��JoL,8Ƴ�Ffw�i{�,f����cSk�18ͨ�R��:�$��r���מ-�cs��Pzoe��8~>R�t<3�gM�u��0�fOL�p!�"5�a���#�(2yO�4an��T��Bz�Ǜ!��|�{H�5U�c���ln�16ݐ���Q��7�$�B����1`R� ��D�ȼn�Hf��ry���"��mb$/qP�������,�]T���r�&�|1ita���v�7��N�K  �q#��6	<0�o�4���4�QN�t$��xXY+�}L#]	�7���$�t<;�5�@�p�K���c��Vu��3
��)��a�� ��{��M����t���gĳ7.�U���]YE� ����er�����b��d���dox���t(t������=��7�U%�.�|@.��c�O�1�|�����U�hX���e��Ș�m��F)V،�Z5}ߜ/����1�54��	%�r�#7O��(ꊵ��"e�}���rQ�w��7�w��PP`ELˈi�9P��§�7e���Axߗf�>]1Ҍt~,u�1�FB�ߺ��SU1~¹��LBz��K\�[����3Lz���k,Q�Q.|�c�a�[�k��ݿ���d�ߍ�0|��(���#�����[�G�sƓvy[�v8w��	~�`q(VP���2��+�r�@AYԮ9�CQ�ǀ�v���'�Z*C�瑩dK�C
	�|g��Ʃy�=M�'��X���ʨ R��D������6%��U9��5��0��V�Uԧ(��>	`���������q!���6(S�?���uy�x=�o$e���Ó�1�_�Wy8�yA�b����Ȅ�l�L�o3,��mou�Lb�c��e!x��k
Q��r�[��=P�dh�<7�e�:��!K^�bcp�ϧ�qXû���Z�}M�~1�7� n��8<g�qB>`�x�W lQ][��3X���G ��x#/һ���v
�s�f�l;}�k	�;.OLѴlۇ떫yfZ�;�W�.بq�`Ne�鯮����䉿�ƪ���~�W�l4j��6��k��v�(rpUb����)�͌Z`� 1�&9�|�?��D��k��3
ɕ�W��B���y�M|�8{3����zU�_�x@b����
_��]�~�4L����ݤ��O�+�#4�������yK���/���V̈́_�cE/���<`'�Ir�RyYw�����Z��l�Q&4f�sG������>(n�-p����#)��.�W3tt�E���ﳀI	�/�qX�n��^'��*�L��)8�M�(@	,��wb�У�}��&B���\C�JO�qW"T����3$^�shL�TsM�.ƕ��� O��*���d�Iǥ.���g�F��ٮ�é�o)#9�KFjK]:V�5�������%|���~ ||����$�4q��W(\�mA�Rjg0GK>b�����4��ZOnj��$������9���t�R��.�q�P���4<sb'#H���=@f��)B��b���Q�u��^�
#��O�=�z�d�n�e�(WNP2g��ۨ�a�\�zA*���C�Q 3G���H�4����q�6�˟ ���:��$�W�፧(�&].�V�u^��>c���v��Rxx�᯦�I�5�F��I�
�	�O�iuצ�i�f]7o؇V7�X\;��HcInՋ����t"��Og_��f35��ʈ$r%���}Xx,��M�(Z�z�Y|��7���M:���[�ц���4�������ob��^s1�=]n�W�q�jG�j"��E� 1lj���x���s�8�t��APyW-?���Bo�C�g� ����]�Iuk���ǑĂ;2)Y sp:8�l�'ؼ�c[�_p�d�hX����X��H)CL�N?�1/��_�E�춷�ӿ�oi�׫��5� �#�zG�r�!z��k<���0�F���s�Ucaź`�4����y�9��0�/+.2�q.�������^C�<9��{jj�j�Vi/�4�w-Rl�\��ҵsX�1E:�cN��si��s��=Ʊe����7
��/s~T5�&Re����?���B�?��@
�b4��ƙ��$h�ZD�!�|E�����I�q>�]�����9�߃` �`r}����� �j�wg����P2,ُ�g�V}m_���۟ Q����P��dj͘���oL��As`��}e�V���dgŋw%��z��WL�r٨� �.�`\ٳ���r��c�SR�m���%�c���dx:��;����\%��*�+<���Uƪ��ђ8)<P��>��;��.7!q�����n/�Q�U�O�E�Ա�9�Y���%��m	�fI-��'�e�Iw��ˏ׹f�}�I���IamMo�z��hq�sI�Q�������o�Z��Ձ�T������<d���]����H��S��-ڢRv8|x'bp@:R:�4]i:����kS��~y�5 7�5#Aϥ��2�<#�����_���� �Y��t*/��1��v1p8Zo�>rcf�u��/���2�K�a���y�L�t�}��fD�7�L'��|&�\���4�W9�9�U�-�=��I�0�wٸ��ǆ�I��4�*P�T�D�1A�BCOe�G�!�O��_j�tӱ����%��F�	:��7�6?�J��F�j[�Ze���!܍n�r�Oǹ/
�����^#�N&�\���zO	&��iD2�u:%«ҽ���}Z�f>�L�x��me}����0٪		:�:$�f5nI �r\�V�dG��?J�{����7��0��B�k���`δmc��y�W K�U=�����1i옳�
G��pӛ���t&�Pq�v� ��"4�oZѹ� 8����?>��&k��;�G�TH�h�q��W��sW����]�	�3#�$���!��Up�d��6d���>�ۚ���`�^}���s�ѹ��W�+6��V'��[���F�!�L[������ڗՓ�:[˔\B�C����C��7{��S����-�CV�͍��U~�k�z�)��y���Z����rh.�M�W|[�D����?��x�\H���,}o��7"p+X���39"�&Xt����v&���x4�"h��;'�c� }t�%QET��_:��6�A�xd��j������1:s��3�L���ր��8�x��Uy��d"��P�2�F�-���
.0������E�+�.*��mY�{p�V�*������@�;L7�����kīz�/$���o�4�u�ߊ"����g���Y��aX)C��j��Riځ����h:M_;d�LSz��Z�~��]�?���J���מ#�I�S:�yg#������W:��Q^s�L6I�ƭ��ڴ�a�{,�'�����H�3�;�	�XGe/ݎ�B�hv�b��#�M]^�S�Q��(I#g���ρ��(�wE��|�,�!f�4�)���,;�����9�l@�G]��l��Y����.B�`���ō��j��P�tY��5P�lķVp�X����n.#�}�7M&5!|g��k&������P������ 5G��8ZaG��au�ǎK��������Z>�X��������H�?Si6������G�'�E��ZS���r�D̮S��3C��Fll[�[�Oº���w�VD�LҒ��l��t�y̡�X"r�Ӻѝ� �Z!��i��·Ba�bQ}�w��!��O+�|����Q7�{jz��جKôy�N8'����IK`Ս��v��Yi��E��u=����{���|�<�Xt���q���!|
޻
��u*��(���c�n��(���R���g��L# �շ��F�\�?�눐��X��J�^�=���]�*�E��~ǻ];����,m]1+
�=�*�]�Z���1a�V����D�+�����R�$�;A=ROo]��$x�R���s��Z�U���e�M������+�T�/��1u��=(�%3g������(j�$��ؘ��%�˱�۶1�����Jʃ�41g�5�^��6��:4$.�,笏}��\�Ho��"b,oi�ͣ�����\lEh����,�:<��(&�Z�Wo�z�����ۥ��l�)��� ��@}�m���SvW�*%�ꂟ�P�C5C�%�F f�s��9�����ɋ�[jb����#�Q8���؊Fc�n�0~Q��}�*(j�P�
H�N��8�Yj7$�#���� }B�y%�?�{O�čS��A��N�S�:i���i<�|��h�V?A�A��D�=�TdEЊoIR�B�o����3r�ײ6�7��>�>N�@��ݴ.$�%0 ��v�?�}�� |`�,P��B��l"�d��_M�T��,Y��t5�I��r���gL<-ZIȆ�;�����+�$��h�햿t��B�W��zs��E��^��M�P�/P�|^p
.<���Od������S2,a����*q�F�����#fU����эp��+<�����-�j���(&(㸩������}���b���{�&�n������y����=33�Iu�JEđǒZ�����Z�U$9�&�}4p_3<�|/�>��{��]�v�X�����||>$0n1�!�7��jWcF]��Հm��Ab��f���ǞR�n�����h���A�-���=�]}���I'�k��'ѬC�Wu��ov�at�gT�eU��y�X�`q""<�K�6D`.�*����9����+$��CC�X����CW׈�(?�>��[3h��{3�� �����D?|�@���2^ppBU!;�
8ъTN7���v��qY��wwR��?��l	OH�U?#���`*RR���	�S��e(`ό4�U��e�`��%']P��1�E��z�"�N��;��5ґv���|���ˁ��>t=��V���C�q�1+e��X���/$�&��Fc#:��|���99���A�
���,ǃ�� ~�U�\�'0)D�����v��0ʳBjH�V� �{7�r�V㓀�w�ā��i._,?Y�x�|=���,!�T�OY���X�3�M�iҎ���cb��z?��w���{]���~ɰ�Nb��i�=a�"����;���m=���F�뙙���h�oT\g�
�U�t:�.�M�b�E\���r�W����kjm���t�WFU񇽓7z՘���<i�h����&F6h@ ˮ,�2�۹=�A4 >�5L�ٜ�|�L��"���Pu;��r�|-Bv�)	�o��d�����[��ǭl8��{�>��rn�0�����E��p�8P��2����ӛ�����<����+֤��<S5-vZ�Q���
1Be�6̲��7��7����vH�����7��B�8�j�c��$�u n��~�P'q��l��~Zm0{s�
��t�u>�Q�3��k�#�'���aX�"�z�O g�%���/i�5��T�l��I��8&�	a�O��zR� :"uiaɌ�b5��8�0����$�|����@��´�Q�ο%7���"��	�Hz]e��5��k�b�ah���kYp�	-���h��1Ӓ�7Ps���F�sv&8�^�| �p!?�+�d���=�s�i���{�V�h��$�k��+��cB�]��r�q����x�UHl��7+6�C��y�쿟>3h5��(�ՙN�,x��禯q�	�o�|�����(�^<4���?�Y�Fks�<H��X�C������,�W3�֕l�n�2D�N������u���"��@���R$�/�0oit3�Yړ�*ɠ6��
���}��3p���ʝ������i��;Ge,�����������E�Ӿ�2s"�����z� �xU�� ��m2'������f��m�/�P�΅�ҳ3���k��42}�\`iKP/R������ay�Q*G�O��RAߺ}M��I�������Ji7�`�V��ӫ����W�%�u�"�CG�����|$%K�駕y���7?����5|%i�W��
G��t/�nc��9>o-M��)ڽ�9�&?��r�K���+�f���_�Q����#�̞���C��$�ԩU$��'���-��B�ʌ+�Ʉq�G}R�cp���:ب劜C6zK����?ʙߦ��#19Z��O�u��w��I�%o��0������d
�E$gשNt����f�qʶ�����ZE���*��żc�(���RG�xX�	�	CtP� �ͭlR��{���i�60��g�L�{!���=�؞�K��+�t8�5�a�27ؾ�<�����ʐ�*fJ9��ݰ0����#T)�4�6���흿�����^|	x϶�P1��g��e��JO�M>�x���-v�����`u�t��r�q��Ҟqh-���NDyĈ����zȑ���i@�_�ϊ��d������T;V��|��B_�W ��U��P{�'y{9��xQR}����'��(x4�I���W�V�fz��>0j!�v��i�X�YGo-�3H���U@���?'����Vw� ]}��1[B�(ޭ�ZG�6�w���Lzw�TO$m�ޣ?~�BV?/B\Ư��C����,�G҃�6��ö�jO1��:W�8AQ���H6�j���~t,��#�"ܯ�0Mp�Bw��8࢟�,��-������������s���QK�ߡ��0)��/�1]Q/>���^����(C�Qf�-�(��W;�y�fr4=��'UQ{�
���"�+�B)��t~X��\I�N٘|[({�����b6�h��=t"d<N���m�M&x�4��l�Q�ɴ�:�tF7=5���,���Nw4�9�O0�{�DOoOS��ڢ�P1:�����	�;�<)�͘�!����DτN�s`�R����\Ċ��1�a�8��k	��;��rvʭ��~Y�����T\]xpyV(��ufm�?@���V~�=��d��	���A��8�i�[����-�ծ2N�p����Iڐ�=jZ�F${� )W�� ��6��&����Z�8��H��9�A�ۅ�0\q���ҹ�8��El��h��}<��NUR^Tx#)��^��i� a�I���61��e������_�:gڻ�]eV�S������fL�0$N]�ΉA���u���0n&r�+�D��HJ@��5?��(hr��A :R�g|���V@Y�m?���p��*��1R�us�~Dj�);ǥۋ�K���Z�d���v���*HQ	h"e����pw2N�;�dD+��Κ�j�`���@n˓��I������w�p#������(��0�
�t-�2J�q_N�xah(����v+j
+�a`�4N9떷<�KR��y�ڮ����MW+�,�Q蒩62�$R�s/�{˻��i�(���z������(�j{��&5}4L&�m��ʜ�˩?��W�|V�ʣ5<�bN)�%��:	����`5�;���"^���h��G�Z�VP��<�d{ah5�g�9�>P�-Q�X�m)'�OU�?�2�ڂ��~uve�@��b�\,/��`�LC����(fۛ�q%{�v��@��B2Ep58��^9�`t"@�@�|�u���_����/�׆�Pl荜�LSg�*�D͜�P;e��cQ�Bf��-��!i�7]����o2 �Я�3�����>-��(�r!yAM:�1�ͪu]\ j�k�F���e���&f�c�]d���)�V�U�����Ǐ��@Y���Ձ�,������[�؝���8��̒s�5;@]�1�}�*��P�W���Cϴ`kKx�GO�Ii^f#�#{z9� B�kC��g�J.�n�Ճ�m}�aGx��~����.����r�[6Go<�0FQ
�znr�پjiN������J�9���O��E\�Ԕ�z��S(�XB?1X�YJ�z���CQ�+nz��`8���%��&��۸+'��s�U��av�}��Ź�m}�|�̸�{��Mꪋ�bw�66Q/�y$ĔU�L������ ���)�V���2=.�	+oL''%���+O��zw?@���ԑ���:a����s�	c��h�
��6�f��q��if�4�h����e�n��r+<�AuBu�\Dͪ<"ymj�74y�9����!��w�tֹz�wӮ�M�T�j씆��#�V�,�j]��7�m�;>��w��*�ŧ�m,b��&D�Пps��;�0�%[Z�y��N�xf�>�~����F�a\H�P�8-a�"��{�/_Eũ��!��\|�V����^�F��1�0%գ$W���ET��(ǒ�k�0B����;��.��2�d���f)��=�K��^�#4,;����~J7K"N����ܟ��3(�Ine�����\�C��'UB��i��थ}��6�יɸԸ�E����O`�*R	�����'f[���+T�i��gZ	��z�����O�������D��u��V�Z5�a5zߓVO�I?�u�rG�]k��G�f �2�E����=#�b�	�'�'�7i
tI�Ͻ�i�RV7Lc�m�T��snS=��8��ip���l���A�%졈Z�m�u~P������,�F�T{qR�"�R��S|d~�Y�e0�QQ�Q~��x�DY�N�y�������-9��r\x��v~~ph�'����;���.���'�?��n�:�j�����[F�MV�#�/�OsA�����'?*cB����O�3N-��No�|�}L���a����'�'# 9C�f���K�*W��j8��T���^��`���)��m�c�ҭ�X�J�D34���S��[�-�y���2�CzG>�2uN���ΪQ��R��O��z��P^�g�YXk:,:v�%G$��W�����������,Y��g����%~��A�,����>z]�W#��L,��_'�d��o�c��:�8�~�Vͦ;s輊Wb�;t���̾j��䯚����d����6��@RS҆�l�u����ӳ("L����hR��@���Utv��1&cl�mN�&{�LƋK��?����EsJ8���uX�ow��OI2��9ـ�C�����:�T�����˰Z<)�@��1N�d6���o] d�3*��!BMB9�G7��1 Y^�,�uR�m(k��Gܾ�DcQ�y�̀����� M��)i�}�y2�D��g� �`^(��P�d@�~k����se��#�u�8� ��Ǆ�����B�v-^��-��������N��h��� H�H�8�8:]%�?H�mb��}xN`5�0�b(F�:H�f�Ă�ՙ�G�;�~o�o'j��)�Tё��obEW>������NQ��}#��(�qoť�2�s��l�'2P(����$�br� �0�����B���)�z�"�����
La�3��ƄEś2Pv����
l��R	 T���z��q��s�]�'u-'����H���̠�n`(���z��*��ϋ�s����t�x�Bg�#�HhE��$��D
O�g��E�+Wz��IE��CW�q֒�w4�7���,V����̷��u�j��8���}��'�Hݽ�:�]L�8`��Ð%�:��%\'�>m��G_������Sh3���[�3��/�=�9�f�16��>�T�wb%�����}�� �1�Os��ۅ�b�����*KxH�o�)-�U��N�0w��'^H'�ůZ��~;����s&�6�m�+PѢ�`�����gxgv�|�i�=q�#@�Ml$}艮3�%}I�w�O�(L0a<6_��%S��mI$�_	�l�!�`@?��\V���)�<�R~��,�u ��F�Jܠv}t��d��j&�6Vvúd�f��,ɠۂiWS�����(\�i�C�^"n+�ޗ��hlmY�ǡl�����`�ha�*�d��z���v�;j�S�An��>�W8)ؒ���qfff+�R�xS�	z$�����X�x����Q��꡴��?\�i�b�h���_�3�ԙP	���L��h9�M�~3p�:P�6L}��y����D|ʭ�6] @p�4m[���T��R��+�e�0Ë�1cȟ�ȭI�i��+2uj����S���@ǹ<r9��F�*F.�`��)v��g��������ɏ}��+�f����F2�`�Z�q�F�?����l���}x@�ĥ���׈���eׁ_���T8 �\3ߙ�Љ�{���cF���1¶⥐��C�ӊ�Y8�`�:��Ҟ}�['O?������']�@D5IX��ԍ{�]�4~�M(�������A��	�{��&��G����o�
9ʤ:�^RJ{������Ks8�qt��d(L,�c�L ��8�u'�?���:��:�k��{I�T�����@�Q[nh�d�����/��s�#�m��6d쉻F���M�Oh'ʜ�^�I�~�3���3V
rKCD̲������S�����%j�o�F���_�.t +8����*�R�8
�c��r�Q5�Sv�U0-�d�K��o�>���v�Ǒ����|_Ni�c�Qa�h�uR�s��_�7'B�?���Y�w����\�A��?��HԠ�'��L~l|�I�fEޘ��H}i)��5ʱ��M��ˉ�R�W�Z�V����V�\�b�2'f	��S"f����о)7�W"���Z�qL$���B����-�#������ڼ֋��E�@ؽ�Ѻ�XSג��ss���
@4��%�t��/z���!����k��}EÖyyS�d��7U*$f�����7�7���@Օ�w?R�}� ebn,�1�^F�n��?uqB��2Lk@6<��S:`�M��r�'6x���\������qO���~��{�	�	�����S��A�w��c��C���j�����b�ӸG筮ے��_����e`G����'7�����FQ�8��C��W8�T�����4.�׸Caz]��G{"pu)�Yk'�ٯ��&��cM�E�Ši�z�� ���RP�#��������wI7d�y=_s�����[P�Y���~+��ç�r���
�����`�gӣ��I�3+ %2��U4�C�}�a��+l{f8�ɦ �`�lĎ�|��c�E�W�z�҅���׻�T��x,�t�w�r�Ʒ�<�"��w>�n������H�>�R�J��}|v:R���^����� �O��������� �l�hG��ϕ/���-ӡ78#.۞n6�A�D����SB�&��b�P}S�f�~���2o�--5D�����#���F*��˪ͭ-��P�y��5/�����Q�"}�DNM1�V��G#��p���#�>�͜�;�6Y^�9j�i�F�S������b��yT|,������Z�6���QR��̲rc.���-��F�{p���_ ��!��#ʱ���"$rF::����ż�g%\�V�b+w(!�馺���:��3�y�������l��|�fM8g��v{��O\,��Ih��C��xձ�KU�$���Oڌ�c�����(u"�'�<��s��+aҢ���rhK	�2**EF����4V�#HӺ64>�r��J����-����v��X��نƴބ�`�{�x+�
ѣ��ögF�zE6w�7
[f�+cqY;F2�u|����qи0�5��}�=5�@�:W��s�eU������x3������EgA�}/��H�TR�ڨ���H��1���L��޶�����txm5p�Đߐ�gV�]g��'�Ѥׯ�;S��^d����0x���m�l�6䣟��	���܃�b��w��m��~Cբ.jM����<�z1^�-���~�xt�.ݣ@ ����!!V#B�
R/�A��z4B��z	��1�5�`���eu��(z@��NH
���ò�}1�x	�]#n(޶���,�C]�m�UPM�8����]a:6"',ٓf��E��@��v��O�Sa$;�Lw�W�^� ���<V*Yj��b�r
8H��J�as)�Ã��i/��"�s�����G�P��CN&<�3	�h��-g�s�F�EW�5���>���J)��`��1?��U�X~R�̚���a�~�+:nL���"8��$�;d[L�����4c���ܶ�Hǭv�{q�co7D�ЩH�D'c�<�ԭG��[d$�9�!�E����63�`�be���Ky���ޡ{�����`���M�W]Y!�0%���0��	UpI������r:����>f�{����/�q�d���HT}��J<��d9��] �R4�J;��ƴ�@A۲�G��1�r�3�7�s���/�J���>���X+�L������p%����4����5�
y:��N/T���$�GTf9����ӷJy����׬�	Rm=���+��Ia��������>9=�]��CL������������P��{n��>m���Iz���.�ᯮ�1�ަ�=��)'��]��K�B���4p�U�R��ʤ�I�w�Y2��b�O����7&Hċ����@�U6�?��_?T}�
��m��.�,�W�9#ЫWNV7���m4�4%�ڸ\� �M7���b�n�@q���RM�UvY�N;ꑣi���̡�c̸��%�kU+�/d����L*ND�CGN�ؼ#�󾆔�S���נ�7e��l��I�&�I0p��߂�Oo���m���5vϲ �^$z�v�s��Ro4����xj��N���1j�ӑ?3����Ŷc��K�QA1DT.�.��z��5^�݋Z�y�X���m�qX� *��'3�ivԎ����4 ��q��_�nѫ��e�~C+�Zz�"p�� 6���>�?VW=ܩ�xG�x��H"��j-���=�;9�+��u�c$K�����:��.��#�2���Ύ���,��XZ:�<氠���p��n�n
T��;��a�%������Ќ��1���^��R�(��_svBM��v�@���|KRA��0TA�r^U`���+H��)��a���"o_L�R(����ePI�Ahl �}%�,<;�vH���:��^�dE;���B(���f7~3���3-�1]�O���;Hr�p(n���2	�b��\��e�~��B�<NدT,8Rq
���h�-�A��{<��s(u���7��GD=��F�`^H�O}�����A7���X;��6ū��e���V���{wؕ��%�����}���lIy ��N�E�[Zr=m���m&1�A5|�]�m�\����^������u�/%_C�@6+c=3@����#f��!c��=���+]������8�Q���<ݼE�7�6쑧�]^��p�ي��i01�h[7���iG~Ѥ/Ps�E�p��6�/fH����T���:���Z@�%n�[=~K���y����fWvt!�v�������ɮ��d�v<	�R��[4Kk�G6���<r�6��*rJS��4�>O�s��2�ر?Z���6�ι�ҝ������5G��i�P$�+"H	�^�25w
�*�5!qW�����_�i�,�y�5��y���pP/�������T0��%�#E �!b��BV#�'���y��H�w(����Tǯ��!�e��Z	����xF�B��y�F�p�ogɞ����>��)J��	�{�����opnz�v�[q
�
�I�0�����2�`�P"����b=�4�f��l+���X�\�8E�,�j�s�QUm{����bi+��7%c[�I�;$�I���MqP�J��#(�y�F��x���j���P�-�?y�R8�լ�3����l�%{m���Q�"��j�G�Xd��n�J��~��wf�}_�L)��������M3�Z��}#�<ђ�Z���b��m�����J���~�Z��1l�����Ǭ�]b�gA|���}�'�-�]%��F�P*J���l �n��m��7��Ғ���H721��#�}��FFqmj�$9~�G�XhMx�����d��ElZ����e��\/��1�y�,�hk4*)ƥC���,=*S���-÷Dy�%�^���'+a�t�$��I�	QP��޺��ol!��l��/u�R_�B.ˎ�V��@�+a��>_.k8��7�
��ڏ4�  ���5��(�U�6��^޳i�#βAn �Ih���W��ɶ�E������6#.�>1�8z�'��\�5E3z.�R�g)-)q�D��A�&7�m��릫��MX�?���h˫Ro0�<\�"ت7�s��) r$h�N����[>*W��R2 _h.|n����3�ݍ�qN^\����0s\�Y��U%x���������
	F�N���m I>������G���4��Y�Q�\��F�Q�Ŏnl�9��Ic9^����77��+ZG����P��X�R�%�¹%�y�6eA���o_\�-��'� �h����r�ƕ�)4=��*�%�շ�;��5������r�Җ��W�9ov[c���bw�
;@�G���Af��eQ�H�:���fꟹ˶�ǡx��b��Qp�C��ShO}�N�`���
4Z�'g�~�ߏ퇧������w��ˈ0J���#����9��pBǦ��Q߉~UztLkD+��J��1���ND�ssl}?8��$X�(�t���nס�8L�_y�;�Џ��jH-�\:�~��4E�'B��)��E����,G����v�?�sD~�8;�h]*����R��N��%S ��a8(�
N�|n��
��;�����!�¦�ᙤ���z���I�be8O�$�^��!b�)>���$O>P�\ɾ��4W����V�� �*���S�d��M�e����kd�Q�53�.μBP�1[�2�[B{x^�v�2�Ħ����AY��n�,�kt5a�'��8u?���|$�����OJ	6ʿj뮡�?������W��BZ<dn�˫<���Vg[�]'��8+���`����V���0���#��\���Fy�*"s���,�i���[K�.�0���P�;{��AƵd������L��1��� I��ύ����$�j�Z�!�F�i�p��1�]����3��7���y���ǯ�kr�*B�(5'��
�@4���S9k�Ӹc#Uh��G��	�W������DKg1{�����p���r_q9��������'��ģ��Ut�F�h~������S��>�3_�p�����wh�eޯ�o\1w�}�B;0\º2Xm89W`?�S������:�\��`T���G �'�,l�U/��/5S�s��N@_�\��g��=��*��R0>����T*��|ʳ�@k�?��Uϑ��:�$T�v(��΀7�=�ۋ�ɁP;���U/�N���2G|��$�U�|-O�C>��h����:Q`�ٻY1�8(����t�_l��[s��RA�o��@]��3�v�I�_�=�(�g�����x�M�x5%�<z��Z���9��FوW�����F(:	P�h��/Ut[�J���|�˾�5hq7����#�N�u/��"�31v���j�粻�M��%kV�m�ɝd��Ljq��+�yܔ?��D�� OD��c8없z�-�h�ף�ec�,<��0�ܫ�t���E�S]y�ܦ��+t�I��k"�א�,Ļ2wC�P4���ǝ�(�K{����J4&�ꈵIJ��#�J�]g�b)ݝ
���ǖ3g��˩�|	�s�[��-��Җ�P�Oa�q�&��%�A��'� �2�=Cbx��V#/���4��Ms`��gw�څex�$�LvpS�V<"�g��	ed�O�nƤm�����|�V�	��\)�x�[��8�v�k�)���m�����=���~>���ه&��`��5��=�}hT��6�%f�#���/��hW�d�q6���Vpa=����oo�!D�uo��axG�@�z!P�*����f&�����+�s�8<^�@&�>�<[{	�^^4y�_����d�x#�-x8qT0��c	7�k=����� $�C\~bp�ե��m	�;�Rq�� ������
�mbFF(��	�a��[�m�������P7��qՖH2�����s!��nP��N�^�v����fI*����av���I+�p�����@co�I����i�	2�&��,��k/���;ː'����5���\@b�Q7՚&�i��]�Վ(F*���&�����&�#�>5��z��G�ǜ�ND���n	���M��$�5R#(��C�"0��CQ�=1�$�F����@�T�E�������ry���	��t3U���_QbL���k��R�u.E�w#�pd��W}څ!	� ?��@��룠w��T�K�6��EE����*@\�\������
ѫD��5�"�5��.ftx�b��"��#��=py��g~_©VR�H�{����E�ė2�'��Lu��&����rՁ�(���\MR�k�}�caJ�Z:�o�᧘%r�'��՞`�������_�<����uC�xK�-���fK�m�|K�m��/X�k�X��0�=��j��4ZZ�/��<!\�D����2~I~�`�.�E��pW��ǔ���j�4Rj���1s��������2Pޭ�_���y�'w R�,�uw��cB�M�qr	#�W�R�ν�k)h[T������n�,d�S+�/E��tH�Q3�s�9K�~��B!��M��=�z�;�C��=AJ]`&PQq��Q�j9Ou��P��8?w�CN%�A��פ���Rǫ�m������O��޲4;��7HB��O�0֙�ؠ�ш�E�T3&�J΅7�� ����xqJ9!gD��yj{��$.��*��>h@[� ���_�4��������'2Dk���4&;�@a�u��jm�B�cm_��~�B/a�?i�4&�u��mq�:ĿP��A���x0���^�����������<��Nڊ��z0͆z$E{B�������!�\8���3���(�s�>O��/�z�//0����E����cP5��VAG؃��*�}��&�i��j��M;���T��P�X�B�d�?�[�]B�#nW߇�+5�A����{/�9��؆훧3�D�Q���e[���kZm��>�
o'H�Z�|�"0�J:�d�|��X΀L9�}��DU(���狁��Y+���	��y�$���d���(l���s���S2�꽅9,����s�9�%r��W�`H���4��ʘ���h�eO s$P?�)����I���Sۦ��%����Ǣ>�G4�B���U&�JU�Dq9ao��T� ��Lό���C!)D�TЎ��t(��&"����м���PY�2z8'����KiC�e�;Wܕ�j��ĵ���PsF����5��X͔Eb��=C�h��Y�H��I�[�1�R��(R:�N?f��b�2��GZ�c���8�oy� ]k6X�W�^Wej
"r{.`d5�g�fܑ���k�ܑt.D
�t�����7I׭�0yW7�k�!54u�)�^t@t��:d�?˗��LW�.��q����/5rګ��
�p!ƫ�H_���q
\K�s"��!�D4���ǟ��-�GJ���&N7C�Q�d/R���H�j�]y��-������J�U���V#��G77�@�`$䰘�`������ �:1wz��bAOI����F��k�R��"�G+�g���&TE�i�x��6�mu(�$y��.��η�� �!����cP�Uh����&���ml�y�ƃ%1m�m��כ�J2�*�uߔ�$P�6�^��g�9+��L�K�������� �H��K�VF�&4Ԝ����¥�UN�O��0����z��-h��F/�L�hk����"���$S�-z�����ķ�y~�(�T�Ζ.6zN9)���2�c����_����v������Xe�k��2E�}�S�Q��?<�,��� �k�|L�*r���\FP���^�e��#�;ܴ�#�bd\r�mW��A��C6�c�
/��z�h���f�=��[B����9��w�;E��������9����Ԉ���<R���Լ2s8g��1���݄�p�b�ZQ:,�c��H��m�,�c!�?VK!=_"8�������.�*~�����v^��ߠ$W�Xv�G��i�c"�۹�
a�(�6��%�|��Asi��z�V�\'�Y��O�6w4��!#s�*0�L���]Bpz��S^�h�K�<��Ūy��iQsG�̺|?��o.;V��ڬw2��ڇ|��e[5!�_-7�6���Y��Q{��oP�\8hZi���B�8	��q4aQA��]cZ'r���>ɞ1����e�>o�:.�?Zŝ������~����e���^�׏cax��4p/����
�����c�-����hc�tm���h�MD���(����Zd=���r���n���_�V�<��,*g��p	�c}���ߜ]#��[�T�6Z�m��#QF۶����Ԩu�ٶ���-��Xn.��&�#Bt���T
�@� ���N�� ���Yd�����e
�:ూ^�<Uz���(���ն�'������ܘ���@���s;K��y�&t�R�� M t�G��@�Jj�^j��B1�"^c�xQ�׽�zGP8C��U!J����$�CP,�9��X�#��Ǵ�no9��)>}� �����A.�H��;�����bDs�y��B�/`��/��i�ģp�{ۋ��[oN�/M��C u��n��5�1�uW?�4jۖ��VxZDi�����O}�uǿ�6��b���+b��c�,���B�\)��;-�7(��g��@����j���<����8�(���u�x�n�����:z�H$h-��˚x5�%t�����;ѐʍ�(���"te�����}"�7z�8���V���H�xkB:����w[�UE�
oN?��
��t��̙�@����L�_W}�]�{;����\@��p�ĩ�+�H�����8����-7��(��	��1��"h�fD]eW>���>hCl�-���ׂ41M,�y�]B�Q_}��W�(���6s�0X���� l��k�-nck�l���h�F�z��;ˢP�W}��0�Ə,qoo���]�V�E�I� ��k4�͆�˭9Ͱ$,��H�vE�Ѵ,wf{<��z�#�����Ie����r��豲��;lR��}�ю���'U��wt�"l���V���=]�ߥT��u�����|ZҰ��3V��m�K`=�'�ხђ�k�b3~%
��ZP8n�O��N6�}������ ���p	J^�x0XD��~��wv�� ��#��R�0�|����/��*��˰Ud������ę�R���n����jt�P�G��"WI�-���,���I?�+��WۭR.ظ�Q�Ð���.���]e�uV�B1rj"�4Q��N��������7��
"2a~.i�m�Mt[ߝ/[�^JbKx]|�_;7�
=��7U�]&��J$.�\��fc^���9tG�Z��4��rn��v�n ���0�~2����5/�RC�bDѸ�	�w�|���]_��V���ZjM��37��+&��4�^M}&��m�|{\\�4����Fa֤řPo��O���nE@�Å�i�f��C2Y�f�[��H�7��}�D��R�y�s��wW\[��n;6T����!ĭZ��C����_כ_�]����(F-B	w^{x��a�.RV&��_bA?��|L�S��:)�B�t>K�H��R�BB��+��\��o���>Ff�/#&�Rn����I�fyl��H�1�hR&|�)�2��k�H�%T��:	^�婬�Y���eٸ#[�~Hœ����Z��E����(f�+I�t�Q�rl��
OGRj�VMc��۪W]�6��5 CM���;TO7[��!��]���B�el�8iCS��
�a���� I�fh=�f��׊����[Zȼ~�z1N��v�/_�͙�?���X��).�x�+�d��Z.�-|�Z��J��ŲS��R�l�6k�V�{-R�&g9�Q*`˻>ҿW��Ԡ�ۉ�ճ�`S�a�N҃c�0��אd{�pf��!7�ܯO�����P� n��~�N<�ʙ�@�:o7/�ֿ�����=m�ܴY3f�Q��q�B,Z��Q�_GN�Z�g�]vC�"��;t+��$8dz�h�M�<����D-$r|>5���o��Z�g�xIM��ux,��T�?�".F:�@P��])z!��S�Jq_񢳛t����F#��g�G�txxj'Wۂol�����I�Y �`)bI�C-k������*��J�)��Q(Y|f|=��<j�\���S���q����]�2K�O��.���آ�H�ޕ��D�2�2�*Y�pP�)�B�ys�C(t�HEn��xF�����^z�G��#�uӒ�����k��r+��m�������(F[�J�Gs⩂�-��4���=c+���k�^�_�%+�%�y�������#����+~�4ڹ��Q�AHE�wsva5b���yC(>k�F��)�
�	�2ﭮnI�] �9.�A_n�Y*.am�B�i�q���3��g?�^�4��`{Q�%w�~���E����&=q�#i��~�nY׬(R�3T�����"�.��ڙ��~�B�rF�'ZE�Dn �W4-|I�Ny?�������&HH�g�?b3�������Jvlbs!Z��|�q��(]m�g�<"x�rC��������)7C2Ѓ"�Τ�ǈw�	��zu���$� ���W
��}��<�J�I &2��W�F��{F�C�$]�"֊�Ƭ�J,����a��zNi�#�_6�BhqN��텦��%银 �g�]�k� O£.r����_}D�E->���L���ۼڄ��&,�� 8�����Y�� w���V8��I�j(ژ�7Ր�Q��Vԋd8�%*�� C��"�F;QX�؆a��yW?��D��. �,
n�����
׺;�w���,�%bA%���b�|�.rls��v��ISf�]8a�M�/M�B%E�kv��y����
�}۶���:�9^��ѡ�0�D Z�mќ�O8�u�c4	����q�l��w��#+�>Vk��_�$�w����=i�7��6�N����D���K�歾Rþ��63ˤ?���kS[��J��>8��Q�ս�@�>�R�ٕE��92έ9���:�z��erdT��re�d�1�,6&��d�~�X|�t�tPc��7"�1��B�xo;��`. �`z��|U[��0����(:��V��&��M�TL�휖�l��r��w��>t���4<"8���Px��놳��$_9��:r���I����-�E��x�]gw�E�w�h�S����6-�h�Ŀ���@@���-Ǫ���[L� 2�����m��>��q��AjPPlQTj��[0�[��c��������o<`�AՕd�
%�rN%N����(r����m�4������k>��>N<}y�LЗy��08���w�5��@�'��MNo�M�1]�5�m�L��#�Aڽ�y�U9���i�.-89T��� ���s�I�~3���:=:�ӉN�I �%@"V6|/U�b��B�9n)#���hmz�}4։H�#���*q�Լ�ՉQK�D;u�x�5O��11h�Xb �h�^^Z!����e��v�ݭx��ƫ�s�����9.��T�]u�[���ǚ)pa��4���mCd��9�RHD��H�5�]�1��x$���,�qU ��~|�Dݿ]�ak|��.�&�1+chg0��?�?���d[��K�k�~�)I:2�&���-d#5��<��	��L7�=6��7�����fۭW���r�yC�Ŀ��W��&�� �	�n��0��q�n��W���=���ӕ�	��([CE�G*�#��`�H2\K�r����`̶�@�9�Ǵ#!9>���AXǰK�]ib~Fo��pl"���d��������������1B��`�	?P��%]��?yv�sL���E�]~����$5���d�R�&J�$yL����T�D�(j�-T�*�N�O��S#�=}ୡ^^$W8��xMZ�W�Li���L���T���K��a��E�k��ñ־��[��6��`�Z饷�Ji���B�븘�T9h���QKlZ��[P�ur�o .w�0���+/�~'p��F��x�e9�ξ��6hS���7�7#�0�e_��A"&�]�;O��G�\c��P0�WΘ���Zk3�~XM����ha0��eA��&�Է� �9�!]:��Ff�q�hCBbdц�'U�"�� ���-�k7�7u��<yĲ�j�)�~�����$Ew��ğ�x��N���A��Uz��{�+� o.����/&�����������r����q������v«��2w_�]��d/h�Νi�����Ilp���O����4�S>���R#"������|��?�Gip�UM��a���f���aX.!�O�S
��پ�N�����"&����Ê�M٠)�����5ş/w5;)�w3�do۷�0���G���w7���~���c��!�R�diR�-�kT@R���_��!lօ�}�:|�*�랍�$��!q��&�t��� ܶ�'���ޠѨ��c���S�KO5!��X~�p�Z�u>^��.b�RU�R�S�
�	��CJ*��"��ʃtE�l�y�%V���M���*@��������4H�O��k��u�eiϻY�y߽T1��M;��:��k�.[wn���W]%�ZH��/��T�U[	���~�7_R�{���&����9�������d
_�OMP92;u��o�5�D��a��g���lN���T,�r'����,Me&�)�w0t�ǥ%������w�{3���J��z��X��ɡ�D��[��j��M+�j#R�~4^#Ӊ'�& F�t֍ �.5�N�(N[Ri���I��l��]k|T�͹@�/ p�𞳥�W\8����**���&t�g��I7�NNÖ�o #�K�\��q;��M+��5�� A��:�W�N݌����l�@m3>Z��ha'��s}�-D��*B\�y�E����f��Su�aNQQ�hU�.ޜz����d��oIK��:���Q͆_+�+55IW���v���Ţy�����%��=�� �L!���}T�X�ִ7T���=�9�����/~5p[���l��r��*�zhSrF����@������avf�b'�=���$��X�3�uԨ[QC��dj��JW���ҕ���уS||@-���E�5S�}|�9P�qdG8SFҤi���x����ΥB8��bʰO*Hg��P��δ�H2f�?EVp�ĭ��y�.$�;q;���s�ò�B=r�\��籫x:<h���2Z�{
�,1�MMT[<-�V�NWʔ9�"�}�uN*�V�NNƩ��*A!p�$���ޭ#���[-h��I�B�]�d]`x�H(U���HrۄHJ9�;Y���sXe�pQ6&�m�\d_Zdo���x�م=Q��>���.�6�U��ۑ*H��t$�9ܱ���ŀc�ȯ�+��u��7����
Ѧ�m�8|��hy09��'��J����=�Hq�k���{��x��l��f�i�ގo$Ë$� 8�����0�{W 5I��VC�N��ZI��O
)��3���Hd>��y��K ��S��n�p��7��M����	�)���;���ODkÏF��Q��e��}������*G�T�#�s^׀��L�����y���!4���U_G�2�S1�W�I�]hQ���J�2M�L��GN�ە�3����e��*��S'��cd���V�:jo,�4����
�-L����w��*h���)�/���N��H�k[�p0ö(���~i�d�d�uhs�f�BT@����ΡBg�ᣒ�V5����2�.�ϝ[B�a�*?̯��E,����V��YG��.%�?٧�s�M0�Z�u�{�>�mI>�i�%�uW�\͇����ʉ�\�I]�~��!@;�����������F$�o�	��ST����=&d�h+�)[~K��Z{������y�4F*�p�.;����u�BLi����%"��p�����J&����[D�w���z�Ze�E��x�8F�x��ؖ�`�I�E���G��a���z��Z{T9W���G����֪�`��U���i#Z*�=|�'�a�O���@�CO�;e/�S<��m�i��D�HA_���?�$)��6*�hdi񗋽��;:\���F��A�E.��-�;���mL�f���&u�1�$���3]T�w+)XX+����#��,���b/�ݑLVt����<ë|c�m���F`1`���f�h�fm0�^|w��� G2~��O!��N �ǉ��{�yse�h
^B��FdEjr����ם�a){M/���¬6��q�q�`'�ά��n�uRADa&���I�J���'�'��(L�I�*4�)��U�\�c'�s�lJy�#�b�g�ǉ�Y{Cċ��Q��E#����nE��d1�X ϑ�_��Hz\;���uS"�$�ڟsZzZj�.�ͦ �Z=f�.pViF]ȫ����u�B{��m�rN�+A�RuK��!0 ����2At`>A^*�������I�����H���������<gL8O���n�`���/�ߤ�n���[I���W$��P�I\������<gk��Q01���ź䠻�c!kExJ�&8D\;��I��D�z*�~�M��d+m�Ll���:����G�7-�,�6R&��f�*(���������;l*�cdSo5��u�F�:Y�XA�.+\��{"�6������)���y����Ջ_^�nɨf���	
$�~���8|6�)}kP�?�3��ɟ9m9G��-���7@G�z�u�9YN�;ܽDA�-ٰn�;�2��հ:}nԷ�u����i�4@��c2�̉��&Tb�����McOt7����	󶜳���{��D,�.�.ʜ�e!l�B�W�����x������1�'�Z̺�)����~BAc�e��sJ$�b���]?*�a7�9�mO5;��jhҿ����:�Y���z��>f�mo������d��h�7��
t;��%��%�J"ѫ�ژ�b�Y�t�ƒ��i("���Z��+��7=�Q7���/jl�h��xn,�3+��b$� ����3�d�4@�v_�� � ��;��x����b�?���z�gE����%���$-�_�u��:�0"��M����xήW��Z���f����˒w�����~�<��&��Nt��m������[�G+�!����q�ٮ�Vx�B�1W$h���鉽w}E�O��"G����:����@��?1o\A�4� �v�k���z�UU�p	�Tհ��x���`��G���>��J��@#y?|g��fݗ�����|m����Z���` �x���.�ū[`�e:�j�7:���ɸj�����;ď�
��B�i�����L1�<�A���HP�8��%�j�^���+ई�r!�G�}�ᷟS���!����p�椡���S�HO-���)�(�^W������7��>��?�Xh��16�}#sD�8�-<��D��j{9+ծ�;[Msy���sĨ�S�=?�0f��I�w8=���[�V���e�i���Hz�.��=��گ/�� ��y2��`<�n���~��$�[g��}�"m;�d�O�Ľ�`���`<�iՋ��?�3#T��>$�M[��܆Չ���k���ӡ7ᒤ��!P!����i�f2�nf;	���ֆNW��w�1sB�s�L�"�Aj$D�uĽ˟>���y�R��4!�D�:g.��w�7�ձI����e����F�Pt�͢�K��/���|-аW�N{�q4��Y��8 ~B��	 �����@��U����T������9�"�����vZ��tj�6�)lƐP��@2$nfH�{͈|귩�c��
x�L�r"7�e�N~�@��;�z�ݣ��ݏC�3���:;,K94j�j{��]��3
I��ጕ.ˢ�FIb������"5}<�嬆�%P��yp��n]�J�M��Ub#.h�q�<�@�&=6�a��a;�q����$��S��iQ��k`YKv�63��w�)�l�&��~Z���Fن?�)��шYn*ʨ^�L~Zl;^���H`F�R��HP���f�|���+H�1�X�wU�~8��e�h.��ǫ)k�����UWz%ҥ��[�rd�z�|KЬ���E<h�=�jq��Vѵ�lb��J�1�IS��>kw����%�`^x��;?��5#eg���<p	��&��$�;��gf��~���(��g�i�ش9K��|�#K^KH�B�N~Q���J"�}��Vi5���ʊ(%����f��ɺ���W�+Y�_?�֑���b���Da ��4A�N�*$������c�rZ�cOۛ`1gԖ�L�;�!L�)&��	ͪ% ��Q����Ǧ*TÚ�<!��/
W�g��շ�9QXM)u������D�'���^��;����N�O(�oC�b��zq#��Z-�[�<�EZ����N�D���j	"K`\B�<�6�tJ��xT?lU�-�`�Ne��44�5G�鹢�?��|�j�b��?��|׵�HpБ�딢�<��3L��cT�T.h��މ�����];p�)�5�7�=:�n�a6g�d��ZJ�%��М�:U�3}+{�����_���x��!i�_�eAs<-L{�f���^�$a�"�t��˧���\�/U*��F>=��[��jb��+��sP툅9SרZN1��ܘ�)��.�M��&M����۲o��&Ty�tut�|��6f��%8d�Ky6�U�2�PpK|��e�^K���^�.�&��t���.�C��q��x@��RR�����%Cn����U� ��"d�}QP3N(�E9�k���}A�E��mU���fi���n�͓�Ka�%�WG���ry��	��n@���ӑ��}-L(>"�ZuDotwFO(*>�w�q �c��>�rs9�7�	!Hp����_',~oQA7�2 �бX�� ����JRJ�wC�g8�Fޢ_�]&2���*[j�
���mӾY��/������O��^r=����v���$J���G�O]'yY�sAf�kq�՝J&;X����~�y��%�#|��z�ofs+�����?T��D�~k��nRi5�X�~�JL���������Z�������3��{�+��v�t�����z�������~�̈́YG7�����0���{8�^�U�֦+���mP��V��{K1U-,I�u?��|Gݮ&�-��e�Vɶ��P�Bވ*�q��񢛞���!�5��7B7���H�]S�	^l"��*�RR,|���+e�d��� s�T�u8�c������M!)<�ݿ��m��/�u_R�]{�H?��U(��%����E�Ԕ۹��-_c�M~OLT�|c�����(I�P�N���`A��W ']����Ih�d��~���=� )�:��C����P�����p�Ǟ��ʄ]�>�sz��:Ǭ%��F7=r��l=�權�~C�2�N:��([J1�܌I�����|�/:�U�B%JWS�'���\���4,��Fd�0��{�̢&&3~l>���(�	G� R��qC"�xo�������D�mz\"����y�i l)Z�'�5�Y��]@y&��IZ��$nm�	B���D����@�L���l�ؔ3�i�y7m��e����4�dv��$��q3�%����'�
�P�L7�^������FG�(�������@J�0m�c͵����s�;����nNJv���O�j��`�AD���03'a�2���l����ha8||�f��0�Sw���%*wwMX�&�:j�Ϧ��{��i��}	��\�Ç��q�(� x��V��G �b����{�<�R�4}=����8��wZ��On��j�M��U�.�����Z?�&%pwu��/|m���Hj7��S�ݚ��R��������N�%�޴���³4:V���}�1�B���������Y�r��
M��1|�������
:zh</�	�
�KmC��h��[�Lx�v�d�n9�iC��^R�\/&0��iĥ�N)��ժb[Cנ��
�K�& �,��t86{�+.v�Ȃ�$������߁�	]�P �>2��5C����L��'�����O#(7f��}I�C�T5+yRj�ʿ�u��2j�/D�Rc����=�K�[�/�a�~�˟�����I)a�[ܭ)՚PC�����+3��IFLI�N({<������ශs�MR�uv늧I�Y|����\PP�ǀ-?Op�<,��a%.~^�\�K�@\V��[�/'�=u�o�L�9��Ԑ���4i,K� П�`&ᄷ[�(����z�t#�Z�.��#��B;1���&�ֳ'0Q�Z)�p��(q�d�rߥ�:8����-�����s/`�풐�h��5E�)S�X�1�Ųm[�j]���>�?%��I��+� ����H#s^�\O:>���8��J蚟ﱦ���E��E���/4�������{�g��8ZH��Hr����O�����ǲ��p�7/z%+�ŗV��#�ٗ��||O݃>qrd�>):ʘ���@�ޚ��B.2���N��[.���]��INعL�N~��`�m4e�1�M���$���D�=���� d%�Ќ;f��*w
%=?�|��e9%	�WR�@87��31�l��(k��n����V��q��
c�]O���v=�{���	M� _���,rdz� eE�_C �]�HoW�oGS���|��ʘ�}=�L�"+�n� DP��h��|���ߟ��QKM�ƶ�Ep��L�B$�wZ_���!*hT�6r�W30�Y"�~Ȭ`���%0Ҷ���s�u�Z�|��P��#h��v����iy\�NnJ	�q�T��jZ���X�[N�I��/�v�y	��A��Yq<�5R�͖��c��Y���|���ɇ��8�ǂ�%����x��8���]��4Y�<��QaU��2�?\I�"]��L�N,mQ�gk�K�$iL�"8�d��,�m�t�7������ҙ�p�	ȩ��̞TOw�>X��4�~���mC��_a��x՗'pSR���>��7�O��~��58��������MV��0�?G��n
��!%���$3� �Oa�˓ԝ�w5`�>��C��e��}��8i'z-NS��I�Ǚ���| %.Y|�]�EP�S��(5���F��+�
~qٸh��nXV��J�"�����0�>74�r�=t�m�ɤP��mEV@K��3�D�O�|�e��sIk�>Tw��Mc��8��b�z���PO	��?�{�5�.Y;�ļ;��O�y�yv,�V�)��Z�\~���5���0�ƪ�Y��Ho�V��-U{|곲�_2��;���/��"���m~Q�T���^{U�n0;���-f,�:لy�A��;��ו4��	�K��� ����F��0/>�?�Ө��o�3�����Gn��Ȼ�!M�J���
��b?���rZ0�<n���:�aL�YV������@��u�<��1o%�.��ݏP�m$%�ܷ�������"�{t�L��۟9�Rq�@1�زB�QmE�`vd��t�if똇�`���?F�W%u�ƻ�1�g����k���A��A�r�B[��t���A�|��E`�'H~��\�wE������J�gEt.j���*� S��KOq^N	��&E�)|C5�+nWS߽�N�xlt�%�m.f�Y���X,c�� E��n�^^�5y�3r��A��$������6�.��{dcu�:915��˻��>�Z��Q 	S�@ blE�G��w;����&�*��cbܵ�*�^r���ۄ3�-�L-�����|�塇7��v����[�C�X����A#�T�]PYF��p8�C'J��𙇵��W\M�=�B(��&t�w.[%۞(*X`5-�ΘR�Y���r��S� r�)�����d�m�U4�0X-}ZޓH��r����s�<q�F.m)�$Gwz"I��c����Ӵ�L��4�W�)ok[�q���p&���y�����u�.��k���Ҙ�E�#�j-���/{��>��bg6�A�����-/�/g��Ծ�ֿ�`���Jm�[�Hi9���n�7�[Xr���+��p��"YБ���@�Q���Oy����]Y����� q/�%��7&�Tc=!�ސ��(o����U'��Y�XP����]͌R��1��ћ��/I;�'��_��л�K���gCZ`�HLj�j��a]ڨ)��p���%[U��r֍�@>ܢ�Mf&��[��6��u����Q�V��Ɖ� �(7]��d?�hf�W����|e����FR�xŹ�r�Tw�¡m]_(ic�BG"�]�-���{w�A�*G:��Rq`�2��Oz�j.�6y�F�:f-�Jޑ*�
3��L�Z�)�T$`����=W��XQb`L�����Ė9P�>�f,��ެ�4�շN=J�i�a<�p)�;w7������%���5x��V;Cu�������T��[�$U�6�H�С,��^���� ���)�k��*d�4X��C'����o�)�	����w�׀�����ʠ�d�9����W%
_��%�&`
"mN���@Z�<y����]�D���Uzb��Q���`?��S�� c�*�fZz�5+�d��X��(0�ޱ����.aS���TG���׏[���(�ԤG��PRz<`��!Ξ�n�d��[�E*�w��S��|�|�����Y�1I�&���[Ù�4릍�ݽҖ��h�
�1JdΨ���z@ƇD�\�Nc�]�G�^��kc]��`��T7-.Jk7��5���X8L�Q�Y��<��/-�Ҽ�s'0��R��x�����>Άpԍ�m��gT��n���t�����6N S?@c2O�k�5̂����1*W���"�tV�8�K�stٺ����;�v'�iw������G���諓���T � ɩt��R�P
N	���e5c�cӚP?���$K�8`�)�K��!�
��_��% ��&[jc�1Eϴ5�_\eܪ��F���)Ȩ2;~����u�&!���5?W����4��w�أ���K�>ؓ備u����i�%�h��
YJލ���s���Fw��>�5�o����ل�a9�q��Nw��nKNE}�ׂǕ��m�ڠQ�R����B9":ǯ�Kc�vh��$R�S_�C�K�g�D'w��\xG�L�֝�c69��.�eY	~�+���sM:���~���I̙Z6q% 4��IXv�?��V̏��JH�T����P��ZB��P6-Т:ADϹ��.���H뮜5������<͂,	�I�hlέ`�q}�(ƞ�&��V>�`C�yf0�[߬�G�p��[P����Z�e�Kr3j}��4S6ڬ-�-�u��̬�=	E#x���y�g������I"��Q���yYc�<z�f5�-j��鮈����	Q1^�R]5��ݯ�0�9����UX��=�Ii���->d-V.����|?�+I}�Ns�F�]�E5���0�L�c6,�]�E։GZ
~�w>��z�^wRO#B�a:�rU��cw{���# 4�?��צ1`�.�_w�$��O�� �Se���FϷ� ��y��+2.p�_*p��^�uajP�VR���Q5�e���U������ ��y'C�~�AG�=��&�?��M0��yW��Y�N�x����$�eF"�zS�Wg��ϭ�L��{���.��4_F��t!�h�z�Ʈw�yr�sfZ�b�i^E���u�݉�S�Z>_�hE��ԫ'ʵ���_�R�`�_��u�����o�/Y��<�x� i�\l�B��6E+�=	�xQ�|�"��A�88eA��_p���Y5jwܛ�_>I�x�����ћM���o	$9�������q2*⩡s-�4�C@&��������l<<��/yfI�*Uܤ���u>b���8������2;���2)b������"?�O���=.p�`2Si�����WD���I���`!j�|ex��D���E�d`O���Sd0ũ�8�$��I5�q����;\}ӧnS+�-7��b�~?3���r���p�p�9���\��bi-c����r��łև��_o{U+Ps^�9"���>#!�C]^��@$l��㬌����п��4u#���1%6ql�)_R� �#P�)�=i<b��	�K�7MN�e�����a2!����,y#�金�>�Ӊ�`�i"�z3e~�O�/Q9v�k%���`Jqy��_mi��>�!��5�2��~W�� �̃��K�N�*�H�"��1�T�6t	۱;r�ԠVu��T��U�-��y��/7<��#�Pd�M_�1惰ԅwh�����J�H��d����(@�}� ����,(��f��E`�S�pB�\����u�Oe~B8��K�x�\��U�>$�Bz��K��s�i�AEM��Ɲz�(����J����nA �Q�P��xGB)P gF�>b���n�w�T�螔�K���Jcr�\=�7�լ�Ȃ�o2�lBl��mqF����]���weqoT�#�Ԥqp���!��F��$��g�Z�d�g,�Rn;���G:oZ��BP�����W�ڏ���S�d�}��>�/6�:���c�U尒{w���J �� ��\F��W���;A�vsl�\oT�[�$PW@6�E�uM!�DI%�\S#�.[q��"u7i��I�ܩ�A:iڅ�s0+��<Tjh��,d
ZO����cz+Mu
���Z�]Šgv��Ab��\l�*��i�D�$���o� 	!�N���ʮ��4��E���tĈJ�bfP.�lO�Z������H�Rc�����o��g���ǟ�E�y����LB�j���HfJ��笎:��<A�}@c̱%�S�Vk9N7�L#d#G���:�0a�0&�֐=�r��a�!si8���kH�k��*g�d��{�o�n��X������g+�/�@�KEs�/��+HK(���r��'GeŰ٫:+��٩����a�~{�5F��XNX@*,>���儁�?���F��h��R;��b|���`kj����[Y6W���A1dd��@J���Di���.Ћ��o�ђo�c���&O��~3��^�����(2��k�#�5�����q��p�/3�Hq7a&JOސp )c(��PW_-ӊ�Ç'a�聆�oA`��E���:���bI�D��	*Ys�d�����l�_P_���s]�N���Cl|���e}�M�����!��j�.�;s^L�Ύ⮙����1h'c�@4�&�t��2�O&x�hWo�1�YRa�J�6����]P���җέ#'�nc��ӧ�ϑ�v�]U�<U�++��I����7�n�{xm�	�C�nB�P��dN�伐S`l\�Uտ�N��Ĉ}̏iJx��b˹��y[�ˌ��v���ٞr��`�]k7��Xb`[��xD{[�=Fȿ��ש՝~���YӮL�`F&�4� �T�ǜO��H����.�{��
�0P;���2�U�n�n�?fy/'�T�Y�E���;j�I��ϱ�B�Y�-z�j�Hm����Ll_�T�!g��S���_�Bǫ�yc�kl*�?'܇�~� ��}�b�^d1�)����F�9��7IG����x�j��J�ݡ�.ՔYu�}pk�����)<Ā�Թ�K��*����Z�a��7�W����~��^{J�f�I���7؞l�ޗ2>���~���<�|Ux$��*5�j���e�}������ʆִ��=��߿N$��6�)!���sQ3�O��n���/Ծ�֗5j�����TC����U���á���N��=/��Plڃ���%9���QO7�2�`͓���B1ѥP��� � )b�Q�Hz^�SѬ(�Jn�L�p�V�}Q���AB-|E��`-j��	�Nj�5lڨ�^���Ec�ЦW�Tz	U����	��5WZW��j�К�&}���
P꾏��\B�_�w����o}t���V�T�%W������P&��|�㶙L���1_I��;܃(����D�jc���t1�c+2E�h���`m�Q�㭤B�+��
Q�}��f�Ů'Kʢ��������g���9!b�@b{����!���;�LMְ�'d��g���1\0��=��p^�)�E!��nB0X�ֽ��������Q��ī�U&#ϟT&�|ʸidDu?	еۮ�f��8�ǨE4S$4::ϸw��z0�3/x��ѳ\��o���H 2oF���I�$[���S�WG	��v�ͽ-�N�MS�H܊@;�%���C��u��:���ʒ��?��ϕ���?�<�{�?����Zpǹ�=���CK�>�`�/��^��{�"x���Ud�n���hϖܣ\�Lh_�T������_O	��2��1��S�>�L���f���k�����@T,�WpZ��c�*LC��uOΞX�9�M�7v䖩�OY���qa�������]�$}0n}�1�[�N��%���W�%Ao<� ����\����|����L�����j�JM�w.O~���=95��b���GLЀ��5��q�ԉ�da'l�H=���hk+�j�D}��Y�j�1�Lۛz��_ĕؖ��;��e���ƨ~����D(���ā�W��mD//XԄ3jd�.��f֕|&���"�(�-��-��]��3�,4jXJth2��(��9�0"!���ԍ?�����ub� ��`f�w��������n�ݸS�A#�l��t�-�hgtc���c{���,WT!?R9�� sY,��b�Q�}-G���-��T���^���(V,�2Ew�F#�$�R6}�k���G�������bƬ�Ð�Fp�.��X�$�69��@qz�}h�M���VS��ͣ�H��7�I�X�}u?~v��פh4TM��߅Mظ\ۤ����q�r|N������%��t� �iy@�r��B�N&����<vd�ܖ�2�f�˺3�CB/��qG��m3�s]�B��G����ix�Yf����J��!{M�)�H���Qy4�/8� V�s�=%$�bAm��G�/-�z��S/����p���B��I�T<�E,��X�IVN̓w�k�V�	i0�9��o&��/ꫣ��B��c��D��~ &����x۝k�s)�?��o���7�%t��!�0��㖔,���c�1��\d&���GC����W�E��Ȑ�a��ݣQB��B����v��#WX�^=f�h;�����Y�"����g��\S�*�79��3�m��ǩ-6<���s� '��N�/�_�+m�r=�D�۳�J�j�>�x���z��0�)�P	Ov>�`���<-R�r�q�=*���I6Focz#��|[՝$ƍқF����'����m�M�0����u�hf�Dc":!.���c݉M٩DܵX����d�����hE�GEV��L��9�.�0���S���̉"�����l���H��t|��įƫ�s���72[�&t��Ř-��)!{,cӊ���s=����[(s��a��hw�7u�~��hG�k�65��ڽ��٧u�a��YW|��Γ�؝B�m.��I��V0�ia��H4W��8�]����x�z�q��n�ɟ�;&��{�T4ڐ�@(\ �2� ��l��<��P��.N�� �U�OMn�V�{�Q�4�~F��eٳќӇ~��`g���E0�#Yt���;[�zj�%����co���3$9��_2>l���,�b�4^�WI�H�ۙ(���i@���V�s-/�%���
E���4�X�z`��n��r�&vj�_� \���<�<Z�c����w����,/�`��y��П��5)�a�qO�A�mL߾��Q��q��V�s4y{ީ�~ �y�AYE���@|�6�0E s��\n�dBC���o2�)ɑ��Nwp7	�e�q))��L�_�j�y�J|O��(nYg�I3����Վ*�/�S.��#����0*w�Q?�e3��9εB������8m���G�`�D_>���O���L�ۛ�S[�T���{&Y���z�Z�Bf�2�v����fU�Ωa!4á J��ob�أy0'n���-V�=�<���&d<_�t}n:���ο�N�����O#���ҎC�����9�8�9�`䗥���YS�@��՘ED=����u^�
H�D�yzV֗�2G�j �%J�X�F��D9_��6��v���Φ���5� 8��URN�pRe���b� [��4B/#$�5�lNMy����晴>�)+eg��2ۋ��tp��Y�U���Ӏ�����w�BfC��,稌�F��Ȼ��؂ji�2�B�������]ZKf����<�\�D�;�P�Ԉ�w�o���7G1H�;F߭�I���dS���㳛���4u	i�֤f��2����)cS[i���/6����<b��o�ʓ���/R��梛mݙ45� ���z~�2�N�z�ܟ�;��7�2O��KX��^��'�<�f��8�#�F�/Ck��S8}3���0�C��ܛ䎥+��%�3�(y�A��������k,^�'Ј7�!�f/����y�5|,Ǘ��G`�<��&��6�'�3��F��X<!QEn�xn
D�ɚ�gΓr�K�������G��� �(1;���[�3~�vI�V�I<

�.�I�x����Z�~P�(�����������(�E\͈��S��=�D�34�bX�ݺ>�u�{L�S8װx�
���L!7��{��sH{�`ɁS��J#�F]�����1B��c��n�M�(al"���_|P�G���a�kr�!:���/��� ��޶�SR��@'n9�k[�Yl�l=�Q�z��n�fi�E���@�y+�@��Q,����t>�[�YЙJ3���A��	��*�~2�#v�����M�m�*�S�����S��C1nW~l���K��im%�7;�	a��Z��c�Lo��"��L�ƳK5�r�PϺi �����V���ت�;_x���]<��0�.�5�14����P�����q��OOI��P���������w䁖�h��|j�z�B�^�c�K7w��=�4&:���}Y�����"�pY�"�2_jSH�b�_�T[�F��Z�N� ��`=��վ�f�
D��tK�F���(�3��)��
��>QQ�1���1 ?���}*	�� ���D�M  ��S2��fl��t��ڢ3�_յ�ETO�uL����h��/���4��I��k�=߻:+�K�<���2MS��_����ss�WV���ZY<+��x6�uI۪��	�4�G��q]	�{'C"R��Yd����~�4jŶ�̭s�Č�0B��6ɽ2����z�������S�O����>�M����{wo������Q�m^A��f���F�Y1%[k������ti�D���X/�1D��#���D��h��9l)w��H�F���/�L��f�3R=OXΠξ�k�w����:X#.+��H����7K1!h��a__"�l��쾙�J�\X��e�st�딗9f4#��>�7y����Sf�y�bϻ�P�����bd��*`�����˨+l����;�������o�ߖߜ;��F�a�N�ɺP�TK��̤�+Jc�q�)\�J_�~2�ȯ~-��y
�Q�j)u��
�7R��j���j0��M��Z�*H�ՉNdAz!�=���J��ߔڝ���(�ʀ$��V#]�Z�`xә�U>#�d�.ӑ�� �\��Cpi#^���f!>�q@���ؿ��B�s���M�2.!�'>�*�P��O��/\a���V��A ���d#�������v�{M5���7�f�q��Ӓ�htb��gK��>$&-�+C�s�ɛFG� �+�/�V��z{Nً�.P���)x~#}�U�� \iB����GB��@qˉ/�']�@P�D^�u+��K`��=���>n�)O�Z��/�P�Ƿ�L��̷�;��3�$�Y%)W���o7�92�7%[���ٺ�rAF{	ǧ�i���2DM��^�vh����wgۂ�z0G���&^R����9c���*)��r-(VB����sl�V��Fk/+�ŃR��}���]b�/H�>��. Z[����[�>A��>�����z�.��G�T�,ٲ�Rc�����*��nd3i�];�L=�_�X7���h�(����(8ep5���|<��b�Ԍ�eg�'b�\�f���͖�riƕ��7��M%XT��|l��A�^/Pg~U�
v<���(�E�@� ���eA�}�Mv���R�*��h�{����ۄx]�@�*�)c�<$e�x�.��"�Ou;Ś�^�ܮU�
��Q���U1�Ԛ�	�ޙ�l�+wʇk��?0?�}���%h�NS�#"��|�5�VɁM��\R7G�X��ql�<��4o)o4Wܿ�S���ʶ�3'���ޭg����ѡ���*�߻��ۙ�����1���C�Q7I��؟�� ?0(��(�K1?R�������W�hh�좜�ٺ�E�e�}��`�E��D�M��ط��ݮq�t�LJ��?�e~M�Xg��(�;wV��dRX�?3&خ.��&0���po��#[(z�nJ����-Dd!h���h�e���:-���n��SߺK�/� L2�E-l?F�>Q�!C=��}*X;9��8�N��ٹp����a85'ꁓ6��+/�,�?����yV2���@�ɻ��v�o=L�Wh�sԬ�P�99�L��DL=u\����(\@��h����`L��mD��
W���`>��f�h:��{i�d�fY� [t���V�DxB�������/�_��_d	��m�/Ma<���u�E�N�m�ʍ\ę�~c7v��/d{I5��x|���O��f�m��y>��^�r#�	��˸�� m�
�aEWE��u~�:�UY�SR�����"(0aH�{IN��@�7��d;�b."�oI(-{ķq��j��@z\���<�6�����Uku�2��-a>g�2qwjȣ� ����t��:g7ͮ�7���7��E��;�� �Ƹ��rJ2�K%l���ڴ�p�
���h;��O���\�/�9"�<��P�@�>���L�3��>L��}�*T0@���.G�^2�B�*�����F8��s�? ���iF�#��m�ֆ>�?c()0Dh�!'��в���|Z �i�]��5+���#�r�d�d_��
} ���ƠBc1�A��ESP�ϝAl�$
#`����Q�g������e[Z8O�B��B^@Z����N8kWʽa�H�����&a��	52~���l�o�f	�H�r��ofN�=7C�w�:0z$S�(A�`���B��x�ԁ��/}�{at:���R�%�QM{�Cwe�d5I��BfMš�@�s����@�w�S��g���Ƚ|�ϟ��4ʓ�i�R�Z�:@���M���_	b�]�\fc���T��.>oy�t��&y����(�E��BIޟ[0�x�;�^%1�'�����K��V'�p�u���).~�w�f<֒a$�W y;��A�$�!|Ƶ(zkY��cߡf�hɪ��^r�8h�"A3�G�����C�X��7T�fb�7D;�?2e��{�o���t(� �#��U�t�D6��i1V�ÜU�^��ҳZ���Oi��y��.ض��)Z��%�x���ID�u�F��32�~�#J�?�RD-V;B2_���%s�eU�+�����4���++�;�Q��+*��hh���U@�*���?幉7
�a��}�����v�5�����KnH��.�Wˮ��A�����ou�0N��ɗ��<��6�WK*�#�(��!��`�Ar� *_
¬��ezi�f��A՛��Sɩ�&��;��Py�_��<�W���M=n�som	o7VΑ���6�;�8�۝e���`���9z5�E2��*�E-g�@��b�1ȶ����,�tT������N���[a,���ϸ=:_���I8�$�Ә_�Ҥ���*
	����ob����,5���O�CM�?�RV�1J0�k�~7�MF�#���y%��d{�r�Fi=�ej�'�p���[��X�D�Hx��-x;�����ce-H���KF�����^�����~�m���
�Q���^�qy���ΑGo�\r�؝�zw4	�ftX�z8��/����:{�ŅQ�HzXf��d�;J#���� ���6J_�%�2����]�M���^\yi�34y���S�;���9(�0�7�2@6�o,���>ߐ��_cI�� ��LƱ����G"`�f�2(�hU�@���I�V;0[�iʬ��>�.�i�V7��t�i|2&�7���S-�"ǚ_z~�YU�^Z&��2����ի��8G��Ԩ�v�/�&[b/�F7��7����FD��1����`�>�k�$��n�D�R��IlbN4���Ny�B5����b�=2�@�Ϸq�he��{2Q�T��|F@C��^f�sѕ\_a\l�������NV���A�����)Dw�X��t+HH{U&+��(�:��9���>�4�t�K8n�o}�m������[�{V4 !yy��X�tO,�γ���2���4@�;��	�6aog�����qi�{
�9Féy�g��k���ɱn���׏�'��O�������ϏЫ_tÄ�`b�[�3���pX4ZA���^��/ �"Ⱥ�rF��N�j�6�V��pޣ@�l�e�y6/�k:5�*�A6�G��i�Y	�b!3y��.@��@��/�E��r�ن���r�������[�������y��P>^�J0�b��eI�7�߆f��_��7'�%��'��#��FI(y0���fBo�0�NG䄯�yk�t��� ����%�����@�!�9�v�8�"P8����l�-�η �'�c�ԙJΛ��9Aެ'�ϫ;�m�c��)f�����ȴɫQ���d�7�xQ[���*������7M��a��#��vytl��"e�C�*�
�(盇r�qJ0o���d+�1�%�/�J<���M]&�y�}Q���?+1KQ��Gړ T�%M<(��XT��ā�	8Kr� B�@� ��:�-�B��	(Գ�5�,/;|lQ���������bQ�T|�&�R5���j��A�T. �a5��"��h�qg:�69�'�]7�H�&;E�5�H�
F��� 
rc-m@0��	�ɯ�$�v6������k�%��<&�6�DW�������=���ۻ|�ŭT�_a'c��h�5�X�O���)ũC����a���W��O�Dݚ-� �<:���_��Yo��{O|��h����x��������;���J�zq��>�P~<���$ZbI�nՖ�K��ᴂ_�8�d��\O��d�A�!%O�C�K���+ă��b�\�]:T��Y�R^�z�A.�0�3�ULN\��V�?��<A�F���a0jp��j�R
 ���*�H�*y����i,6wK�SI���JL�l��Z�X[h�K�3�럢�$�G˳�ėDK4d�a�TPH�FJ�S��v�����"5\ϒI�kCm�˸�&�J�(>�m���xa��qqq�{�V�v��s�MC@c�"_��=���z�D`�ٜ+32:�����8e�3�ȾT �3���7�e�Y�޹k�%�?�n���x��
�y}����[�� ��U8�P�X;���~Gx^9ׅy�u�;u5]^{@N���LX|�����y�'G�!���kZ�d$k��آ
�Q�7��A�V�M���wy��]X�j��c���a��$I�HF-E(�qy�hle��3Ix�8R���u"`2R�s��#G�f"�������w=ގ&6���?W��MՃ{W<:4f�wZ6-K�J�=��=���p�/��h����ֹ���j�P��N���a�❹��j�irsB���FJ���B���n'!��En��3�/\�^�3Zvl��m{�Be6+�!�(�;�Ժ�5�.H���0;�.,S��>L�3T�*��X1�����Rf��%��T�;�CGy����r��	m~�B?�d��CB5G�[9��3���⪊�1/����JЛ��w�\�4gpd>�b�a��xK�$l�R�#�P!1��h6ڃ���:|O�5p�`�#A9�N ���Z��[�����p3$��2������[{�g��I�Ӡ��j4@>����(*k.|K��E�2ľ�l����g�A�u�7�\�W"Y"��\�.$�!cu8+��#r�*��SzbIO��F%�W�I֔I�܉�ↀc=~�ü�~\BJfX����1�҇��;�d�T���Z*o��#C^�?���&Lh�U���bD�f0\�
ا,/]��P�ʩCiW�i�G��������	4iY����PC�Ҍ�وdâ@%M%������B7�z�<��d�gD6H�;g>��/o©���� d����ƵYa#�q�������r	�Dn�;��D�P_�*�	c=�S�� �c���lJ ���VS��d��Y	���o"7�:�Q"��òP4���2g�]��}ۧ*��r9ne�1^׶�
�T7N�ҏR����k��z޼.�gzB��5�j���~IJB�Y!��*�ɀ�c3�/f��UU�Ԏ�A0c��1�>���=��9&�������K��btG���\.��ݫ4I�Dx�
�W:E�s�R�N�cf�gW�@��b�lG�Y�x����U�}|zq��$���
L�%�%s�������aH�g^u�ՁS��⎆�ٙN���q�T	�M�>�C'���O��t�������Eg�%%�F62�����-�u��m�Q&��`I����O�Η�|S��j����	��؟w��?Ӡ4����N�\խ��"ю��I���{�!�~h:\�ǍZpmhӹ�U �{K?��Z�smC���JqIEє� 1A����X��\+c�u��O�#��u��H(	�YMG�mk1י(b��Λ�&��}����c�7�_92&��μL��[b��I{c��w��`O��s�=#Q&R�&gW��=zE$Cħ�mח����(�ғt���������M Q�T����1�9�F�������?6T&Z`$�	���4��h�U���]~@�n ъ�Q8/�V�Z�5���D��Q7!�^�������P�7n��|y�ҵ��������c�a�8�f`
U�l *�C�؁{[ވ�`�e�\���������_?� [�y��h����G�D0���90�̔̪�=�5����Α�8�sj�|�*�q?�Ƈ����w�9Üٹ\�_Z5��œ8Bʪ�K�9Jւ��c_�7{���&�WU�Ħ1E�W�2x��0���)�aq��k��P��=�qkPZ�e���O������B�T�,v���W��� &h�A��ٞR$���Z��ӹCi[�������΂����~�s�hIx��@��k.r�	�SLt'21�{t��!>A�З4���rԀ�ԋ�$��s!�D<����;��7��g��-!���������6j�?��|�9�]ר�ʙ!��{�V`W�RĲ_"C�P�p�9ȩx�i�g�J(���6��O:O0fܟ�4j��K.O��kw�n�hf#j�qe9��] �������ud���;!8OX�o��i��f��j��δE1"��k�֫	�&V���LESoÊ@��ڗD0�Pۅ<�]��
��!�`?�5R��CKŒ��6���ih}�U+O|���p����)W���(b���_I"M��/65G�_�ӽ�f�}#��}s����Q������濍�nĐ˫j3�.��ؚ��'�Y��ӓ���C�i/��<#�$<9������Drk)���\a#���55��be7?oc�?�qo|5�h%QrAڴ�s����dY��VR�qQ,e�ݖ�B�pl� �S�5S���S���h��]�[�^��&�]EU��%Peȶ4'bly��]��j��y��)S.M���SX��H¯����U�S�.�Vf	���'@?��a�ը�
�@QP��E�� i�~yH���
�%�^&�G������υ��r�V������~w@Lu#��e�8�k���c�1���M��O�]t�d�L��4D���vR�4Tqe�l��ED��ѯ���`��K��(#߇+�F�l�����KL�Ά��es��A%��#ӱ�>���#����gJ+ꤧ��?6ޜC���א�`Z)Ύ��R���F��>����Z�%�.�L'q�1]���A[r�-�,���p$P��ۉ�/^iRG*��:C=�<m���&r��p�`M�c:�ή��g���Kg���;��݇"����惍�ww�x���y���G/�P8v�I�٭=�[�2�do�7=qq�m�t2��yfu���h13�48��-};0���2u����xw�צ#�R0a����.tV���Lx�o��`�/#�K!���%�=$7�e&�9�����,nf!����`{�z'�Etm�Ƅ���۵D��[�O�7�!�k�]_�M��B��}oI�����3��a/������6͋����g�ֲ�a:�C<�����/�nB�v�s�24�)���!|b9O�'	1����Y��/�QȦJ��/��w�¸�EDFLu$�#g����5�Vs[` <��y�<l���8j�4&u��b@�$C��r�H\d�C6�'7��#V٦=I��A����m`��ݍh#)�:�E�������&��C�8Bv|a��P���x� HP8ˮ��Mk�� ��PTˏ}�?�]Adb�σP������Q��&�HY�R�a���r|W�Zc���y%�L��S�^^��C�֪�P���@���r�vբ�P�����P!S2U4aگ;ȼݺf��Y��鴛4�̥ϖ�8�{��e�
X��2��}�tp�D�U�E�J	Ը���������%����ܼ�Ž��X+� N��E.-w�lDH�	��^eb�n�HN��Pn˟����5VKy֡/�D��s#��%�7a4�?nv�T$=��QmUM�w�>����%K�~���t7+���I����X�8&%��\R�ԝi�*���+P3`���_�%� A�n��2g7d2k�}�����Uh!A�����}E�E��E�=�"��)4uj�0�28�e7z��^|�G�@&�j�7�Z4�.}�*?�<،�	� Lٌ�fl�Gb����"��M5<1����\�$D+��8ʶ�W�P�]J��@34�z���
'�x>�U	O���r��+z�\��pT��O!�F�3O{�-ʸ��^��aB�{.a�mǯ�+����ՠ�����X�t���&�+U���`��9A�J�+a�V�wB�W�@u�}v�If/sD{NLю2��K�z�8�����Q"�c�ӌPs��G�^�I|is�k��K�iG �@�_���"��coDN��%%-d�^7M�`h�d���m.x~�S���2��;紤z-��?��������wk��vxR�r�9[�v�EfTxE$(H=�|��Sgtd]�)��2ڒi	�I��/d�E�l��T,�٨��v�L�Y���FQw�4$��Y�m���6�m��lN�K���p�����ܓu/�].����Ao%4�֑��긬S\�Bs�K;��5(�i�	2�Gi�S2�I�3��\���$�dS[���T+��ʣ�ȏ���omU����R`��k��n/�aG�v�6��(U����[Sӡ>PY^�վ���e��ŀ�`g �y�?培R��VJ��4c���L�8U�3��HO��K�GSjjS&�ǎfH�.�ɝ����i��p��
L�3�L�&CO,�����@�1���H��؝��s���T[���c��]C6��Q	/o>ӹ����#���i<����q{2��܈K3:j����e��4Rr��V��ε{py݄��q�Q7����_���d�k�j�Z�@�.�I{C�mX��gY���l �ഡa˽� -�8�}H�Z�mᣞpb<�I� �^_jV�i���	�g]d���۾,D4����k���0q��Rj:�I�c!�0e���fы*�"�n�kؙ��o�+U5+H�cL�.�UAΐ���s��7�5Ҝ%J�3��=�*S���h�;� �+�m��T�,�H(WʞN�Og��No04�~`����3{Y6���I:{�Ό� o�y-#��W�"�S�k^����o�f5��`��C����2'�׈�>��;�"Yp�N���A��3�;-/j��vk�D�%�cڤ�C8R�D(��Y��dz��0og��{9'(l��Q�4�n��v�W����=��blMl�"r����U�=C5��e&Rc���Xf�*��]��A����Rt� �����p����m�Cm��-�y���e6�G�h
/|	�+����8���h�����:*�WQ�B�3������8R�$[Uf�܏''JDBιI)#AP�v �K^p�+�D�4p��r��V�n�I��j�!c���SU�g�x.��N�p6���M7��u�eѓ��Oh<��L�}VE�'�2�q����RZ����4?��с�j�����{U���/��?!W������_�^w�'Q�X�5NfV�f�/M�r۶�0ь|�|�$�k��@�>��E����!u��L8]yF�F����� [�F��X����Z�O�
0wn���s��뵂N�����^���FqO&��f�2��;Y�?�(r��/Ń�����v�Z2s^����C����+{m���������="��a/��n"a�ԙ�ܞª���DLv��~j�GKu#Ѱ ���>��e��-.�.�3R�D�g,8Y`���x�Pd@��u��W��^��/�K�`xP_)
�a>��rBр�6��>�01Ȅ�в*Q�:�Z0	H·�E=5RS�
�&񹆕|���$��#���uFj�R�Q��ȴ�/��B�5�=r������Ȭ1$�{$8��X�eՄQL@ Ω�1��]	��wۯA�G�OM����(T�˾��?(*�� �2R|�\�ڷ}~IL	T�
�6{{l�-�1�P1�A$��D-G)>��(��B����`����lX{�����OR��&'���"2�Tt����>n�wOqj��?�4�Yd=����j�ǝH哞�j/_xPī7��¢s'zi\=m��[��&}f�x�km!�ˑ<R�!�0w�x.�x�V�ws:�HƂ�¡��U�𚀫΍�-�Y��͓��&	%�`�K�xM% �do���w��I?X��z�tb(�)8xB�s���;{(u~A�8�^�)7���BiaAH�UO�`O�q`�j�?xn�J ��2�ZcH����{y��N`gY|��O��o L:���آ�A���33���͎HJ����j�q@���1S��SE�񦬒ݶ-Q�땰I�P\��q���Ë^��܇ �(�Rz|K�i,E�f����W����@<#wj_�ֈ2E�
�80�/�;~%���(�c�L�'Px��o<6�P��j��!}��[8�ʾi.|�����A-G��'��!̙�Wz����[��Φ���"�?��O�t��_*�A�a�U����ʒ��Dtv�%��	�F7o�ԏ��!i5�W
�ᐰ����y�@��b��Y�n������@+�����(��#hZ�gO�����d]�� ��QZ.�]�4�L?�G?�����7"�Q��S��� W�۳��Sm��7���6X����I��څ\w���'u��h�oh�;��"���������?|�r�ú00H�;�H�!��z\�;1i�%��Oe/I��#���ߪa�~��n����C˽~�ړ�u�X����䎃�S�;���ϥ�҆��V$9��ҭxa�I[Xt����Gj�_O���J����]Q���v٬�eT˔�S��	M��v*g��#����|��ƸS�=�@G�Ut���5<+�2!�rU��C3����Ӳ�6N�CG�XS�W�ES�M�=º �[s��2*���dsq�Z5��t?��������u���g�D�o��2�V�$& *�G��X���K'>BN����BaN���B �grXk��W�"5�:��\7�s��Js[��`S��
閫��Y�D9��D3g�ݏ��ZLQ&L��TM�(�1;0���G�aeҮ����	I��4��GBmt�^N����jy0�6�d�a��z�e�i�V� ���*�8L՞���pɱH%Ib�*	�R)}�q�d�"�b���~%a������a�r=l.�M*�s�3��%L�m�B�*eW��HC�^,����*Ү���_��$�t��u����2ƃ�E�x�)�"̟x{o�r-nv�Y��y�B9;7�n.*�"����a���qY`J�}M^�\M\o`���ȁ$�����iP������4	���0��	ݩiv�bd�Qbɇ�ɒ���Yߦ:�Y9�9�e�5�n9�ɝ"�Nr��u��N僶��x]3�-�׵��3X������uA�c�"�UTg�Zhe��n�ԧσ���Wv� D��M�g�ϳ�'Q8�}� lux�?'O���r�y:�1Ԏa�Vh�UM��'&�2a�/��v�b�j�`��c�I(k�������]����\z3*��#�I,��.�RQ;>�����]�og�k�K!Ud�.���d�$$�N{�r7o��'!:�/�,DC4�v�I-��%�?�䐺h�;H2���X-}���_}I�Q��*`,̓ufg���9olT�l<�$>�YH��J!7�<�m�Bg Ƣ9y��,3���#"�c/^i���O���:��%���o�OyɊYBߝ����e���K�����I�R���DƏ��\����I��i�h.�\��}y�f%.��J��t]�{��62�=�O���R�ñr��x�>��B̴45H-�u��<�Y#�s)	Ȱ���{��Y���|}��C��-�ߪ¾)�
�7�6[�#_�2
��P�L������
&0L5����h�d6�Yst�-S�a�X�d"mIb�_i�@��8?K���30�,��=^��,�Y�L$p� �C)��*=
�VC��8~�"�銷+�������;a����=�(O�����f(Wد�><L�ى�� �*ޭ<��WәMt޸*�
4������}�v�!N`�-{�)Z�K/]�}�k�F���n�b(6�Md���w��^<��UTf���v� ʛV�+��]\��o(�e�/����(�͌�nʏv�碑��G��������K��."	֊86�h��ɪ�Ab�˿�,?�J�G"+�G3A��T��*at	������;�,��V밝��f�S�I\?E�H��[��O���~�^��>"Җ���m3m��7�r��E��"��E��?w�b}����a�n��o4���K��o4x�p7<�I���e2�@���+����%��+��һ��k��XЏ�����(��b��>�V�������!��~V]ʠ�oQ���� ��wip�x~��>��N8�D�=�@��_Sʫ�]�^	,� ��3���_ܬ��jt�;��~dv�=��ɍu�d#���Mg�I��q-#I[Xɕ�j1$���u�O������%�B�𗲉(��iQǥq��-A��<tD��"l���\�A� ��?�HFTL�(��!K�b�,D?ć�f��,!�{�gv���0��/!���k��*�ߖT��WΌ��e�Ϻ+��v~�"��..�#xJ7�FW�l�k^|<Y��{�<�%Qk�7yP�h�����.7�]��AG�R��磅�<�N��]^bI�`0OE�n��d�^1�:�A��ԛރ��z����ԒN����H::�a��bR�c�ѡ( ��1#E-�Tnv�c�Rf��_���D�(Bf��%
�g��JuO�G�t���yPK��@�>f���B:�;S��J�d+�5~\S��d:^�ld8�/�o�)|���.F�N�5T�͐{g5��}��'�-y��_g<�Q+g85����lvP�`���T���������癒��V��8?�X���R���ʿj���f�}d��+��O#ϣ�˟�F����VL�8��8�w���+#q�c��;�/��<�8�i�%�r4���E�h8��N�㤁��z��(.��D�����_���T�1\�+4���E�?m��pw`'J�.�!�'^�x����}Sʹ��drk6Nw-�u;$�fB��h��`��bR��L�5^0K���}�<����{�����A�>�\yf�1Ji��$Cp��)�f���0L�I���p�.nC��S�Y� ��s��r��]��\��E���$�k�x��`����n��[^�Z�8��ϟ���\�#�6�����r���N��s���ӟjG��A�T��#����BٚX7@���M�ڳ��2s��-����LT�՟�������{�̸���z��#��Qx�yѡkO���0_W��v�	�|Y�i
}M�����ܢ�����<Ƨ#��ఓ���k���T��M���E�
*Ϲ=�eɝK�f�D��<����Oc+z+�^�\����7r�_���M]����iM'����c���c��*`Ţ�:�`_ڡ����@	*��Z����:��n�&�E��Dg�2=��x!�ҜL���SpV�s��<k>M���������i�;�x*FDs��~J�����"��eߴ�yM{yU����jd�0��LU��t�NU������V�XH-���Nl����#�M�ez]Zz�e�Փ:���'��m/;g��mǻ����U@�"�֍�KL p���v���")Z�X22�.sZ��hQ�ʊ��s�`���nDU�	H�b!���`ͱm����KbQy5[ug�h�����l�;���5�	!81���eo��9�͵x˰5�B�vtx]�X$�]�3 D�q�Ӓ� �Vm[o��{�1�<}Y����kJ��N���*�A
48��'0����]8oo���2���jg�J�ޏ����e�WZ^`z�eR7#�` �Mh&��À��g5�)�oێ����s��&�.Z?B�8�W���Z������G�	K�
j��M/�Ak��߼�),���ժ$��:;�0�HI��5�4� d�G�E��w5���@�!�D3Z�j�6by�8|߱_FyPL|QE-b�3o��/W����m1.��ƍiO⟌u�6�A�J5�JsWgo�/.�W
5�c�&��n���᝽�5.O[1�J[��xߕ-�$�V��ogA>s�8���*��X�R�� �=x/q�[�㱘(*�Zm\����@� 'T��yo/�4���=���hE}�g�]'�!3j���5zE�����Db��4t郚�r��JA��.#{?�ƿ�Y����g�8����]LHƻܻ+�֫Û�vX����H��j�u�:�+).I*S�G�~R	~)�����Z�����W�l�K�������y��0��=��
�<9�D� �ZY�V��t3��g���:vQ�kH�I�l��Ko�k��M�������q�:u��?V���[�䙻�J �F�7hg�q6��̌4��7(װZ�$>������R�_�Aü�/6���@η��ìF�d�&�v�G8x	�U��a�m�\v�NN:;;q�W�߬��I-�����Y�~����tm����
����H���)Ma���z���+�fG2�s���M2IZ�!-n}�l�L�Q)����I�*#���ʈ�@�4S�yHج��_׸�G�E#B�4��w�Eɰ�l3J����N��캄5+�u�ޖ|�bi_D �̴Ǻ���ͯ��.w�V>{�5@exo�/�o{��$eǨ�:u��Dl����)T�s���p�I��Q�}�k��~V���5*w&����S~�Ʊ"� �삼��ҊX�7���L����ۋ�����GUi�cx�u�����U ����ͬ�#}�]K[a�&�ǁd٘b�J��/w�'|�GI��x�;�ˍЇb��W��� ?Ȃ��F�p-���XH���,zy;d,Ɂ��p��-�%NW���5A�$�/nl�l'�h`b�\$��n�}n��t ��ah���߂�X���v��˦/n8x;�n�4x�T�c#8���oM�����ɲ$I�NLa������ڇ��hЯ3	h��-Eߴ�N?�t�������I�O��a���C��d�\���A6�b���˰�?3]�͵�����V���	֚� ��g�D~|đEC�����ڑ�n��*���Q�4����(u��Π�m$����t�~�O��9�f=�b��FD������H|���	�õ��w)��J�)�����l��.9�K`��"55"�Ƌ\��vh3��,r����U����#���kq����7!����	RI���&6���z�$��/S�WK��"H
~�\J����z㳭Bז���J��+��"���
���E�=���Ԟ�L<�3�9z��ߗǫ�u`��bf���	7,j*��B��:�BӜ	E(���N��*'����(4vڌ�6�=镀^��(J;�r�6�W)���A/4Kۺ�֮Rc�`}����d����C{�r�ijj���{��E�+��f������|p�]2��Ө����$"p%��MX�k8�fӔ�A�[qLzC2� � 9泯�8Kn��\��X�!q����4$��DЅFp��ӆ<�Q�����@�=���g��$-���}j�F��\~�~+�&�յ�BN��P|�^k�-B���QAG���+`��9���te!C�g�7��B/g�Ń��y�dBY�Y�`�i�
�`�򅲤��n_[�$�7_`�a|��#�����.�S���g�P1���	8
�����@�� ��mO���"i��^�H�A㖔n�Y1���g!謳���N����du*&��>� 	��9hH-����(�yv�ƛ�9~:��sb� ��s�N	�2���J���^�МP�ԅ��[2Gho�D��/vcm����K���$%�ؖ�f��(đØ��� ����I�)����uA\��G���J�Pʠ�!Ӛ�2-Ǿ-|��)K5�K}rC@���U?YAJ
O�k�t�W@4K��Cl�Č51Ö^f��m��k�qD�n� �-&oʜz��ڛ�B�0dp�g��8c��F��EU6� b�K�XC�{����'P���c�?�bT��SC�0٩2�88t�x����EP�#H4�3\�9EO��,�B�ꙅzE�	Q��\鷾0@D��������Wn�n�鴷����^}�$��G�q�WVႣ
+��X���7��Lj�}4�z��Z��Ɵ~�߳9|��[����h��(�E�8u�Bp%;��&�j`	��7���VA���񏶔\�r��]������G�A����,z��-gѸ����4k)��4�J�!%���綰g^C���<�t�9�A[����A��W�.LVw����\k�i&0�9](.�*�t���f�j�|�B�6��)o������W`vtؠ��� HwemxͶh�M�t�ǫX @{���(�n�E�m	����9�. ����ڔ;xi���l3s�{����
��&B�Fv'�3F����9�h
�K��<�hw����>�ŮG�f9��֯c�-J�wB�&Y�����lr�5����V���P�Q�}����ʾ������2�-�"�C<� �z"���d��St�_c���8\��Ps%�D�)��J�֌#�d�)G{�J�v! G<�J�(���$�Zd?|ϿQ���r ����~2~���H�V���"�A���n[Y�)���d�Ώ�c�n0��e���F�A��h����� ��j�.w��?��*��o���)pB�*��9Z����|J	x�ᶲ�z(>�K��b=���,Ʀ�h +��)j�S� ����]��e�F����`i�u'���~)�C������+En���r��E'	n�*��q4�T�T����udU�ii����$_�w��R��i�:����L��5d���d�*i�x�ƹ����3���)#Y�� �I������OJq���ݩ�g�wO�������kQޜ:d
����$	M��%��~� @퓲���sX5gMB�����I� `��Řd�3q�	�uz�O���S�ؒ����  䱲� �i�,�?�����|�Fᔅ��G �Wc�c:�>�jd�!~^ق���AA]@J��ˢDŏk��QS�}�V�̊��}�ā���y�N4R��+Z�۲$6K#�Yh~U.�-D�`&B��r��r�KsD���:i=��t�[��L�x����<]"��W�'�=� lP�6��p�!���_�'1�K`���5܁�3U��Ζ�xPf�����'�I[��e���wYM-[�S����T��paA4_���WC�v����$� �鏇�Ч�(�N9���-YՋ∤ᣨ>(	Z
��aǮ�M7J ��W�h�aQ�T��|�&l�LV`���n��i��fs%Q�oF�#S��������	R���\xE�@�@�i�ľÄ,�^$�T"u�%��̩~���������5�cWuJ"��ۿ�>�XS��@��!�\o֐w���D�G�B���$�
�"Y*�yYƣ9ꪗ�!�՜$27�}�V3��Hq��I#>\�k�"����t�x@hVd$N�!��� iY�u�#���=��$��F=�J��6��
�J�� }��Qq��s
�p?:��q�#�:���^�����O�`���8�j�e�âO�3ɝG��A}�&[t�<w�)t�I���Xc:�.6�7$���ޟ,�M'��'�d��\�:�<��Ȍ'�P���jS�����2����F:7���7���S��c�ˡ�?��x�@�}��
�ۉ_�3?�"���T
y����5�fA�Ka]�� ���P�k�>u-O�pq�2�dS�sĤ��'JaP��9��Ê�H�ݲ!�Q��mx��:��|��HOmI��
*�^�<Je�Ž��_=gW�R����u���q�:�:ϯ�'}��0��fmf���t�����Z�Et$��mY��'���V��� =cmH�ޤ���~�T�/����>7���ta��<2X�ݬ�v����II@���#�����"��������=���Z��jh���M ����Glۿ>�l���?<u�kX�N���Y{�;�%22�fd�㲥�"���	%��{����P�%#��>�\+�T�^5�b����ǯ��C�E��2BѳQ�𸺉I�H1y`�`1٠@�1���3^H|�����&'�D������&�"3��������J�K�?M\9�#��B���oیDL�o�"w`b����P@+u�3B��!2;�j�L-�]$Y}
�
H�T��������eƪd��[٠1�A��"?^�F:��Q,�a�W#�j�.]��Nby,g�U�w���@�;��fYB�$�����X�r��#m�_��@s崢����A�D�'�*���9�B�]d��Sn���F���UH�5Q�T�wP�r�P�3`���m�>�|�ܱʮq`w�1˘��ZH ��J�y����w}�x:��p�7����Bh�����
%�[��*F���׻�9ZA�Sۘ1YRV���I�l9ɡ%�¡vB�,����
��N����8��\��̤9l�Zt2��p�ڰS��A�SF-a�N���F)�#�LΥ�b$z�G���Y�r�x��ʫ�K�����;�|���|Y�0 �ׂ���prG`�X��W�����$�&=�1m��N�p1�U�уmy
�Lj�0n�x�I��cӿ\�t5���n邴�'+[׻�.b�S���7��ؖ���:C>��h�R��=!O���$���M��n���K"u�$[јq3��q�b\ܧiL;��b�J�m�z���H��ɽzV��bY-I��Xh��y���b&�L8�w׊��4�6�����ش@�$E'��ဴ�Q�c3U�$�ص��O��XC��#o�=���"ިY��g7�n�K���W��*+��0�-W�a#�*��%��ּ�-��󬕞@�;��9~���p+�J6�֜����~�R�`µX����f�����W����E�_�YM�t�E�W�:���&~��=�4�tf�yU�l��Y_�FM��0�7�P�U_��Zm�����k���)/�)��X�S/f6{� ���@Y��W�}W5��ǟOp���x`T��h�E�Fni���8���|BA��0�!��{A]a\����ߨ˓�)�:]�^�&��Ӷ�;z�8�����#��b�+�};��(p�6E@�7	a�DJoO�U=��G ��2���I%މ)C�>��&����X4�hQ���}��f�Q��I�[)��BƄ�G���:(>6
cE˼�S���m�~�����i_�4��h������c���}��H�om�u�N�΄���
�|��5(J*�гk�G���uKK�[�	I��W�p2#����p��F�%�b>��2Ę_N����eH|�A]���l�W$fVA��+������\��bA�+�B�'*���wd�EX�E�� w��w	�|�����Y�'�C9{�?�p쫏� `���RG�U�Ful�I�t|�#z�貈-��c�g�H4�݁&U#g�ږFc!���L��3JG�.���Q$��1u�'�u��a��RUH2�A�ZeE��7e, :a$9�5Mq[N�����|=n�+���i�P_���K���lF�OUm�C���{"Ի�s�B2W�P��k��L���a�~��v`�`�rҩ�l1@0���.�߈�9�� ��cx&*ژC 1�P̈́�3�V8��Ћ��mN��c];p�pu��v�����9"�zo/�Yb7f����Y��.����k�[�:�>���	�0��՗��y;W~yCѼO�
���7�`�md��M ���V������~6��X�y�2���&'8�05�O})�A��@h�k���f/P�͙O2�U���&n���Rh"��q�RM�2��`�����`DH��)Wy�*�J�r�)OF^jv�������X���F���#�l�m�{����t(�8V	b�S&�""�(�SB�QY���f��YEσ2V��6@�@��NnC�&I�����K#оh�t��*`���,٤����:Z�&�}��D�`�K5���r���+�U"�l��_�)0Y,����1H
��Y�DpQa[��������%	XԊUKk����������yUǔ��ʲ7�S�AE�}!0_�o$��4��o/ⴄi�` K��p%9>�0+�שDIX��a>���/O�[���a@<EAm�6�,�5�f�&�w�ˢvlv&�/{(����4G�Hj�`�>�#,b/d%�2�#�HS^_r�B����Z�Z�Q���L��E�%��&B��C�c;;3����e:�LR�Ҋ�=�b�}�����VN [�P���:q�r�PP��շ
�}��R�Ca��L���(�R#b-�G�`0�KR��Ѷ��N_3J��MS�Q��N_��*h�W�����b�f�f�.��у�����k Yf�P�OT�b�25���*�Ϥ�/�17ۄl}W]�����>�0�慎f}�]1R�@�

�z6YM�u��~e�n���Y��*k8BJ�����r��m
X����\ҚJw�p�� �&sx f���
�2}�߄��J�&,�V�L�Y�@�z	22��x���Z608���LVCw�W��%��əXe��0��#M��61sL<�� ����mC俸��6 Uc|�÷t�n��<dd4��%?hn�2���.��U<YԖ%`޵���z���l�ᄔ@�*�u���Q
��QqF �����9=%��B��fg����|��dJ�������&�i<;ʏ0.�tZyK� �#D���}H�����c�<j�T��h��V1�@ ����d���N���_>�^��&�w������[�Il�)XPpݓ>�PmＬ� �d����Q��� %�=zL:�}{YU�UV�qNp�0υS���a���3��J��n��W{H�շ�B!�/�K��Nmzp
��c�����8=�y�P��m��<��V�A�{v�w�֜�rU��e��r���6�����Ct�z����[ ��/�iL���UO�u%����#��Ui�Oiu�;2�&��H�hc�������pY��8����i�tBĽW�r��Y]?�'D$h!��[��0��q�Ck�#b�W�;���i���<�c�7��ID2�Ș��!LXv��NDC� ����OUkW"ےrQ�3�/���vJ��������]@�`Gp���5Wu]��^ffPl��{�;#�%��R����(�ç+���.#���WGI�������@���0I$>�ᵂs�r��ބ�8xN�	*� �1�Q̺Y��hv뢄E��y'P�+�w�l��9؛�]uZ��EC��8��Kb���JѢV5�t����Ŧ� d}����ؔOdX�B�=����GлWɰ�rk&�H �����d\؁m�4d��>�5e��񖔧���GƬ�����3mXӃ�f��Ş��d�������v
=�
Χ0@�fP�|"����(#���'��A�]�q��e�|�5���ø�h�J��>��.'Y�t��P�@A������W�}O=�G /�C�zIđX�9	�!4�&�v��8 )U�'A��a���,\ ӸVV�G��O��~:Q>⹽n[	�V��EHaɥ��y�=5��p��w��7s6�����s�Ȉ=\Q6Y���V0�AKt<����~����{�V�����Y@>����2�J���kU�p�7�����pG$���?�&�eh@���Fz�1��m�Yq0.d[p~Ϡ�7�������vfYq��N��!�;F�Y�F�1Nl��a?]/��d��OV��bK]���E�%�&0�/]~�x�3�O��k������K$�?�����Z�fʩQ��#윫��2�e˟ J��	�x����s�g���3Fp1.P�]j����C�E������f��!��:o#'���ˢ�ۅ(�`�����5�*a�2~�����m�����!ԃ�����u;�f�ܒ��8"S븯
����L��3(#ާ��Ն�����s{�����"�g�!O��z/(U}�I&��3����$M�xm�pȰH��j�1�����c$
x[ZW�����#H�b�rp��	Y���kE��f��ms�A�c�گ�����ޘ��m��Q����b��ST��R��nQ%D�7>5��։��Յ�9��XD�]t��H�R7'F�����B�5q1��z����?��n;^���*uED=F3�̪��h���r)0�1t  ����et�"�0����کs��f��{/f�DR8���u���;���\���C;:Dx�#�#��}���ނ������W�`[�rT�K��K�u�+F�Sհ�Uj��SJU06C�u�N� y�-�d-�������{@m����K 1����1$�G�!�j]�+�
~T;�0V�m��P��6jn,�!=�¦� +@�T3�5�Ckrd@��'�ԁ��W&�zF}hYH�Ȼ|)����"� �c]:�O��&jO��*�Da�sA���a�����	�6l��f�|��8*�f���Ǟ�hro��G������ʦ�Q�����i�X.���iu7L4nt�H�%s������3���Z��'������q5��1��5��Ӹ<cf��%��v��d2�z��pW�|5�C:_k�8���@�p	c�=+����'}T��-q��.�:�@^�SC�+zXF��3�x�d��O)asq���w�b�g��o��p�z��h�Ad|Ues����^�\��72YDC�p��*�+��;Z=�t���-�G`��-�)��/��݉� �m�W�U֧H}��1 �dL�5���G��	���wT�QS�!*�IH��̔=zzx����{V˰��\uj��|��9}�<5�ۘ�U]�_���S�v�woas�W�x!C)85V�B>�xN
c^�q��&.��<��jgӕ�̵�؎���x_$~N�q�uJ0�)�T�*B��Rs����d�ԾO�*��X
�������v����-���!�%�[��:�q���P&E��C�f]*���h�����-75�>;V�Ml	�Bz����B��cF"rMm`�O/������n>�������Ģ�2Wį�n#��#n�qA]������yҶ�=�/���}���?�(Y#u�ȺW;�O���;�t������]xZ�E����DN����,Vc��JKl�"?���l.�]lX�%(�»�̲��W�
�n����pgg���_(dZ��f�Ջ �,L�&�/�<��5ԉ_[����*.����Dc=�ьIkS�����}�0�}�//L��L!Y�Eo�O:a�W[E[&ꂇ�cO��p�wsdS@g�xD���+����f)~��օ�w�v���w�.[<�ր���F�v�ߧS�N�U
{�U�/�eK��թ�;9ޜ��qz
�f���oGE��	򷋊p�J}�����|��]��Μ�2�z�0"M�\٧����qv�\J��B��~�&�a�2p�u6�L��^��(r5?K\$�EbZRW1�2�#ψQ˱fN��T�8���,b�S&�W*���t���� |�'x����C��g&�� �Z�*=Gi �f�n�G�}{���?������[3��"���r,-���oE^���L4{���r���ﳘ6ZF�c�r���^_:�8*:@JS
Tr�C��46+�.��\��В������u�������/ ¾�> ��oZoo�6Xd��(�/vpfH,{8c(�������ވK�bjt����[�Z]��#y��%Y"�-UQ��n4�bS�S�5/"Hf�Jݱ,��N�>8���i�[8]��Ұ$ى3C2��Y�(�"n#r�I ��F��4Z�4n�!LT���X����#|MW���t~0��j�r`-��WMR%�����Kg��ȗ�x��L:�&�Nr�%R3�K�&;|bE������]e+�QM�_S�U�C"چ��ch�Oߣ��[r�dI��k���{�R�p��n�]��#k�u��|i��jI�:*�`s��v�mW�6,��+6尩��WK���S��>����"K�_K39-�J�&�	|3>m��F�����)����a���_����xK�3�j��|O�o�� �����{�x-��6˧��YIշ��0׮+���ScR�w��zmvL�6��W�!�Ř�������+"���~ Wg��-�B� ��g}7GIQT�$��ھ�s\d 
�.���|8�{v� �Ν��z!�@���a$����ך���q��p}�x�����J3	+�㗸*���Xk1|&ة���a�00�t��v#�@vpm�c���2�9����Mn0�/Ŋƈ����)�o�|"ٵ*Zdc ,�\~~�ХG�'s�b��f����[h%��ju���I��aY�I��4Dy����+�M���0��3� w+􆴮�j2�vkA6ّ�\�:yR��@�U�Y�~W��
��XL�v��I�j:YQ��)m�/����O�ړ�m�����p�����_�����U��.|>�Ǻ��a��a�j0�P�O�ӭ����L^n[�<��dj���F��miE;qMf���V�A6��ݐ��9����=�u.��JFȫz�MGpj���#R�W�;p��<��a�o]�����P�E���EU=�φ��ezc� �1i	���="~�/XGG�I*�qQ�����&�x��\�.�):�S`�p�?�ś�G��@Ll�a��(��m���ُ��o��Y��~����E<�z7LoLx�u�唻AE�v@BQ�s���æ����n4�����O�6�NR��n6�GO5}׹�U�m8#�KHF�Bl?D�.�̝K](q����;�j0D}fT~�Ҧ��cpߤ`�YM
wp�����ҿ�\�{��>���Is�vg�b�ȫ�$;�6������R@�1����1�@��Y)X+����7tZ0��#�) a�������]N��tш��ÑK�p�[M)%�C�e�� #}<�I�X�R�\�>���U�����Pfy@ʜ+�+�|�=�⯀���pR N�<�M��s�\�?�����o���������L�@_W	m7��\�Do6�1#��%w� jM<P�]��7<��E�m����5<[����N�Fۖ_N��ܬ8U6T��:��<��C\^^}j�c���5@l� eqŪ%�@�n���3l�R%C���V�J���E��?��߁2��~0 Q�M���� ���FԒ�N���nUJwicJFȋs$������M��b\�V�g�f"�����H�8ƺ]�H�b���*'�KP�8M���r���0o턻�W��5��p���Vm�0�*Hƚ�%�sh�����-ޭ��5ڒ_�ߢ}F*�nr�Z�[԰�&Y����[�L�0]�,�]P�S�em4���u􍱦��@�Ny��k���hΤ�M�O��5���$$m��e�3��گ{�R�;V�
��<�t]� !��`�2�6���G�(;c��r�Ye�"%�O��)�l�����sƫ��\>m,�W/�#���.�5}Em�v���꠹
**�tУX���tv��|�7�,������^�<��W��f#�+ˌ�N��	���M⬥L�ز�H���S3[���z!P�k��#I�Α��EG<�4h�ᾊ78?l��ΰV��y?��x@a2���`�~5&җ�]7�"���ssj��q�"*(i$(;���/����k��T:p������@��2sV�a�T"���G���zѪ���j�EXt]�D��q�6"_�h���_R���3�N|��Y��:���S���#��'����焦1��`vr3!�7�ݟ{��m0?j��%�b���|���> &�q �X��&X��%$��=Sa�m���O<�K�-�p�u�����P]AkY�/!i1o���㒈E���ۙ2�D��i�h��?�KG�s����e�ޓ��VC����3��2)��p�- ���bҹl+�m[5�4	QN���jF�ͮ�g�j�J���،D����5�22t4�/w�$'�!�ә1]#y�Zwm�f��=�X�\˲�naU�8�N!��l5Yg�wf�� ��A��XK�G	a�F��i�0�Z?0z�uEf��O�9P�Ň�C�7̙���vZ���bY�����4�p�Ru�n�R:�e���0�GX����͒�Y�"7T/&��8�js�1�N�q��x�k��SZ�![P����Ev͑�'oBN�!��`e�`@������������_����1����̽�z®�(��P�*	����3hs�n���e2u ��Y�-��{�G�)Z����%5���&�.�E	vg��y��J 7f:�n e_ ���Ž��O��;m�u�Ҵ9f�<��I2�3�G� c��� m����2KOI�f������Ϊǖ�A����`�4�t����)M��R Z!��=e��s�v@����I�iF�E_����4%���]���<oI�&{�@�� �����q�氄F����k-��Y��5ݔ-��K�n�x�-��&%�mc��To�v���IT#΅rvʯ��a�:��o��p��m���$N��6[����5� ;8�yWQ2T"��4H��dҁ=�m�ܢ7,n?2��	f�l�d����f�ޫh:�yRL���Ϛ�`#�Yb$�zd��f�g/�X�G��V&�E��Y�р�/��+�sA�->P_mk���)��I�ԍ$�3�;�Xu.�zL�'��V�����y2��τp��aw�./��j��ѹx�(��6�x��)F�� GLL}<�|��G
��&$�Sۘ���Q� U,-���!�Ӹ�gIHE�Θ^�"��R�݊d)vӬ$c��V�Pdf���_�"��(xt��]ۋ;^U u' ��W�
�;��#4[�ijM��j>k�2�z91�5�z�9����Ӫ9��T�����XӉ"$D� U:��'�����q��oV�z���$�9�g�lg'D��%���g�����~���6'�(}j^�#��^S2T�Y�U�"M��,�P�yo�G��3��o'o���zP{�� �\�A�f�ɔMV�!�1��ŵ�}"W�@NTrY^r�t-ү,Mٴ�)]���ڭ1�'��6'��PZ��
\�N���Y�:���η��9�1�� �J���;n� ����wf�t��FS�'�j��O��3������UkV𗯭��C��}ݲ����s�ܾ�k^  ,�u݋�����_��6�=��_�ڊ�~�I�]'$(D"�Ҙ-s��n���6L����jkUg>�fD��D�!̥�����&��� ������h�e-{?m~m9��W�Fwq"T=~%P2��EBri+�%�?c@�RY�Wk��G�ސڹ�~h�cU-A���&�?OQ ����ӕ�,̆ߐ3�  ��Y!˿"X:ڝ`��
�uDL�s��?xʅ�q4TxU��ĳic�����������+�J��l����+t~8^P_�~�do��u��[�M:�X���e=�g���`�PE[|p�#��s�e�.]�y����D�{���o0���=�5F5y=��3�f��r��-x(zY��v��P����j����;J�����W��W9�i�1Ff����`~C�c����n�:�uF�16E����Q:���:��RBOQ�U��޽�a%=CX��i'�������[�U%^�_8���@��X�;�� ��Pz�ya�/��/	A��- '�Ek��{[�����!FZ�h-��׻�X�	g����ЦOxO�.)���#_��K����UF�({d ����*�U���;���<d~E1��':��3�7��5SG�&]�X8
�P�5G��L�Xǹ���췝�φ.�9�v�N����@Vw���2v���o�$��ʠMi[��V+ے/��!��8�:�׬���H���3U5H4e\X�x�"��p)Ṳ'q��=Zi_��C� 3�v�g��S*�<��q���^l9g��	'������^�&��N)�k��%Fu�c~B����KI'�v���,��M�ׅEAdż,[����%�WD����n^��\��	R��	8<����B9����0� �Pd��n	P|��q���4I��A�Y�w��i�	C~�R���,C�
Kޚ�я ���Ӄ�N�i"-7
���#:v��|��W��d��h��y�u�0�����T?��4�َȄv-Ox��l5@/����q�n{��@�F����8f�^֙��U���4ʒ��C/���B�4V��&a���<n�hS�]~2�<��h����jg2����!��:��%5p}� ��
�wĔ_��J�k���"��y6�Q
�"p8YjO�t���B��_!-������~pE��F�%��U�m5��j����8~�EO��x���Q�%�	T�K�����K��3~ֹ��-��x��#H�v��ӎqI�-k� m�cc��ˬ
��PRCQ���8�v5��v��y�p%�W+g;�Xxe,:�j����Ļ>�0t<z�m�l�5O '�� !��^��4�W��qC�=J#��:�}��؞���{�0S��N����Lnn��:颈*ĎSM��%Ǥ����T77Z��;X�x:L
�L��ټ�#'���|ۈ,�ǵ��6������F�HZ�.������h�E)o� 4ӑ ��l']�!�!�?*�5^��b���J�ιm�G�'	s�~Y��� �T�$�i����+����߷���{�lu��C������MF���ڝ`�0�O~%�Sy0.��?Y��-( �������� ��S��M�V �[g@�nk�<��mf\��#���S�����˖ 'U} ۥd�q��.�J�ߖ,��,�n�}e�d��2ڀ1X��>\ߧR�q)]�Ц�A~G�z�����i�.o ���/��x�[�`>�+��x�/���TY��ୂ -���{��#o6Y�� ��_a�=V��9Σ`gg��c���b[�>�وq>���X���է��z&�<��=��0�;�,Z-u�4����?XW�<{q�(�l"A��ڵ!;��`��P�ޓ��v�G�I�ؔ=��^{էEJSt���A5�b;�sJ��c`I李y6%=<f��ܛwj�Fт���=3s�rO����� b��w�D+9/��M�'�]$��;O3�$37ה[�d�,��%�0H'�s�V]��CKN��p�6��nz�ڠ�Z��=_�:�K��w+�uڀiy��p�FKp�5͋Ҹ+J�7�`"�\P
�X���}����� ћUux9�g�q�W�GK��£Qt�5�*C�\c�����6"��R��+f�"G�´T�j/p��z���o�;�ۢR�� Ei�|�H�7O%*��2����"���0�_c4e��1�&q�}F��^͘N����V��Úy��?Z�u�F�O��scZf�W�ĉ�f<!��c	(hfy�;�݂���no�4HCY���3�j��J~�T�_�fU���@ǅ�������M@E���qaz�bڱWV��[�pB�5��&�#��]���XZz?c�^,!7֥g^<��fltlŦ���]��Ӟ��޷2���؆#X+����n�#F���T�t�{ٍ�7gr1��A/P/���~W��}��`�ڧ�O��A��?J2j��*t[m&+�]���W������i��kɲ8X���M��C��Z�p��=t��, 3l�Þͦs�)ě�o�7�7<�*��R�����>�l�zo��9һ���!&߳F޳wPS�K_�C��1�����n4����`y��������$i�b�|���+fu��jF9\�
8�!��4u���USn��F_;{��	��s,��Ehw���}PZ�W��iz�߆�j�4v��|s�Wn�Ӊ�t�c��JD!?�҂BX!�o��_�¿㓷|q�<����9�vw]�~9� �r�������Ě������3��7!�Eȷ�_�"�wԤ�#ṃ��q�5�%#�iC}qpe^'�Ɛ@��F̿ �^ʜ2�뚾߬�6~�6�;��/�_�M�H�ۍ�B!t��c���hW�Y#錒����L�y'�Tk����S˵>
�|BqL���wa L<�
�"o�nli�L�Ć<�W!�����F%!{�G:��@Be��4�zk[V��(LUL)���U��q����Lt�}��9�F472#J�!7E�e��5j���GI�<H��Qsv��2|y��_�Ľ�ʸ���@f��]�}uOAt]��Q�$�0>�n.��� �sTx��z������N�*��2��4�7ޢ��dJ��u&v6ꆠ�<����I\
�m~oAz���Obo  GU݈� 7ڠ@�a�%�y� u
X��e�\���7�&��ľy�	)o��E����_���}�\�4ڦ��a 	�|L��+���3��V�yuo����/l+��W��� �۴)Ig��Q�j�D(8@+�ET� ��,��"G�^��#�ic����4�9��ո���#�m6R��T�ܦj�.�n�5�T�)N�4�UQ�_����z-�q���͑��C=h���� H^\�Zԕ[�2�',K�_cɦ�կ��p��bq_�Hu*x.>|�K#I��2볧<l�Yoܖ��e'[�iK�D�)#o>;*G�t`^UJ$ ��kP~C��#�>�.�}E;+�4z�Ҟ��8́@f����^�H׎�z;@4�K�D:���`�����Dh����69(E�~y y�񠄗���c�-D�y!zԗQ|�قzv_Hd0(�{��W]&�<���A&�-WxF.����i^�&��0wT�~_p�5bQ��(��ē�{j���ADFU7_��\��'�bc�LcGC�&�_z㡇�Q�Q�3��{G�j"������~�4�Yݬ��zZd�����aͳ���mr� �\A���Jrn#E���l^��3b۝��?k�9���abx����wњ�w�S�<�E�oڍ���;dT����/Y/f ��|f�g�I ��=Ӽ��?�b���A�����u� ӂ>b�d����� �g�d�@g��G �=�yk�z1[BRT_��2���ٴ4�#��]ib��k�op�O�p
7��Q�wT5;��!V���ol4w(�v1���<��~>w�Q�MR��Tm�??�2�F��I?4*-@��%p�h��0y�*��˓�!"�����|n.]���_��je�<)>_��=7���fY�D]�D|{����ո�W>�\*���n�̻ �?�m������В�S�_�1A��1r�u�-��o�H���d�7B��`�L�{�k�]o\&%�R�9|p���.+�#f\���	���3aZB�=��d"������d�sm�n�1�@
�S��֟�i���0��
�g'3� �|�X/�>~�F���%!��<^pr�-�&�5���*�^\+�go��+�=��b Y(O8���d�`ä�kn��9ZG����T
{i�0�i���a�D��ql��f�?�����ʥ�Ƚ��B|k�'��4���w��\�s��&�3|Fx�)M8��v!���ٵ ����-u��Q��
̳�z�zn~Z�E�&Jzo>Yv7rU��ȘE7�������I�&�nS冊�$���q�_���Wј�b��+.o�O�r��ճrZl}4�mݾ{@��}������4�8A�9���7�c����%(�
��s�>�B�5D�)��=���>�
�fs���QrƇa�O�%٫L	�'�ݚ?�o�vF��7!Wz?>G��Nl�0e����yU�	�����V�eh����՜�����&{��i45��O�iJ@�b�G�u�{e�{���ϊ�E˝/U=���\U�5|�[���*{%o^}�<���w��r�|�F���+d����F�[0@�!��(ר�'��cZ@Ș{����G�xD쯹�Fm:���I�#�+'����P�k.�QW6H��19��Xl�aq��W�sY4|W�i���|h9TBq��n��/����^�߽:���ID���{�0��p��|����V8렺��ɭ��������[�~q��[�K�7�0�Y$Wn�ȹ�R�c� ���7�v��
qi�F����Hs/~�%��o������ɔxЮ	.�jX̔#[�%�H�.YMz0O��Y��@�|�[ӡq��1�R$�L��f�J �+ynkw�h!�
!u_8�����4�bS����`�>1^�H�=64Ws~��FCv��YvL`�ǈ���ڏ����̕��������yd7mÞ�g��<ĳ�깁C��y�yQb(�C�h�����d�<���\l�ժ�N�d�4�%��?�f3 l�ݩ��r������&���4�u�r�5F��]z�YL*T�d�!�X��im�/�N��� uൟ:��Ǘ�c���|q{��J:���L�NSFܳ8��$�G�Ԋ��b�(��Ńe�fo#��W�`��<H������ы�u�����q5B����1�ԁ�A��n�8Ovg�T��R�w�hn���������h"ヱ����2��[�f�#Q��X���K�����Q):;�H&P�4�{��K�g$��	�>�9a��<��b������%V�F!���2
m7Z�2lM
`�(>1^�ݏ�K;͐U�j�x�S��PT��%)�K-�G�A��=���'VOu
�ha�NR��������)d��ߺ�������W�.F���ԧmi�Y���w[?99��]5�� �4��QU�	�岆�#m��ƀpC��7i��؆��V�����M1ܬ��ܹz����[d�z��ֺ
�c4��I�-�m ��-1�a!{�h�{6j˃/.�h��j�k��:T�\�L��Z�6{|��S�(�r��0�|�'�+����<�L�� MZ��Q���FV�c���;�z7	Q�`��!H��C8O�k�2�1\���rW.��w�"z�ѐL, }אx����{#���t$�t���PQ�����M�L��7�"��%`��׋p{�(�I�q��^?d���ݯ���5�c2{�JR@���C�χ��`�$�U��3Qg�%u܄�Sc2����l
��<��1��1d���jJ*�>�4рf�����e�5~��-T�&3Q��L<���Yu��HƉܡ�W����[O�q�n�qM*�Y(��lB�&�N&�||�h"�uX�O�k{�8h�U���a���Fh�	>o��1L�Ǡg�~BUa�H����#��� �7O4�8	�s%�/ө�w�3F�>��`W.4B2��pt�`v��M��'�7�&FsI�'�g�莏`�/^�ab�sa�rY��9�)d7�1��^�L�bx� 7�bw�g�S;p���3��8�:��hA!OR�U�6�{�%-e�+�j��c����}���`vX�6r�<QI�4��D��^��`��H���i�C�� >��h���o_���$Vcaմpt�vr��oF���L\^jmv�v̅��iZ�K�~7�8�;���8�r� �G'E�����AB���׶jյ��j/�V� U�|"��W�Ϸ�1D�J9 ��']�Cb�دH;��6?L��Ͱph�VǸ+�D,~4���潄eq��1n�S.�A��RXN�)����W��T�t��~�P����h' �1r�6\�M-!�TI���:ī���ڲ�`�Kp�?ܷ8��o �x;��W���FQ�� PW6Ӄ�')#e���ܸ�h�97ү�P�J1Þ�=�c�;�l@�X�X߻*s�F�g�d����˞��#m���0�`q�3T-�e�XAtx�]P��O���_��T�=�IS]�ڳ\W�{
��IX���I��r��L���(v]崥��
g��N��5�@��6͇��������S�'О�!*;]P.~�m�}�Y�^��Ur!x��T����	1W<�����ǧ��j&u�ͧ0IGl&l6kB�)G��Pg�[�M:bB�[���c�����OнCU��ۧ_O�w�91|���=�܇h�b#sV�O�H�\���Qd�X�
o*�s%�r��d�Mw6U� U�x�Q�h�N
�� ��+.l�t-�K����n_���ra�a�diM�Eh癃�)i)H������CJ**1�n���.�ą��P���&�����|,=1A�tϧ��B��4p	6U�@D�@�Є������4�@��T����z�ta�c���絕�ժaֳ-��G7W���æ1�XZ�Qo��m����o�?r9y�D@�)����e���QLp�W{��3DlrJ+L����4�2��q΃N���������}�Be���!���F���x�_�>�w"lG�D���X���ok��J�Үҧx�>_nlX7��cu�q'�� �|�g7w�ɱp��̊8"�Հ����RD�y��u�fkHBKk�Woݳ�p�����ۋ5*W�xW\�F�"���W�C1�o��k^x;���4f8I���m>j� ��؛��!���3��g��@y�����y�,��K����͍�o��fK�1j��s&����WN3���'��b�I�"Ar�Ȩ����2Rޭ�%ޅ�`ȁKQt�v�!l5V���pɦ�4.�8�琳�X��n�2n��pj��M?�ʁڌ��"8�x��Č���\��	��E�<���6�A�s�8	! �ioU��!~y�t9�l����̢
) ��n�3��A�IO���O��{t����8���Ft���an����2<�5?�̒�@��$�گ"1��8��ܧ��1�"6�=C��e0S��JdLUVH��(a�z���+��Os��=4�8h!@����+�-��.�'�N\�`��^e�*�N:%������Z�4�7tDN����R��_aW�Bl^rW���n��J�HR��F�ȫ��R�n�<��ڋ��D�M�0��?�Qu~t�dH�}n�N]��Ƙŕ����,@»1	��/�Ò�m� E�1��DwZ�T�<��:�X�_3`�u��'4=)���]�b��x7F�#�ot��F�Ɔ��8��ƺK	HR2��ض�E�x��L,�\\x�a�P���)M��U��_p���l�
�)#�qm/ �<�፾�pԉD��_�g,��|��K��e��W�Bcf�(���:��Oۇ��yo�B!`%���^g��vK����n|�e���"�5�PT'�9�>�ܿ'N�V"��ȶ�Pz�ʥ�f�\nm�u�R���S�]ҩ^M�+�T�e:�����"����2t��'/:y�\(_��i��YW�]3�0=����򮖈�m�N���X.���������MZE�k �����|F�mn�2pgr[����� ��8&1��!�΋�� �IIk�w�[�ӆ%��ؾ���T���2&^ß��z���.�#e��k���2f��A-�/4�`�Fj�E\:���V���5�^�t�+1݁�y62���;̧��48�F���[��NNh�X�T*�|n�?up=<�����Q��陭�(ɪ-܀"�6�'KW��7�l�H��b^�耂�[�t�vÖ��h ���U1:y����F�����H6fbǬśsg�C¥|��?��,��?�"0_t��@~~��^6y����d�1�'ْWI!S���D�S�g���HQ���p�#�rʕ��(�lf+�R'5˶�~�mE�K�*�J�8�0�}3����(�0nt��/�aN(6m��ZQ�O���g�78��Z%~FI�E�#�#S���iiTw�кýW�]��dUl+$���};
*a4k���1vm�������x�e !|� �T��{��C|w�\��xx%P��Q�5�F���m���������Z� �ꎥ��eA�8��vsb�,xS@I�QW�I��6@bۻc����U����a�nd ��7�W�X;ڰ�!�D٣���r��}<S=Ză5u�%Z��o�V������%?'�1��Aw��HP:6���AK1:o��Ko调��km�q$W^�.��W�V�.�q�����_y*�n�@�wX&�x������V�q�_V@а������i��hx��w�B�����h�ܤ����7
F�՜�m4D�5_
4�]��K����R9�N[B��`7����r�P�7R|�;��ޘ3�ҕd*�%�%��ë�"��h�z�gm4�vk�����B{�,c/���Aj�OE����KF�ƍp��:38u�9�[7.�es��rd$����p��;ͱ�_�f�y�ZP�U�X�O�e���=����`��F�ȧգ��ܴ�z(��e��$X���|�o���y�(P�rH� 4$��t|p@^`����%�m^�ͮ�� ?R�>�h���Gd��7Ş�$4Ӗ�'�q�fv�7AR?�5�(<�(��c�p�À�qǉ?,�s_�[9���=�GӍ�X$�m��\C�vhb�PҳvJ��h4����g���GY%�R�EB>$b5$�j���R����ғݘ������kA;�P0���r�a/Xc�n�F��UB��:}�u�yDG+Z2�2�"^����a(a!0t�ep�@�%�x�ٳ5� 1� �N��>��M���:��$��5�g�P�ipM�]wN%&_~
LUOZ���CI���8�3�|���f�2`i�n� ��dΑ����wz�to�<M�1�W5�a� 7����4���=o?��#;V�l�{��j�<,�gkEpէ��K��Mk�U�e��W���,���.�ոIm��rL�`�%�� !��< .bl�l��_"~�`�����<9W��6� D׼;�Z������v[vn�Be,�_<���[����������B.�q�Ao� ����l� =$l4nh������RODعN��n9P�\����M�@U���#&�B�:���S�j��m�<�`���mp�#���bW��\u�J�f�%@��2� a�lx`�2Y ����2�|K��0�B'?ZBm�b�r]���!���^k�T,�	*&������|fd��ɫ�ћsǮ�Wr������0���˶g�6�M�Ȁ���[�ߗ�{�g�w�L�C��+��%9����|S��u�<�\��c�Q���O+�7)J�Ѿ��z#�9}R��vo@�Nx�|�:x�������z���t%�q����O�Dğ�H��3�G�����s���|�E��w�2�	�:=Ny�}�U
%�N�;��=�gş�+x�J=��2��C]�s�{2?���T �ْQ�
�|��z�F�/h�)�M֝;���3 �zO;��z�������k�gK%����Dr~���F=��l�(]���S�>{��E=��}c0�v��u$�M6���}��@�a=�z���F��T�9*/�Kc���C*�H�n)~��M	L< L�x�T����A�P@��<y���=n����u|� �;W����G�r5���^���T'���	�����Q��kq5?Qj���:~]�?O�T����]t/^!�\����$:��I���8��x�c���x/��u�{��f]��=�2.�[�I��F��X����&�}�_#��`�\=B)������B{*7O�)wK{]�J�.��O�hZ����P�����.:�3�l�(�\��v�A����&��$xԁiּ���R��eAҨ:yT�@�� '�E���,�|�wA�l��Ua�����$�%Y��m8t��h}H�{�Fp���z�7r[�͵]@��rg��*͈,Ei�o�~}�k=��\�`{݁�TTQ��C>Єb 3��ѽA��V
�������p�k��D� F�}�Z1Ĩ��0P�"A1K"�КZ���O�c����d����H�<�����넞P3<>@�+��t��4I�A�\���p�}�l�vf��U3^1�~�Ԟ<�Vj�;FW'��3�s��AE̱>�6��������hŖ9e��#�ΈWVr4����x��1C�r�(8�5\��Rϧ�sBf��u�<�JLg��J��Yu(H/#���$��Q� �<��6u��J�<0�;Y�z|�ݡ�ڢ�^���Y�fE��QC���Þ�=ڹ<9�R��0��[xĬ|�m�"��6��Di�Z���?uO8[n%w�/bY���dp�a��_��zr� *u/Q�ο�g��4�@6���V�0;w� ,�P�Ĩ�ȼxs'��Nr�A7���������f�J��r5YR�6z�)t��᳙�X�W����ʔ��������^]�D���?�+�A[���Hm�B�ɮ_e&��}�g��-X$d���Ux�����
��tnum#��:>�� �5�PǪ�s:����O�	`�)��?��	��QO�P!�B\6��\�u����J�R|�fL~+Û�mD[I�(��4��8�"G�~�F3����B����I�9���c�"�l��O�:^O��H�;\�7א��[����p�K!��5�&~p�޹��y�o�jx~~�7���0y��%�U��ͥ�|�*�$+�=o�vu�`�̫	��`�g���v7������05-N,�خ���w��TN;�%��B����P[��Gb���7A@�-	B5�u���lϜ7��e��:NQ��~ˊ�ŢZ�('�<�ͻ��;W���"��w�+�(י!��t��GW��k*���O�aC�˞bi�"w.Q�X����AV�7�ꈣ�C/oٸ��<W��:���3�u��h�ba�^�KAa�Qv��W�y;�P�C��Y{�ɗ���Zcm���o�$����@�TƧ`�m�O`I�4�ԍ�)�({��a1w/(5\~��ʏVҹ>�/���H!�P��0���L��e3�+��	b;�`�W����f[�g�`��ݟ�[�j&�Տw^ �������q`�`y����=��b/�B��@�	���p�+�L��e��������Ө�2�v�T����o܍�7B,kTc�	�P�+!at�{�:Y��L��T'������h����x۲=}��3\Q�~�(d�|Rwą̟��������+��ba	6ɏ���M�	|�!��HֽI���FE�U��X���E�N��h�u�C�19V�64���M9���f�2�c�s �Ȉ�.�qXJ�~��g	>�ʒw�j�!�G�s�9��4F�������C���D��[I�V��D��d�*q#lN�kAqz�������8%�?7�*sh�<v=�F��H棔3�.�فb�\����#r Ψš Κ��3��"S6غ�@`��౼���+�W(��&6
���ضC	��1�1@���x�k�h�SRo��p����������)�?��o�$�u(��ON��`=��Ǡm�G)�˧Hh��SJ1��U1���R������l���q��d�����|w=ª���-���''P�(V^�	��B��4Q$T����HD��%.R�� ��]Y�f���-w���R�	��!:�
d�E-z}2`,G��-~=���d}��읒S�2%���1)I�[A��Ϟ>��Y��a�RJ�r?��:n�4�GQ����:ҡ��?K��p�
��_{��D\����EU�F�+
Wb���A�y5�s�[ 0��a,�1Uf��$�;C��3\�2�;=�w"��y�C��r�
�fn8�{�Үg/�q�v�ƀ.gZ^aiu��A��d�?��8e�K]f������i������;�OZB7����f�e^Ad��95K�ϱu /�0��O�3��^�۱�V�J׿7n**I���"��V<�t�V�lb	w��Mk�cǢ����[�,�P��� ��M���#ӳ�P�X�{k�}���[��hubb۪p���AD84ma�`F���i]Õ��� PgL��4�����H��*ص��S`ᇟ*�l~�X���8�mFg�����p�_����Ĕȼ��zMAc�f9��#������	/آ �F������/�R����K��ݨTy��ǌC�����\1L��p����ϤL�º2�s1 �ߋ4�7pt*�HxGY�F%	H�]eo_��e�>��ʫ�k��A2�nbӘ��B� ?��"!�T=���N�L9�O���G-v����J��,�LS� p������'��3��P��}LH>sN����߽�W�ƿ*[�B�u�W�ܙI���5�Kj�l��]��P��X�Ki�nEq@*���.6� �[��5/���"|oW	>~xw�HB_��2�,>�Z/�{�ĻI�\�c<��Сd����[EeS������I��VѪ��-;��~j����
�V��*�H����������x>>��*��ꜢG]~ȯ�t�ջ6}���uh�Y��4k�w���I���� u��N�&�#2I����vy�G������W�C�Iw}}	����ǡR6�=���`�$߷f�[��Xs��v�(a�_�S�թh�E$w�K��@0I�9��R ��	������c4���fS�dg�y?3*�l�T'�}�a��_P[t
㺇�`|0�ؼ�1�`cXMo�o��+��'ݲ�����(�"��<ر��j�hh%��WT�B��N����BuQ�]�b�K��O�,�L���Ҥ�U����o����`;�� �Y�[1"��3����BY��i���Zg�5�Ȑyݏ�z?�-eԸy������5d��x�P:��GY޻� |`�}��۽���`�M8ŉ{k�^b=s@��nUTY��(u��dɭ�i7������Vٮ�Ԗ�9��Z�Gp|\p��YB�:�?�B��ёq���B���Q���ϳAK�̙�;P�٦�������i��,�$sr����4h��M��0ͺ���h=6�A�����i�#�h�ǌ�n ���>�������Sz��4
M3\�3d��I$XCԖR�U�3� ���a�C�4q0���Gp��V<c9zaM��Ai�%�aE��āY�!��i[�td[��xȁ���Hgͤ�%��ء���3�������?Pzݙ�c��hѻm(Ջ����߫�'��h8Z>���k;<�M=��I*	Kcָr	*�!T[�J���Ev�������*��Ոkƭ�'w��@.9=�.g����С�1*w�fV�����Bz�3�$E��b|�<em:������2�mn���?�  ![ŵ��q�h�#Z��R���X���y1{�O��Vj�k�����5�J/<�tD
d��a����m:ҟ�4KY��mRGk��R�%'�n�3�y#�����eA�ܴ8�C"�����r�4�~H���tn��\\���Ki��J�h��P��ۼ������_!g��)��9܍�΁�MA�l��&��k[@�A�众+��7�,r������޹fI���i��K�/M��{4�;SF;r8�H�؂a�I,۠^�˝<G�}1���0L�T���o05�\R�b ���b����ۢ�7��~d��c�I�Ug�U6��|���S��{���;t�Hnꄛ.y�Vg����&w��G�>�ǱG��\_2Z����	�|	�~t�]�Т�]�D��w�V>>J���ԛ�q�R�Նn�[�b�a�*���9��܋ŭ�i���K�à�̌3��0Mҫ��۔M�����N�i.��j��L '	���x,uq�h
* �]t�43�ۍWi�����OSL��Sx��H��\��U3F*�j�Ώ/`�`4p�	ݾd �𱮦ߑ	��>��o\V+A�^�L$ \ށ-�g���NA�m�ɷ�O�j��f���d����3L���Ǯ,�|l����ao��cE��d��]��h�����VV��վ���^~=d���aJ�3�j�64��[("uQ�'M���?�Ιw�<��?X�=�6�J��!�;�S������rvȓ�ES��D��[#���a29�/r�_���f|�dV�g ��~�I��2ۿ	��^J�!6��)5j���r�0�▲F�]c�~�m��CT�vb
p��I]��uHC�L�ɀ�(����!;�/��E�P~]m|; ����!wBt��X;>���aN�Z�����;Ͼ7��ySR�ї�r�b�l�׈֑��Y=��j���\��m�.����ߩ��pN�ZUS���E�3~p|�L')A�	;���~N(^�gW���a{_�&(jR� ��9�7_���[;t�~�x�4�0h�@jEmjm�҄;׸P�V��y�կ f��]��#��v»�]F�M����qF���'g_��MC�h��+�7��viVϖ栐 �vI��r�t)yN��z��b��?!�h��XM��r�RJT�+�3�PD�/-�g[�p���y�W<o��C�����HۚP���~�u-|�G�\q&V�w�#��b5H�VX��l3뎗�l�.Y��EB������^D�E1ъ��1���@.��C��"����Y��/�u�}	����$r,,2�钖�iFQ����7��ds�����h�)��f��i"���&m6�v_UJn���џװZ�R0��b
Yc�7'bBl6�q�?�e;�.�o�h��뾙"�W��ZW����2�U��=�~(ƥC�1�ȅ����ý���Kf��"����t��l�����N��^�G�e�Z��W's�n;O��<���E���0��=1�=+��X6-Xr �}8;f���D";���y���x�Ŧ�^���&��u�h�T�W���|I[.�du�4¯J��5�e.�Ago�96�LNAbu�[�2�Vw��Q���xmpB:�M�SEi����%cF0f�P�@Ǟq���k�T7s��
�ϻ�
�9��	M57��VAf��_Q;���Zxp�z�.�-���iW�o��S�i�(�j�b1����Aƶ��C��F��K����&m�fˆBf����IVb���6w��g���йQ$<s�[��%+�����z!�Sn��n�1{s�>vݗXQ�f������P�2Tjk�B.����`1��C�J�
�xX��9g�#�V���D8?'�3]=�{��F�U���Uz�"�}�Wr����B�%��j1�j{):Z��֭���X8����,�9��<g'_I� ��M��{�{���ϾNZi��b������@"��������gȦ��dV�2P����*��4LӬռ�����)��Ќ�em!e��p�p0��wV�2�_�i��1�j 	�،��]%�ghUhV4��P���:yq���Tj��7Ǿ{մ�7bu'SF�C���N��w����b4�#SW�DK�G)��1�{L3|<Ֆ]�0>�V�gw����l��TO��L�֋��� �ן	����K�T�7"��Ӝ ��ˆ �`�z��e&;<�B"���,��% œ^�n�e���a�w�6�~m�F�/�d��/ڪ�'����	�A�uXu{���/aJ���>�5tlgP�hd&^+}W=�f�	׬Bd!)z&#T'���'Va:
!� UK�Ǽ��h��&N���GK��P�N,���B8��5�&������9Y������8C��z�U.<5��T	���i<�;�~�΃dg��%bJ`_E���,aR�,r%��_�A��bw��A�5Y҉�f�d�Hܷ�5%�����߁٧�o|s������G���'�=:��I������ȅ�Q���0��Z�䯶
;8!�j.�6�ܐF���Ѭ�5q�׆C��^��+�4d�P! H�f�C#�V�Q�	��a�d%�"V�1����A���3*�wH'�����Ku$S�S��~U�?���.hLxg��4ݞ��S�=b���H��"j�<A�F���1�}�p�ި�CE�T5����v���
`�o��m��7�B�{��Qqdo&yՊN�:*h��x�e�?����"ܖ	�Ύ�YO&|�I��j�JHי.�j��z)��	V�:�A#r$�M���'G�t��v� |�!�R�@`�r�o;��f�@��/�OR�&�n�1��1PR�F�	�"�:�)��ˣ*Wi�z�B��2kݥ�E�v��ń u%�Vy��һ4t�ז���d����M�u�*fCe��~asn��虗�T;r�QLo�f����}�rtCV�jĒ.˭�r�[\�1����]@G{je4��Qj����a�OLC��ȟ��v�� �W��ҍ��Yv����8ڝB�,[�"Q���pN����E4� ������,�Ρ��N?�\
�Po����3c<w���$B�1m�cNb�E�^Xͣ��1�4bc�JB���,K����LR�;ްס��oƀ/��瓼�jZ<��*����c�ٴ�"���-U���
��]�!��*zM"j.�@n�{�D�ܱ��	��V��d�8���(5_7���B�訵`���+N�����������t�mL�Edʆ��SR}y�W�ཟ�p���w+Z��,����'%x���P8���`+�=	��d���'�X=2i�}ܭ�r˧T���=�О��.�%#n�6w��|%1����/񁖗���B�9�&�*�/���@���bP���7��	|`6� T'�����&8Q$�"�/���6����<��bY�M�8z��z
�iL�R���
�����bG�{�7�M9��;Im�#7{ch���r��!�Ğ����q �}��A��޹ B��
w�B�,��6X�w��f�E㒫k��]�p�z���ZD��[����%^��^?<!^^Os���Ń���^��8��w���yn�A�$N�4�Ɋ:�e�(�d�@�-��T��]�)g���}pCt�Am���^�]�À��.u��	����aY'"m(
WR,fE�G~�j[Z>����o����/��L""�h��, <U���.�r����o+1�&):��Z�5������=�ޒ��q8R�Nki9�]�YW����V��h��7�G�[�:���ۜ���������1xyꏖe�.���E��G�͈�~]
z@���S���+|*_2�L�{va�8��R�KW����"Jm��6y"�g�>[��Y�4PS�k.��rm�����<�u���C�ɧ�t��"?t�2�2�Fd�?
|^
���}��{3� ��%v�<7-Q�&�?n�2�� �Ŭ�?��`�vG�zx�J�&WWDK >Zu|�� 9���Ğ��e�n:6(y�O��6�k F��Lr-��xy#�To�/��KYë���:�W��& h�C��#��p<�\�����&�B�/;p�40xآ�p;�����W�Ѝ{?�~H�z��!dp|oxi9z*����D���+����7ŁP�8^�����S�Bz�g�͊�cr�u����ة��t��Y�vl�IN�L�)����R�ցK�fv�Ϯc���'��������/4m�п%U���;��ä�;��+�Ð5�G��V��GL�f╎�2p���<9d*y"���`���ܭU(X�`L_$@�|;�]ߘ��	�q�'���?�mX�. a��s���&֖z�&njd���'2嶠Q�#��4+��؆�X����8ͪI�:/�w� ��c�xRF�yxv���د{'g%R87�NuH��@��5���!�&X�?3��_%�uY,���O-�̀z�
���uP�u���4Sp���Hc�������Y�w�Q�D���C�D���x�����U��_m��Xu����6����l��mi<4�"�kR��S��1��,���8b�S�k������<���F��&��뽘+� l�u�c��h��|����x'��9�X�$o�%�������!,�/�6_�L��$j��Y��KV����7��g���VB��UM��Q�:�"�?�aVz��a����YG��稔��=ԉ�J�U2�$[�����c�� �S=��5=?�L
�3UY��O�kɼ�~=J�EYyfՍhx+��ڤ4���y&�UEE0��o�xߞV�5��0_Cd�F� >`4�D��t�,۔�C��A{Ag��]8L#!ǖ�`$':z��-�^<m�66Ÿ/"�]��:ZUfV�3�es�37�v�u�k� G�+`��Agڒ��ò�A���S��(�pS�öOT��A���QĹ�P�sV�7�!��ˢ%e�9�Q�YN�qx�SWi�_!\�SO��f��/o;b�_�c⿷�L�H�ϏMl�w+e�������D�̽�{��k�.`�~���_񉑸Rl�
J�uz!]
H�K�SU��'�F�tl(�&D�mq�#"J8�����;MHg��%�~SJ�?#]��G��:Cps+�%�W�	!@ֽ1����A�t��5#�@E�;��`��6d#�]�W6*=7��76\�-��>"�&�������`���9�S�0�')Gz5�,r\�ä��8wS�Rf*-����,���Q!��eT/�>v�ߗd�g���C(X��D-�zs�j�N�5G|L�}�6t�h/��R�`K���>fksl��`�����[��*;�I<f�U�+>��uu+���]�>�mRUTN��4��l�FU7:�=�]a��ϊ��ރa�I,e�&[� �	.�e7߃Q3�*�z�0�ضm6�MT�ͬ'g�*P;���:�Ƕ�O:�D�).N��P����r*��k�e�^��J�J�7-���O&�2lQY�v���!wV���bѿ��Q�h���UuJ�W�Zث�r]��x��̬�&��:aM'dk�gP����x�gg�[S���M��};�/�*�a˹�Q��5����a~���tZ�Kp��ŏ��J>v�ђ��o_=���k�G�I�W�k�g�͉��LQ��0�'�C�W��B��Tw��WKEhr��DV�� k��"��^5�E���j�u�%�j�x�66E�(�����J()�O�<tMl� ��/7���KtK<מ
GQ���:Df�$��a�H�&�&6F�����W���`!9�*BTT ��D�n��˥��=� ��=���	�mұ�)	9on�����V�Y9O^��wK�>^�T�)l��gl��g��szyo�-.$�����o�L���0�8R�c����[k!������7[eD��Hi��P)��r0�xӌr0��@>��i�a6=�=,V�P��y��3�bh�<H�>rc��mi���-zn��T��P7�������l4ECtCAة8d�!g.��Sq��A��0�}L�]}[�(,�������)���i���n!Xak�n�P��Zv���;��3������3��G�"��\�Tʅ2���+J��`!�"�3Ŕ��S;��"k��j���?�������c܆q� �@Ǩ{��_�pv��eV9����%b��Y#����x�.��q&4
�w�Z>B�+k� e�h�����F�n7I��۷���!UY�86�p�2O�=�\��4.��0�8F��6���H��V"�R��F$�c�{&��z�����4���q.�`4�=��o]?��]��\�аSߒ#n�FYs$��}�d�"�k+tt�u�S��|hb�6�5<%��_`跁r��}�&0
'�N�b��`������󜫵>��Ǣw|�������4�p$����Ǵ��N�w�g�>�Z l�s����#�ќ����
qt.,����~<��L�K�`��M3:k���A��|�8���:���+N� �`���S0ߟ����Y��J^�F�����l(���1��E׸=,<z2�wŧ"_�싽+����`�p ��s�.�7l�g%�Z	�Y���?�hy<��6���l�;`�^�)5��h�<b���F��ɏt��lR�<I����aN`Z诓�nS�-K�좐S&: ���D�DV��Nefb�J�VWzQog�(̦���.z��H�g0E�vn�^��{�0>
J���a�gL��>�XI���̓-������H�U7���c�S�qf��H�/�L5���ȾD���~A��Dv#_�Ɨ�	5�m>&����έO����3h	��~Dk�R����S+�<.��݂Lﯪ�c���1`�t����$�ys�!`0������6�٨��R�5�?εo���2�4}���h��Q���:L�}����aU
~d�5�RZQ	R��:8Q�Jȕ��!�"�
e�����ٙ���ah�=�tq��՗nVt� �f`��U����[L���t���H;j�UhgُK�]`��}m~������>�~�F�<FM�6��~��ql�  4�a+��1d�G��6�|�Ø^Rh�5���r�n�ղo^��}�;{��-"x��ݚ�^O��>
G��r�|�>�D]<gh%�C�� ��z����1Ep�(��*J��}pG5���**�j���$�^زeI����TC��<c<jK�J�L^˃��֏�,��[,4�^mX �b�	<�	i��5�6����ٸɵ�t.��"���#Dy�L�Ƭγ��%��K�T*���(���PWW����d��&��(��LM�5P#�{�ː�7�3zB�ϩ���lh��$+e�����a���x;��-�����A�Ӗ�=���� ��l�x�<����hGC+Y=��!�j��>偊�ưb��)��Im�:���*㲝p_�`L,����P�-�Ҩd�ʡL�-G��?�P0�������yܸ�ͷ��Lی������d��:�89�C��Ѩ|��ޙl6IWز$�BÆ�Z����hO�*�Þ&	�,�୔��x:z fW��E����(�D��]�k/�fi�<La8�a�����<cı�y�.j���9˚i1����4�=�>�nfB��Da
��!�R��5��>�T�
�L"9{�p������'�x@�1�CUu�� ���mÎ��w��9�zU���*��bi��Vf3}�\B�;0�n�@o�Sd�dC�f� �-��(Ca�� ���/Af�����vz($gj������Q�`��Ɋ��&kWe.��p�+-�G�cu�o��qC���a��ak�zA��K�ls	��{KgR�5�C��$��E�9�mi��\ZT�� �5�Dk\YL2��B�wN�;�D�%!�0B�<�O��Gd*�L�=mNί�M�iR�3��NO�H�6oa��N�T+�����������RA�g�u��&��9�eF
���_��~4r����\� k�V[��m���[�J:�E>���*$�_��A�]}�a������b�.�59�AYI��ݨ��e~w5�������le����� �v%��c+!;u�r9�VO��Q�ѱ�^L~~�6?�Z<�I�#��J�� ���~O\v�X�iP�V��n�ލ�5μ��I5�'h���2Z���������
a��B�� Rc	��bC�F�d0g-D�#V���j�x�GK�qD�
�NM�_�ͺb=K �IC�&��<��\��Q'��nz��I�������|g��}o r��yM�;+ځ���N�}�MO_墨���l�*�/A5�Å�Dh�� �tT,#���J1�� �-B�7-��U�[lW�y�c��Q�q�k�������a�B"�²{�i~B�Amq�<��jΏ� Q^���p�^C0���R�!�!���s#�3V#=	��Wq����WH�܀ڹC�k���L�,�0�n��- X����4�E����|�P���_�}�]�'^����*�L]y_hz��@R`�<�����A�:��I:����3�o�^J1�����޼�|p��|W̆��{P[ =#��B�Xgn
&����+�ע�T*���e����gB�`����eM�������8�0b�~K����>1�����q� �>�n-�|W�G�
^j�E�ؒ�(`������۟7�@}}�V����h�?0���K�PhBcT����KP��ߣ�t����G��Ĭo4*ϧ�ܧ��Q�p�#�J*��.�'w�%��|�<*�7�P����_m��'@����Yfy��C'{�iI?����3'��;;f=R�^L���=��)8@��%S���Q����E5�k���u�x���]�wf�7�]��V�S��D�D�D�݇���/��z�����+��^G4a��s\.�I�P���пf�.QH�q�Gz�KH��(�+�p�# ��qI��0�ׅ��9�pEt+�=���4�\O��"�Z*�}r����6�g�<�{\�|�@���V�Q�d���Κ�4d�#�l5�%-��[k��x�/�͟�s���J�d�ѳz�g�db��:`BӺ�C�MO�?��K>���e�M��e7��D%`.����Y�<y��`2�>�H#X��T�m�uSpJ4���C��� `u�SG�+��8��ɫ�A�EWX-<��p�ub��=� (��?�v��a�0�ʗ��Pʐ7"Q����u��
z5�q<-b�%��L��"���P3VVT��0����F�,N�"�F�7ƶ�`LY79)�V}C=�n�\���Xv�����FYc���uf��@U�����B'xX��V��z���U��a
��Ȑ���hУ_�s�|�a~_iq��qO�~§���⪊��0/�k��H�ݏ]�~T��,�	`C�۱⡬�_�O�R0$����2�q�~l���Z�0X�Z�}��p}�������kH�}�:B��c��Y#�s��B5yp��H���Q���{���-Y��@�bWLM� �hs�#��7�1������ؔ��$l�6��#�� �Q���vd�*���	{6&QiPUs[m��6�=G�:�DU�e2t�o�(6	;�c�r��M���8��L�w)1���E�}!w��Sɋg�B/$�tHO�$�{�"�a.?�S_	�E��u\�n��k�ب���z��JT����O'P��/�9��l�����6�,Y&u�L�l�j��L¢[� q�j��w�(�'w�o�@�(I�O�-��)�sy]�9����.�D��*\;@��M�P=�5����L������ܰ�𑰲�V��C,�l��!1cS�z�����/������������0�3�"���m�?���yZtS�^J��:� \ۣ�	}���B){�*��0�\�<��d�"�c�:
��<8W�;���d�ٕ�M�s
�{%)�TU��hۓkNj^�\G� >�X�d]���d���`
/������-"�ʌ���cC�PU� >�����R��^�/٢��.H�^�)V�	�/r���������D?H�!��剏 ǓW���j�X�lR{$�.�>�9��7Q�mn�:J�n��D��wz��0���%��'�������YŮ�$��f��'�q�ǉZ��7W�l��]�xt%�6��=�??��	�D������e8�z^�R׈J��@!�S8�Q�i��3�9��2���W�~;+��Xz3z�:�ӑ@����*�<R\N9�u����#�����h�_�B��z�����G`0�UX;f���n�}�:`Y���hd"FӺ'�X��n1��78��\��a�k�ލ4�+$�qI�*O[��û�MU/�dW!O�:��!W$ƕO�d��S�}fyH����Lq���t���\2$�:L���xD��2��HAh��Klq�<�VZN���o�w�:k�X��"�c��-���?Uo\��V���;B
�3�k]3�}^�M�k.�� ��̨�q�\�O���M�HfZ࣢��f�+\��	+�궛9���
�p�u~d6��6�p�/_\���gC���Q�^����ŹPx�L��sT*D,A�F�T�-��	j��/!s틂W�#=�'{!����]5��vA���W�� �yx�([�+�#��~�u�r�f�w�r@iǜ�&�,����;�4��!dN�:s�PW<.�/-E��|.�Mv����%��K��^�i_����?^��I|?���^�N�D��Gۯ ���x<8%�6|��I1�MC�	��G��aPU������A�]xյ蓭x�hA����䚚q~�<UqVN^i'o���vM�q ��i?�}��p�s@��4 (���%�_��A�'�� 1�y�'�U�)D��x/�����_0�ˆQwьC�6G�j�ܱ��,���{��C!o<L�c:���5��wL#��3Y��>�%�*�(�lVLX�=���^
��V yE���
�L�/$����U�B�|�łP{!�|�3�c�<��ឿ�1,�Ҽ�վVb�T:O������6�u�9��)�ۻVX�I�Ǳ�`S���5 $=�}!n5�1�5���)�l����n۲Ϲ��3��:� ����E�j^��}�^/�ޗ��^ؒ���}3n/�`s��.Yf�ቪs\��ⶫ3������C�3,#G0����|^��j\��d�_���9ݠ��}ˤҒ�ڬ����X��Idl�Ð`�i�|Pܽz4l%"O�z��qh}�Z�-3�S���E�����9~L����PPj�Yʘ\/�J�}���EF��k�*�n�T�J>�;3S�+��v���Y��%��B��A]����]��*�7�闃���2������ԍ1�v��r��sV�H)��h��<���/�+�v�@�Ng������[��109�yJ�9	����^��$g�t>t=�-|�nb�!��6��:��k�%C��=TI9yw��p�1���v�}�!�{�'��Q�!p�Η��c���Cʎ݊��[����	��D�>ECz����.6�N�珞<t�'>��8[���m���nA��{Z��Q�9_ ����.�T�0���N�Y��M�R�|�z��<�4q��i�u�wA��﯐�g�<Sl+��jA)��㖲5�+���8��r�ih~�	?��G�^�i�aLo�3���=Љ�i.,�3��5�e��&�*��>M�k�C�#����1�&Ƌb�l�IBᤢܲ�>.M4�*��p��!�!��ջ���
�T3�Nx�4tm��M&��.�U�S���8�P�i;�S��g��nq��B|�܃�Q���笐-���.ս�Fݐ�� Zc��T*uy�3X���I���K�uvolDPӝ��H��:�(W��+F�|�X�+�q��0z6SV�!|���#P�F�-ӛ�Q	x��ڈ�-���>����a2&8���, �y�s�����~���IZ�#2rJB�w�-�y� �0I�os��r��n��'�hP�uw�~R)T-�u�	�� ~�U�?_s*"��_��MMp)��}s��A����2p���8��#��G�;^k^Z�-������N^����0*�󕇏��t��V�s��q�DB�4w+k�3q�������.�(�n���\y�S6����V
ב>E�h�3yj8r*�7��}�5�4�Ȗ+y�SP%���~���Y�s� 4��|`Rzao�S�i<w��=�U�Q��Dрb|��28��o_��i�����4�=9�s��0��fX��ye���G�$�����0:����.��g~��@"' 9���0S�4`H��Ǔl}/����<�������-t\g&����R��<2 C���YR�V`�.��늲Bдև����G�v������a�=͆I��ev��� O��#i�j�e�ĩB��0��M��s������K
`���1P��A2�k5˅���!D���JQ�i�Vߨ��u�ZT�Iy<�R����8k��s����\۫��qx�vW"w�NZ㕷�TX=�n"��?��=.���)���$�
���z�|8w�������a�ּ@�uO/M� ���ڀ7]޳��'s�&?k>�����L�'cg�j����s�^�/�R�6���M�|��T��^��̳��:	(�����}��V�)�:9x|�'� d�i��Q!�^�>D�S
�gUGNTg2��(k��Ũ�ʫ�Hѧ�ǈ(�W���|Ǔ^����I~ݛE��^�]�����:�yyR_��ǯ����6L�ϸ߈As� �mÛE(��nG��{L�P�.�uq;n!�/�]�����V�hQ��N-��.]���m \D\��1ϐ %%��J�l@�.�M�tz�@7=�_��|�G�Z	���t*2���R�Zo��#pv.g��M��"��&�/�N�nÍ�'��	�p���flUa�-9��@�UVh�/�"M)Qx��ť��(�W�~�_�����湐�v���7�+U��Qr����cqL>�i�T&���[�}��Y ��e~�����^ɨ�}����s��h�֍l�(S�y����8Q�D{_Jbgr:��2��Y%ęC���*	�s�����;sM~��wr���ڂg�ǝ[i��̝���*'�v,�%��Tk+\����	����p,�\c��#�fI�jBܾ9�m
��H��M0���7��ϴWg�����+����[�b�4	�Gߗ�9oldW, ��s~gb6Զ��m� �vx#���b�n׼�zAQ"�,QS�\3�Nl�lW������x"aV�,M^�+���8�)��a�9�שwYOa��M	Q]�N��<�g���g��rK���UZ��>9�=]�6W��z0`�������
�i ��2@`��Yg��ā��](��e�w��"A!ret�P�\�l�ZU�j�x�`����}�#�`���qu���<Ģ��S�Q�`��O�<�k� W�}���Y%�e�E,���@�X�3߄o���T��2a˛>\���e��r�4{�~O�����+[\=��D�h*oI��&��Ĵɏ]���e�e�ϟ`+�8�d:�U_�İY�C9N����+T�DP"�^�BKӯ\�r�em�^���m�z$8�I�X&��N;�������o�,d��������8�2��Ş����Q<|t�a\S� [�6�I��z�������.@�b����pD6d��؅s��v^^�)�I;���D���!Sܘ�@���C]����IH��6o�C&�b:N����/�n�0�!�=��k�����+`����q��o?��q�;V���5Iѩe�4�TS��bY-�I�N�X�R��x�:A	$}���S|�r�9��BY\fQ�#p�&y�xt�"ӈƈ9�w�l�}\��o>}�D�T��1sqjɇ#�k�D�sD�_#��o�˳/��ٯ��Wz�v��X�Ew���$����URQh/
�dgH\p�UM�n�h�����-ySɊ��{ԣ]{�m�(R�Mg�(�:@��۲[
d���VA��g4������o�� ;�v:��K��%XzȠ��|�rk������b�!A��O��>H*�kEɊ���w��Kz�_le��"���%�f��~�#�o���}�X�:f{��Z�?ӛ�L�l��s$��\��`|��7�|v %e�켍�p�|G���-� �b^-�6�J:kƤ��J�OrFyh���<��s?��C���:��M+� ���tKp�����e�x�NM��ki@�9�.��|e:�E�!���&$vm�H�e��$I� Dv4��z�؆"�^��˃bc[�WI{�S/2�n�V��,��(��x��#�KKܙ��ʣ�����*t��&J�۴A!yd��1B׬��.�W:c;v�U�Q�J��Kp�]����}q�)�g�^���(
���ꏪT܏ԇ����k+:�Y�Emd��'��:8֢�g�&*E.���܏�_�����g9u&�l�;4l���=:�Ζ����0�_�/ 2�<i�4�p7[߭����5��,��5Wg7�0�D#����s�