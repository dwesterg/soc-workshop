��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��/E���3Vʅ�����v���p��A�̠m}������"�|7g�f 9�����9y�ކ�������M�罘O�{j[_Qg>�1�89Q��v4ac�ʋ�Ȍ�b\8����W������K����R����s��i�vrr���ܴ�<%5�s'Y�G�ӣ>�$s����
�נ��{�%&����d����m�kB8^9�ҏ��R�nL'qn4N_�����l�C��l����l�J�>�Qv���|V y�e��݇�ъ%�=!; $K�/Q�]w��{�<�r�$fC�=&	��@DKd� ̮wuV�>d�ǝcm��oe���I��Y��c"�!�L��ޞ-(���װ�z2xz�S�L�U�1��5�t-K��:55s���AV��
��x��ԇ_�@;9��e�:e�SQ�������N_��$��0yK��Em �p�U,�ܴi��;?9�-�:��nz�6�"x�6C��;�cV��L�:��4`��0�U<w�?`���,�31!��M�=!(F��}�#UF��J��Xx^KXV
�	��^%�_�7bq&�1Ь:ܹ"�\�H����J��1�H���e?q���P)!ْY�#��h�}��E?���U��� {��n�L��3�~Z���1&�5t�޿�̬}��m1�0T;��EI���9�_�
�C-G/[Z�wI�C������m	 V��Gу�1���fW��|�����u���:�\��3/��0,Զ�ed槉>�7h>��t��T�6;Umd%��uuE}�X����<'�⋕4�Y�෦�ve��i���t���Z��W錐I`��ȫXe�9��K*B�*�:�ɣ*���~���m�,���*�.,E�]yQC�\��c�:��x~3��C�t�{�et�<{�rގ��jL2.ڀr��c�H��Z��`�dm�*��i04��xwy��:�{c�]���*�ˉ�;F⹴=�.�~_�-�-�A<�b��� ���L�t�ĿN�>g䞻���yG$|�&}�'3����22��0���'K��v�K��S���&Z��&Uθ����̵u� �����D�P#�P�rr�z�%�,�T]{�FC�xU,q��K`�� y$��1���,f�`�"WOKG�fG��o�ř��OY6-p<�ĕ|���X�3�r+�x��n�P����(f��5�:�b.��Gt��i����[,�l/��n	�y����Q9h���[O���;����?}�~��p�.���;@9���%7�`�o�� _[@鯬����u�K�Wr�+��^@�qM�?:�%�ݽA>>�+2�F��4A�}�F%�?����]S偣̇��iAl�c���x+o�
(�ά�0�Mt��U�+Q��$�J VS�J�� �9�v�+�x|}6�
�Q;�T��Ĉ	����GJg��Oϣ �qL���4r^���̖v豱��:'wkLڒЕj����>O���OL>�PZ�ǫ8�MބwJ��պ|mN��nn�5l������`�b� ����%�����k��חg";P���RmI����]=\��n��2)&����	��?69lugB�|��'_�n\��H��N�.,�om�x6�ψ�2=�Ƭ�҆8,of�F����)��Rؕ��+m�� �i�(��j.3%�a�U��@�˸(�*w�fv�6�V��	���7�y���G���΋�u��j�W�Ld�n{ƛ�Z��s>V�H��_��_��Ë�lb��(�Ǜf�ӗ�;��͞���H¬�%o��p�����k���K0k�����d��k܂�������f�W����<�ayqĽ�1�U���0�v��X����@+F����'����]�Vt���%I��S�\��k�����C�]P�<`P��� �BY�"�٩ �:��1���m愤�X�8z���݋g�Я�E~A˶�@މ�H4������4���4+щ���B�Z�l�X;��z�K��_D/�υ�sMƵ��8]��?�Fl� H��.Ρ+�����AN��\3�8nE�n��*,���= �đO?Ƴ2wzj���:����Wa���(�����a��$/-�FMg�CXM�ӿ@�l�=z��?�]���N|�5lV@D^�L�h�.Ffs��,}+�����՝v�#�������Y
kR���w�H��c�y� ����<�5��.�ʭ%��E��Vhp�_���(h�W��~�o��>G]p 9< [�n����S~?��j��_����״q�K:���Hl;~%w�!��Ӊ{/:>x�[�����/I��[$�Al®z��'ӡ��'M����5{�lT���w�/(%�������Zt{��j	vV���
'�%��L4����x�vwz�����L��\��=S���#��V5.ޯ_M���/< ���~����Z�������1X|R�y9Q�ЪëB���dJQZ*�� ax��E�i�ș�%]#')bih�Vla��I���N��?9|��p�Ѝ���7y�f��������Q�;��������T=��޷��om��$��5Leǈ`�6�lP��rM,#{��[�h�PvsP�+�s�������:<�͐̐f]��@�d6�8mߠ��L����W��)5Fr����D>����V��j\�#�{-���B���S�۷�{T��+�a$R,�#��`��������ǻ���R��^9ؙK4�V5�M"�N�f��엝��H��"�����`�X�wJ���
I�}3�d�E6_r����8�/�e�p>,�o�{�g�Lʆ�Ǟ��P�$iZ���t���h|
궀��U�_[�|�V{؏hvGi-�0a^7d!~��֖�P�jq�X¢�#Z%\B�N�Y	���&��x���eK��eZy�re٢Xe[t
]�Q��O������B��kG��@q���*���ء(�<���_#lA��q���o}�o^Df}�N 	D���Ky<�B�lv��%E(�f5��rD��G18sk��H4�P,�]@��������K��������7��I�Q��
�
�����%���b|��y�Hpv�튟�����"������h��\o�L-����%-�U@L�[�P��:B��''���Jy��1=Z�pH�M)k�{�yi5Ă�<��ߪv�w�@�hk�,�jb���&{dKه��ys�`
U-�J�F"��u����?A����UӪ�?g6�x8�h��.�M�`F���\�[d�L�XTd$J]7��v��Z���CB��Z��@���!+z ��Ge¿�f�*��u��
�B2k��w�~k��^Y�	��)���>IÞ?��uF���Њ	e��9�(d ���(]-�2��7]v�#�+�տ��	Z�~��M�Ξ��Hߩ>]/��W.��K�rM90�1��T�Ŕsy��?��t���}�:��ӫ��Xrĳ�{�+1�r#Є,s��j��s��6��h��M�{�L4����n� ow"�_�&�	h��C [l~.�k�v���d��p����E%:�`�o]�u*����U�����A�m���ͨ0, 0���҉M�����ݟ�tθ�eMn"�'��/�` �T��ؚ�'[�Z�?����8�0�@`['�7��u��Pq5�d|ݞ��.����� h�8;������%mX�D���YQnitB�܄�TM��y��{gS��XQj���|GvZ2V���jzkkۈ"6�E�LH�r�JٻDA+4/�X&�Q\"��V�ۂ��Π%�혙L`�eN����díD�R=}ջ�U'����]����iz?�z~��|hd�1ҝ�H�jj��k����8/������%Y92I����5 JP����1��eAw���q��IbӃd��#)�k��+�$���h�P����?d�E���k4�X9��8T�'TH�I��8 罬G�A��=}��s�c��.l���?��\�> @��nI�XJߘ�*@��N3Y�S�׶��D]4l���XQ���8�'���$�WQG��|rv�GRh�g�AMD栗J��ew18p$쑂�Q�d��2�v4�=��W�����G�d���蝇"H����׵���#Q9 ֱ|�%��r�W!�4�z�^�wh#����i�������p�h�-�_�(�nrJ{�5�H�C$I�5,;W�d���2����n��x)=�������2�*
@�QA�hUT�:@�"޼B������yz'���\��Z��怡ߋ���$���bW�]�*�7�ZM�}Mh��W�]Wc_
�*2cCJ��%��)x�~��]@<���{Cqf�Q�G�yX<��B��6��ĸM4l�.�����nB�ʑ��}���3�.���Yd��a�w�F۵�b��ۈ�� �p��/y�I��=]���fJs����C��f�w��k�J���>�]0B�4P��ø�ɧ\��Y��\�-���gٵ���?3�m�&y31�{�J��R�.��?i�w��bhS_؜���5n_�iԟ��2�k�+��<���9�2�m�	.�̭�^'_�.r&�B0P�zN3�lq��в�~��?BS~�NFe�����^4mj�m�`�;�O��x}����U��BRw}�-n��y��j�{�Zi�Ŏ�@���=<��4$z�x�x^�`M���Ig�-�ИШ9jt)*���yq��¯�'��$+�jA`���N2������Tm�d��J�6��ۅP7}	%c���h��+��!����T�'�`\\�p5$%R����M�oq����@ 4ץ`��Ҍ�#g�����`,�a������tф�&��X@��%���N��D�Q3\
?p[�P_zg�*�X�Uh�7�����6E�Xv�:����4�7�-3
���g�;�E��G�g�sʌ�,v�9e�,r��@����.��[�1�&ݛ���Z"?mp"U_�M�t�`�#�+3��=ψcX2w�{�o�����_�-�=��>�YB�޸x�|!�,��)��U1�}�TDjz��[��_Y�U�B4Vhu��D��Ou�t���`��&: !�+a�YL�	vS��щ�0����F������x�����-�������c�>��r��Rk�p+�\�5\��IP^弄�pp������ˆ:^�a���;iN��J�MCO�M�=rެ*l6kQ�������MCY�]@m���N/{�;�$�����Z������y}�1�T�~P�'���=�٣s�,�~�{8�%V2Eү�'7��q�\�s�r��=�%��2�K�B�E���,T�;���C_�o��4+J�3�^U��p7�BS�&wB����P�L��T�,i�ɯ5D5s�kJ�ߔ�>�dI_�B��(���&ȱd\�`��pb�^.��b`��Jց -�Σ �C�J��g�C���/���4؜���l������<i!����7�z� _g@���BL��b|Jt��"������!�ܧ�[��S�:g�!�5f7&�O^˦�>���EHM�w�Z��Ԩh�����a���]����Z��^�ۮFL�r���0�~��yS���,�x��g���s���/$�*�XZ��������!U�h8k�IX�=%.��P�I�98ξ���n��:^�򻌕;�+u�D�'�~�u����³݂�՘x�}�5������hd�P	tpk���g(�~�1-6��G �<~��ҟO5V��������A�W`�L"G�أ�:��y'�����a԰����jD�(�%$ٳ��:�Hc��N�� �YU5�
���Ǔ��o�y��J�?���W����73�[q��`�jތ�:��o��i���T�}�W�i����#VP���mF�<He���Q*h��2I"S�
]���  UƬ�� ҡϧ���#���
�� m3���6:TN�vk\�k_�_��M6#޲�>eP��(%B���O�ͫw�wAb��}d���s������w��B�p8��6K�=�ś�=��z���u0�� }=�ğ`�)�%�J\ĉq�'_li�B���`����k�;�{�H6�qe�Z�s�� i���Яtg=�Ճ�S3����;LQ�����$��p�G��Ǐ��M�.�[���,Y��DB���P?���g�j�J5��6��&�r�u.�i�d�n6@#�
����N��,�0�#FR3��C��D�0���H=������SNe���	��M�������(����tk����h�e����k��d%Rr��w�?{,^�����Sʕ�&!���r�'�ؑH���5�8#���BQ6+�X���c1<.&���؛,����ƬZP]!�V޳m�r�]3�ʟ|�}��z�W��qE�*=B��������~�(=¥n)�<�=��X'�ly�A[�~��l@�˞é���K	��<��TLNP�Ϊd��J$��>W=H�x��lڭJ�CT� ������T�fb��Rc������P��oF+f�8�g�.��cX!�����;tqq�o&�/B/�E�<OpD��'�E�V��lz���5��ȧ�$�9H��c[$��n�A�EF[��=����ؖ�[��L������x�X �M$��u�'z��ʥ����-��xތ�#]��s�������q�ZW��R�Sݠ���X�/V�jb*g&�jx���	�X[��5|��p��,oP@���O�9�J�b�~�jf�L�=��g���N-M	А�P'�J� �����Z 9��e2�ӹU]��x�V���JQٹKu��l���:������2sm�Ʌ�I�u
p����_�B��
؛$h�21#n+�0=��{^�z�jDd}>�wo�:���k�
���X˥������
W�5�l�3�%���?J?e��]7��9�){|�K�ڡ��M��N�W�G}�(���f>*P�t��2���˽��ؙ�����갚g[�����c���ʷ�5h{8r�BJ6�,�Ƣ	�6lfy��/�$�2u�\�d�W�tprBU���\������ `���u~$�U�/���{#+�#RH�%m���'����L,�T�w�ߪU([F{��-~��{�lO\��CbQ����i%Cۙ�ߖځ��'G²H:�����ͅ�;4���=-�@;�^��C�u9J1���ͫX��9,�1�O���6`ȝ-b��ˁ��`��\*���e���unE��E��ږ'"�a�q�`�(I�++�nL2�����I�vqE�������M!��]?�����Dsz�J�Td@M�*��0������t�u-��o����B�&qv�S�ogXs4��Ԝ������r*_R傭�<���EQm�g���A~G������Ȭ��k���90,�a������1`��{�"������7���l�WT��,g���R�x��9rvd�-u�X���?�B��{���S�`+�ҬG�X����s�����&l��_N�u�X��SBR`�C�㻵ĬM����OGB7b��a-?B���o�o���c���D"|���VFc+Wq�S�����������v�g��&�P��"�:V�k%��~ �X����b���i*�ә#�U��`r���^�R��@<���AO{�u�Nm��P@�IG����	WMq����Ɲ�Q�a��b���@h�Kk�+���B;���?���g(ܲ~���	�� ;��MJ_�dF;5�L;l+�썌1�8��'Ө��1��5`b8��6���@B;����T��*m8��X	Q�9d��8��5;޻�q�f}��r4��QY ���.�>�_�k�Δ�},~y�LS͐;H��� ��� ,��x���ΘM7�
���/ɫp�{��z�	�B�u�&\�ҷ2�(�`��5�4)�u�8�i}��(48�����V(�7&���D��(s-��CF �}����>�n�����%,ѥ�:� pu���+;ƛ$���3�<C��z��4LnL�(�C����B�I��OGTw��=��e8�1)*?�.k�4�⧎H�d��<��B5���d]�pd�2�ޅ?]e��Ǻ����!�yO�kt+2hh�-%�h�Dy��	��=Oڀ��g,����ЌҰ;�r�����QHXJ��Bdz�^��GK*��0e��E�HM��!�dz�D�C�8+݋0*OU{�w��$[�e�c�'�PC�cYz�B<
��Cy���M�{�w��Ty��,��W�QV�������d$
�^��IzG=�_A� o,x#%��X���1AT�Z�$��3̓[��SV�,��~�^z1G��J��� ��������
���W\n������C��R�Q�+1�@9ƴ���å r���&�<Ho�$��x(ɱE�&Fx����;i������9 [Ig�E�j�'��sb��v���m�Sf߀�e�1�v+&]�q�9?;�F����茒NnD�pl�ԉ�j�z�:����Zi&���Բ��Q�`wJ����'4z���T%�JC��Q>̣����1X|����Bg+��R��y�Nv�eIoWwO�:d.6�4���S|�P3�H��n':E�RPv�˕Oz���`� ��D��U܁7�kx�q��"}��޽3�����Xa��"��ץO�f^D�8�H	t��B���S�I�S�1�esdX��%��z�W��8�N�A�F���G��,���
`Vd}��{����~�����3T`a@���/�Kwi���ńqrk�:��}G���G�xh��w�0T�l��!���"����s��zW�gp6B�Q=c5��������Q�_B(ƣs��6~�KYKлL>L\&s žσ�պoW�,t����0E
H���W��Pn��$�����N��.��!�u� .���N\�q���
�8��S����i�	A�)-�ԥ&f�����E�`~־H%��v*�I[��{j̀�Fb�D�P���|6�����JL�M �G>�MO�YR�O�ޘzx8�RB=nY�rP����R�
'@�#G/3T�#�:�V��ِ4��Zk�I��K��y�eߎ�ѵ�X�� ��j�&����Lxg��C���p )��ܙ���~0��ޗy��e�H|6#�j�"渥����1�Y�&ѩ�~f؇U�y����"5��2 M��gO,�x��(}�fr9ÿ��ڶ��O���`b�[��k@ ���1��=V�qq�f�Gt�}��8�`�QDp��򖦜:�&7��	�-x^k\Ep�x9Ja�w�I��źm&�5*N~$�*�c��������u�֏�Z�	(��P�_����w��_����#�a3:`Sw�d���"�����sHf���w�'͑�OX&�_u��ڕ�\êS���׈+�2O����g�ԗ�-��T0%v�G
�
�T�±RaC�5��R󁅝����QPZ7������I���>�1�� P�0i��h�Ʊ�3���k7n��Խ�H�`�B4��j3���2ł�]���r�g�w�i1Z�t�B���E���@��,-�Ho�)Qc�r: ����jQ5tJ���#g
Y�������x�x����N*˓6�	�1&M��RoX3$�"K�S�����~Ŷ�����eR&�d�G B�Q�U�0������f���J�����zS�>7�h��,��E+�O���Fύ��Fb�&�v�$cV<�X�-�`I��(!��\z$�u鯸�q��)�m����ĞE����Z�"�ˡ��Z���#�iӹTE6��*��.	]z5x�����i�Z�@`�*�Nn�I��}�����2��!@�"��63��9�U�}�̵�$_�B������nV���#'�6\� mi+&γ�^�s߂.���B0�T�➬������Z��B��LvZJ��e����HElf�҃��o��ZSMzF�a �JN]T H�O�������^$��J�ܯ�`
�Z����8m��k�F␒f�0c�[���
��Y�TX�§q���~ݱ�܎]e�ѱ��
��Nd��˗�`r��v@q�����ڇ.K�Ь�}3.��*Nq{��!O5fP�U'L�|��"��ƨ`%[�U���;.E_�����%N�+�9(	�b��=��`T�.�"������d�����"Ȣ�"CjoS���^e�7����_&e_�-�5�.�6��h4c=��N���O�Ȭ����Ԛa���+���1���%�X���X%FZ�5���&���SD��I��p���;�4(�u��=�>[��1���M�}�KQ*u@c��َ̢�F@��-"Cv�5��h:V��-JO�T������5e����]p1{7p�C�0C20��·	"b�����BS_��!G�Vy"� .�����	-6ue�^`�:�{0��3�����{ >�vxo('[O6X������)�ʃBX7$Ҩc��PF|��)���5�����i�S�,�%V��#<3Ӊ]���m?�k�u��=)&�����4����)+�J�łi��/���Cg#���z[��h��j{]a�E@7Qˏ�!ӡ�q4��_xB��E˛`�if�=mO�^�b�oP�R*2�jc+a
g�zeV2:��o��q��5ek례��#�{S����V��0�O����C�[���̿]��b�]2��!e	�g-G���?h/Kj� }�!U��ۡ����`C�i?�sK7��--�n�� 
�u���K+0�N9fiJ9�̡�eq=e�k�y��(bܷY?��1��L������*��U�$�A	�'4o@~~Z�r~�٠�2#�(�5P�Xr�F�\�[m_`��Yn�Ω}O�a�� ��n��uX�A��1�\�gs�Ǘo���V���4貢�8�%�:F[,��x��+�O��Zi�T=��l>�d�x���yr6�R��	��Qwk�:�j��˃F���|�f�am�,q��\��/3*��f��l��� �7BR>���S�,������N|�DI�wr�������i䮺�x��'�	� ���l�i맄�5�G�{���aR�/g�5����5��Jps���-�7������}�Å�l0�F�Ae��'�sTR��p��ѷ$�Ƃ�_���?���(�}�?�!ف�' ��]�p���K�7��<�j�u����T�R�ijgk�B47[��hwc�u������P�}��Ɠ�vl�-�1�T�r���π�ƀ&�ٌd���H�,�";��s�o̗��vn0����/8�d���(�9P�u�k�HT�5{I�!:��r}o������ _�,��^٪$�|7�D�8�1�2�|�^L�ņ©ޖ3��tUu��z�bb0?�eO��G9ʥ�%�F�y-}�ڳ�V?J��&؆g���^�b�����������6D�k�� ��?�&�?�I&у��D��m�W��S�و+`��ثT^��xU}��D��\�D��]j��Q���myztRw/�$h���� )����i�J��2$ ��uI��1h�#f��j���\�����b�+�0^�/JT������,�(�R)��ނ��[N�Nζ�B��o�x���ƚ1�	�51A�E�����#Upz;�n��_!�[��D�U�!j�0�ëjD2�;>SQ$Yr)��[P ��6j�o%%�ϛ�,�����5j���a�t+�R��@aғ�}y� ������ƫ�>��k�>� o �R�D^�=Na���7-
!���W�>����Ϭ�X4�!�6E� 9��C��" ���dN�a�)\�Y��}�|˧O&o,���6��D�N\w��}���۲��m�GG?��L;�l;>k2nQ���,��8}ݼ��y?U^8%�ƌ;�ĶqV�f��q����NQ zc{��L���+-��������X���`���%�bB�٨�nX��{�kި R�Ș�T\�[-�I[�SkMG&�.�z�7��m���� =��x�q�����"�J�p��L�$�4��!|