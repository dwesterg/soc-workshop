��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:Z��� �B5�&��jIK�0���װ���p�%��1�
�+\�w&;����W�bx�>��?�%��D��.�"l|�T�0ӷ�����%~��+� �h�o�Gf�{<3+�8����]|���*�C�7���C����@�LB�!f`��@��h���5Ȉ\��o�����y��ԛ�ͷM����h�I�}~>��J��ByD�l���Hx�����Ln��q�w�e#YW�����S(���3H�1�f�
h<���LI�;��Bӽ]�BI�gks�]�c�^}�ZQI���x3z���7ڏ$Vݪ�);�zAnKR>hY�S��8��Prؑ������%	O8�i��g��UK�Z:�y������}��{�%���/j��D��x�Rfs�4����֚="�6���Si��7}#�'{�4sޢ�ɯx�M�r�8�@w�k
���P��c+\l��|�C�`-�2jnBHj"�0���]	d`���{�D6Ps��3J/�U�����%1i����6	Z����Ժy���ϭ��/�31��q�RӿaD��X��K.}q�F z�#�i��J�)�:�C��>���D�C'0�7
��v���>�Z�mʺg��x�T%�/��g���.#��o���e�y�&��{صeO5׃!�[��U8Ј���ڶ���&�g��Q��|'�7��ݳ�.#��έn����ч�Գ�8d��*��<j	t�/-�K^l�}"�=Э�A`i�G��_s�9Wއ\��b9��z%�6��|
�L���!_�j��@FT��9ɗJe]��rb�fp:���%��5s��T��'���X3n�7����.�O5���V���/�������
�%i��*�6@Kނd��f'�F#D?�ҖhH��E�ꌣ�5�U=8k��� ���mPo'�Mw�}%㗯��R6��>V*=	N9�fR��g�o�Sc�I3<ǥ�[�� �׾j�5E��~Q��ܞ�1Fѕ@�al06������7��k�ޱ�̾2�ч����v*w�Q9�UZ�%���2O6�Z�T)�G0�d����/׻�+�.Bnu��k8���`h����mz��e�}�������Z�q,��sed\����x�}IX�L/p��(4R���o��`!OG4 �@m����zO���:%��X��������Q���'zΥ:��y3�`�M���w-���Y��NW���H��MfD�[��e4����l�����}�zL��e�Lт�q�����a��?Q�a���]����p�y�n��N�O�ʋ��H�vn����<AM�p&���hs9܎ۑ�B��3Q�^��~R,$�A� ^4j�G�J�騟��գ��#�� "h ����6�^�J�2f�ɛt�
V3T�+���@���n��!�z
d�T�G�7nEo�竹����a[��Ѓ�7u�ɶ�nٽ4N��C�)�,����{^�Z����_��r�h{�>֫����x�;`�co�f�-ܡ)�ަmĪ�<��=��e���=���]!�G]��ܰ��x��^ZǑ}�%�!Y��=��Sj�W_e��#���/4��l��F��9��0��ld �6֩ݝ��D>R��Y�a��I�T��0��j ȉ�|����uٛ6|fV7�=�Xo�"8H�cyy&���|6�*0L]ƊG7x{���|��&���	L��N	�\��V��@�8B�t��`Q+s,��7��O��p<�����lޔ�"�0Dv"����hW�K��h�p��4����R�"���M�u��)1�29������c!~��(9���4d����bsWD�p��#$Cx���dp{*y뺠N;����L��~m�N��
��R�y��}L��	{#)\�_ݲ���W�dI�l=��F��q�[�p.��t� ����Ӫ����U�_(�Ȏ��F��@T%�/�|o�m>R���c�T��ﴸ���kC����f��� eY��Ӱ�J�aϏ��qh<���9������3ӍvF���������\��B�PIj�
���I�'H\�[�-2b��Pj�	��6ŗ��դuk�8<���WnB"Y�R��y.�#�e �N��]p,�7��U���\�i�)��:��큐��~�Y����#���UC�Y'��v�AB;h�nM�aIx G���<'�7�f�j����$��֮N��l��~�JJr!����\�Rz�Ԃ��R�B:e:ֹ��Xv��])2��t$
g��N�T�L8�q/ݶ,�d�u'_��׭����݅ɺ�׿�A�G4U	4���F3�
��vE�=lĆ�����n�Ai[��r��]�Bo����6H�vC�ǣ'H����6�}2ww�}9��x)� 2���@��,b<fv��j�rM�N�]��Z�o��P䞧+����,�&>�Z�{0������r�p�P7�s촀{��y����*�d7661������l����m�N~4rc����*�4i��0����A�)�]�zӞq�B�TXލ��֢�'c}f/�����z���Zv>A S�Ab�R7���nY��bjA�\T�L��}��,�]dݘ�5TeuY��N�� 9����vc�=��W������ƞ�O=D��<G`�*�/V�٬�M�y��(�L��/=��~v�˛�Q�e�C�@R$����Ͻ�������-�EsC3��!�?7�d0�;�<��yG煂�4 ��D ���N[R�H���-9G��4��F�6np���v�b0�t�k��M\ѡNk��j�h����O��|O_N>o�@�ܕ�,&�,�Ґ�!�6u���<*4I���|�s���&Y{R�/ͅ���~��C'΋#�#'Q<'>6�3ׇ)u� 
ZIxFJ�����М4�A��u�X���qb�Bp}Pj� 2ԩ��2�<����p���)�}R��[r�n�˹��q7��p���0>��׺�{������Х�S1y�vI4������Q0D���5Ll���4L�V����ľ�0X�L%�u�s�����{�~߭q�#�e����rW�9k��]]~�
�c�ď��,�W2�� ��0S�>�N�6S�$��;�g���(#Z$F[�����u �tj���Y�����{C��e��O *�~�����5�v"����R�}���7h�,�@�y�A�"��(��>�{*^�J�bZ�P�}�F���O����8��QsZ��/����b��T��s�X7f|��i��*��s��zMs��R��t:��{ w��#]{���'"��nB!OZ��box�w^�-�4c�)nO��M��1n�L(�;��B�d������͵ e�A�]�r<���SU��F�sq��4���.�ܑ)L7�,�{BY7j�N�l�KΖ��A�������4�2�2���_]}�B�i�ԐC
����S}i�J�h���V���z������ܦR\tƞ�_7�]�*j�4�㍉�	t��boFˤE���0m�li�%I��I������K�H�u�\1\5�)���3��b<�� ��l�Rk*'����y���$��N�ؖK�O�
����4[��O��&|Q,�k@__�Ru��d�,W��^��3ּ+����3t57�]�1�á��f��n�Q���?����+�+�
釪��$~89�'�a�W�0\Do����^�L��`!��
e�=�[0���W�F��)J
HL������kJ^<uA�( 1�1�,�K�ܳ+���n�$B���sH �E6��!�n�3Et.����[u؞�_�O6�D�q�Ý� ��[���.����6�J� ���i�"�1��]��-���|��4��D ����l]�]w|j@_]|���h��$��o���������Z�)}��'��dS�t0ƶ_�w�j�s���Rn>��q�!~6a��Eűtkd�����_���B+Y��焠\~S�'8����vK�,J?��5�����Ԓ����99���3\�