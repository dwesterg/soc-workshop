��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ�wL#������8�4sFx�� yo�"��ş��gÛY���"��G]�z��`XǙ�8vm	��r�K��%f5���	���!y�e��{Z��S��)�T��%�RMi+������l��(��Ё���(�J�e�� �T�E��6���m2Q��<�h^�v�m!-�ޓ#��p���uti��z��8��3�Xv�$�0�L�b
���\]���=Q�������oo��k �W����*D���W�H�t�B8g�k?N�O\Gj��P��<�C��H�����8��X��b�����K�EϬ�C�.���^::�7!o|���{�=�o�T����O�)�^h�k���Ie�G��K�$�B �g�9�=���މ�S�n�:Yr��|J���9��ί�Ud��ݞ=�貿��&6X┣8[�	ڍ�y/�>ێ���8�{X@\N`�#�����b�D�I��KH�a�t���/o�I\��\����˓�؅��Xut��=��܈6(�Ve xv�,��J�I�����r�b2�~~kBJ�œ�7��AA���
Jj�?NJ��dG��\�j@�R��͆��Y���vO��`�QZ�,	F �[��Ҧ��̖��)tQ��ۺ*vO���%^5c�[�0���>\��y���vb��B��ʎ��E�&m]��`��(v�����%k6O�W�Akj�10"�r%�k�R�B���ƪ�I=��ҕ���D��p�eSC  c���+��5�ݔ*��_�rl93��!�mb9��l=ò:����`$%q>��l1���㑵쮙m�o��J�֯�d
97�B�!|IӔrf�M|İ��q�S�bJb�zItEZ�ԙQ݅v#��%'Pҧ�S�PN݃����1(�v��S�h���_�CNQ *��}��d9U�iH��#��Ȗos��ꤘB��Q	ڕ����ch��ܿ�a-��B��:�|\ARO]J:F�M�j V?I�!J2	�|1����6j���/�;������e�_T0�CT>x�?C���k�mWɀ$�[(y����'M�C�N�.&v�(�pϮ�	$���_4�k5+YO]m��z���2#P�q�Qض�l{��g����y�k�O�j�d|B�P�S���A�}�M 
�oH����1�E$����ʠ��+A���by�- �nWH��gҊe�:����}�1��&���y�^���q�����*�.X�F���:SXh�+��E�j>/3��`ѳvo�$��x�r�i�!�U>���x`����Ѩp�E�Y��c����*	.	�-&o3��I�59�3��k�e��W(Ռ����[hC�苠B��8���/�������y��������ӽ�C�ǟe7o�z��_i>B�#׺b-�݋cm��j�'}[��up��z�R'`�I~��Bj����	��EO"��re#U������S�%� Қ�X꛺P&z��s��هſ'%cѥ�@��4��Q�*���~z[g�󖁸��360L�/C~��Ҋ��e)E��)�@PR��L+�g1�|}�c�*������,���}���z���qQ��|�F@�CM�&E�K�(WwP��F!�����A�%�B�5�B=��ēQ~J]�x�/P�]V�_��5�"k�A0n&�S��+������S]-!���й\�\���$�@>�W��r�%�_'|w��*��X�3'�[¥X �G7� �_�~�,-���1�"�.�wJ�ܧTW.l�S�tk�-���z�3)�������8fkG
Xю�Q"����������� ���PU��F̝K/8�*��2U��T�f�[ݟ�`�C��n��?�73}����i$e�:'�t=��3�k�#��>��<�G#O܀m4i�BY�YB׎qK?�P�l��,���=�4edYZ��w�?q�����'n���g ��a���c;qSyE�������
�P�(�2L����휔��j������ݒ?S��K��-!��M�J�)��Y����n�D����V���5B��<��	ENI��5��R��.��4-i�&(]F�;��-m����"B����	껄H�N��S8��e=�8?���7�"��2uɕ	�!��_���|�;_�>_��jyD�(md�ND�L�EOb�|��JnLDY��+H����E&�0�>TH�`�9�ϕ�{SL�������diZ㟚�����*�lQ�~/[��$�J��F�Dlnŭ���v�Ғ���#���&w!�0�d����<Р��L9)J-� �������c6)�/��7y�.����6�\	�Ne�_��s�-2���8���0'%�,��o�z� }�$dJcw]ۘ��)�Tqz-a��yh~��hYi��%����C�.�R�5E�R
�$A[3z�gg+I8R:��mAZ@�<��(���gl�*���77L0¥�̧CI���&���&b?�\���zH�� %�-�H�[���-���Yp�ٓ~�§�]�Qs�����aLr�� Γ�QL	�`_E�:�R��D����RʏS�+�ɢc�΅+l�ȴ����Oȁv"VY�F�j��z��f<G�/��y	s&��f�`6t�Yy~��<�>v��nDĨ�/%1D�ȟ�m����PņfR��O��o{��s6KF~������V�._xz��ح=Q�T�"X���)Ρ�,q�ȯ����I��N�5�,
�e��N5-�K�F`��������iu[2�F���L�lA��R�s 	tb�$.Pח���������D�~���R+��M�vR�7���/A��,�Z�L7~|	d؄f #V&���х�+�	ۡ��/�c�;,�t��JI���5{.����t��F~e0�"S��g`��҂�?ɠ���ѺNx $�[���Q�BZ�ˡl+X}��0w��M��՚�8ݚKeJ�7m�o����[��[�C�����ڋ蕧�DnOp%�L��uB���I�����a%P��C����]��G]uӃ���y�<���IyR�,��!|�̱U����M��='q�b�b��t�"wWNlq|�k9���gJ��T�r xh4\��P�\"V%!�k�a[���K���bv�=3ai�g�(az�&�o������VQ����sx����Bq����Ѓ�N��Vب�kH5��j0�`�������Һ? & ���|��@��S�4G�.m�mc�g�Z�Ί�_�M#����F� ,	�^�6�Zb�,�Z�.�c5	k����ȗ��to*/k%����w�eb���ٍ~|��[���'����V��*��������x�*�rb���|b}$��"?���I�	_t�ޛ�Z)�k�/���0f����G�1��0�^�X��m��o�E�jE�7�ۣ���*��\�x<�{'q(������cR�b���ZU�#��E�[����ɗ]�)�{^i13,Qm��m�lV��w��:)��e,b�
;�d�o2-Ѻ̾��0;�5��:��҂,���nxH��^?�s����O�t�`+ر�� �>b�eɫcx�P�����B���NvKg�*�
2NN!9<uE89�fkIg�Ya��MH=��=��X��Ժ�C�/De9���`���ǋa�KO�݇J�����|; �%CL��#L�D���=q��'�XKG�9b`�'��ǻ��P����=�=����_O,��E<285�	U�x@Z�i�e�gx׻ pAĒ��*���B����