��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t����z�2w���*ٓ�����y]����p$��o����:r�RwN�ӻ��i{�N�k�wɣ�i���Ýa�3�be���+�kM����Ò��A��L��C1�Ý^^?C�R�/��Տ���fqj���O
��ÿא�Q��-��C�R�P��"�(�	��a�-�u����Y3�H�������� �|Fg������(��#2�2e
9����562k�jܝ����QjM �2�݁ ��7)Y�%�<��������/�|����Q^�k�l�kl�e?tr��n�)~z�ɴ�J�!a`��!�	�\��k�zqǌ_QL|���1{��>�8x�.��zz��u��F���5�E�^�V:�y�*���q���k�Yv5�I]W)�~rps쩭M�$�AC�^�D�ci��C뻠��n9���ZO�x�Qr�"���t�7�0o�5YED8ܟ�PR���?�Q����|��$f}jw��*P�ub�8t��I�FM�-k8���{{))۾GDs0���<3o��6�x|Ev��v(`ge��s���e{XU�\��yz!-�aݙ��wPS+U�QǠ-��ŗ�]��8-2F��{�H��v�Y���e���y���tJ�jCQ��J�c��5���	[���(IHd�-Kp��]-�J�E�C���9U�1%��Uo^�bX���|����@<�k��lv�t%č:����-M��@�j��݇��r[��&h��h���59�ؿ�����:�;P��9',��(�S���褍�. ��b5���,,M,V���_�u�����z�>�# �|����^OԲ�X���(bq�=��WD����Q�O������=�G����A�E�ha�������D��lU�[U{�#Y�����/B�6 1��Li#n��j�vm���L��\����G��6���I�y�|m���S�U9ȝ��@�I�S2�����E�X'v�^fd�&�a�b�(�߃kxFH�\t&-��֫��^{��$��]i�	\+��3h�(�F+�,��~oxH�Z�j��cR*1��p����l��Y���6@MCW��^�~C1�%�,A4$kx� �A�W��IK�t��(rWK [�[P�d����U���,�h0Ǧ�����) �C�Q��-��0I
]��#���:4�}^�(��X�u)D�������i���#�]F�\s�d����w�"���N�(�ٝv���(�'��'���nī�'aM�:����Z]g&��>~���\0m=C�š/����}�˥S5%�a�,s��L@O��i�G��j�2���=�C��ZNբ؏W������>:��n4�3h��6��oE�F���Q�Qmv��$����WT�1ZK5��"l�EWu<�]�7z�zO��G� �]��ђ�G��87e�������mɥǔ�L��qkVkt�l���t�*�d���!����n���ܫ�7r^���lP�*�X.��e�>/X���8^NM�1Gѝ�C�� D!Ϟ��e��c���j'������)It��c(e��p"F%�rC�7��jY{J�R��ր�̱�\a�AL%������V3�!��0��bՒ��liY�B���ͦ;?�Je��W���g$~٤��MݝKҺ��S��ξaa���1�t�Q&�/�w�xw��/�.�Bh`�̘�ǁ3��&3�X��;`@���&b-u_��%X�83&F��y�;W��;���d^Y%����%�Q4�2e�$�T෿��/sn���i�v4�4�7�왮��L/��KLA!Z���s���MN��{������7hv�KntZ����]��|��
�9�5��,s�X\[��:�||2����iB�����=@����2��t��$hѼ~���W"y	����̤~l�o]�s�U�PB���W��h��;vt���? 3���QY���m�nsXkt��k���;W�s��?��1�/#���ަ�õ��}�
�Q�+_���4��
H7���a���PZyS)CPE�����ߨ������dV���IU�4Rm`�If���r7�#���r`��6�D�c�p����4�J/Ӫ>nl�'�%����&�-e��!��wMN����2�}��U7��Q��L��x=��O��^7ѝ 	�)|;'ں��29�u6ָ� ����ss�U4��0O�@x�d���;���c�vk�1�<�'$��Uʴ�h
}E�)�Z0�6d���PD4'�]�<�zf�a�	�]?�CRj�JA0.b��/�s�Y���@����S��҆�>�ձ��+QQx�t��[�$�Xp���M|,���`�ÚK�9��N�����Gخ%�sv��Q��b,ϐ�S�b���C�b��n����^np:�����XS�[�BeI�r=�`�a&����z��VV���e@hKE�s�%q�Ŋ>�!�N�ם��e�G�,/�4�� l{H26F�"�$�CX��N��T��OG�G���.�GG��)��s���9�p0W�gv�v�jD�@pj	�^�a-_�}R�恹C����.��z��a�GBj�L"5X3A��=��{�W����QF<�t-���{4|�l]�����:�R?���/�h�.t����8��vdk^ϊ�^�%%ך{Db�C&�މ����7���l�<>�E��,�������)�k�Z����A�"�x�U�������Gu�!���C�%�h����J��H���T�iZ�n07E� �u���e��-5|�1�v7���ţ_(�!�TV;�Kě��9���WM�d���E�ɶ6����:�T3>Qz^�%(��i_��!t]��;���*���\���{6�<�HU�P�z[�?i]1q��K3ۃ��t}���L~R �y��c%o@�r?i�M���2�1/�o��1�����l�OF	k��<GgBxM�JR)KMj�08<�oȟ�	��6e�nAT-��A�V����[�R���3fԪ�"����[�'������o��3��r4���$ǶB�Gxj���Yg�<��#fgb���?w�W(�g��BmBB����k([B扩��O�l��U%ĵ�;q尶�U<S�O�v���7�{�Z<����o�y���F&`���0W�M{�g�(D4f[�%o���|Q�+�CH��4�>lF�� ~\i�^B����r�sз5�2xv�� ?o�>6Zt{��\鲌a��4��i�MN'zb��N���ŗ��l�3:B�^`K�C���m���r-�ML��f4��>K�]��4�=�$rK�;�X���n��%� �v�C�{����_�캣+�b}�kTv+Y�( �-��0 ��LC�-%c�zG;Ē��V���;��#����i`WwT�|A���:�,s�M�Z��`�	�&���*,��9�a3�����D�:0��D#�;I\���-�������Ӌ��Dr�K�9��΅+�� ܈��g�~��rf;���Zu�� �Օ��uj�M@��>�iU����
�N��.�/�-jⵃ�˥ՎV�uh9�ū�[�[g�Ѱ��L^�����8m�&��@d8�����7B[?��/>h�X��"�2C>�����-�A��@t�炤?�����Gc6#ĸ&��>Q{ět�N�:G�`[���l2m�k�Pp���_�N-{Z��A�,zk�y\O�|f������Ğ�o�X`0���d�B7DW/���
]t^(����df���P^�Mp��솿l35������T�M%����u�pHdc�i��Dg�^���v�P߃�4x:cI���
��+k0�l����ǚй�L�!	�W��*'����{��)[����2��WZ��j��Rp9[}�X�\(�}�g��D~��r#S/��"�m¹ iu OuoB4E�O,H���+���|���0}��pi<��/Q����S�}��0��E�$%OT*�������9>c�n�t�9v\C���K�6\�[�?k{{deȮ��n ���p�rÈ����/���F_S�5��vD��Rޢ��������Ca-C��N�p�F-n�5�g�. ����s��WF�?�i"-��X
�O���(��`�|�Y�B�XHu͜��)�� 
�kSSu��z�9/o�ݘz+�`���.x�z^#X*n�R^�!���� 
��kXxP^���J���J�P���5�S]dLi��c��^� ?���I�n�m��k����FS&��_":�p%�y�)n���b�l�{�u'��+f�|��u.��/��¹u��u��>7�a9��T�:�k���3خ�s�ϭ���r���
�/U�_B�$����F����ş�-�(�R�ڄ�����!A7�[�L�����l��	�
Ȋ��}5��tȉ���� ,*��JA%2���MrofO+�*��\���$��?��|6�݂�t�?����q�F��l��	�g�fG<Ǭ��Ԅ�o8��[�ã���u�N����5	M�J����.�P�O��/'��O���Q���[v�_.����/XU�h"�b!���VW����HT]nC�r|�Q��?i9]P�������2�;�)(S�����/{AN,i�Q_�^���
{��(IX��U CXс�k+1.�O�}��'x4�'[�.ˤ�>�m4I�nH�M:�����&^�����j��^\/,S���F�l��(Uo�hmuo���4��+��+�HKG�^������#�`�*���ho'� ��^�����qZ'�i*(X6���eԚ�PK�ߎ�A;���ޫ�
�h��|ꢃ?��6B�|�>�s ��,&�p�K�2��c�������ٖ>ƭxPN8�����+�JAZ� oޚ�
v�H�ո��8�����O#��вV��q��R�=}A��/2�x�E1�ƛ��'nrv�hǎ���ɻ�ŦՒ�hf����!&7ۖ�� �p���*� e[YqȊf ��g��WFe�׊�js�u��B�8���l�M<�9�C��l%|'�CQ�*��K�m >
L|�߅ݏ�!e�r8�iAC�ɑ�]�_N�\֪?Q rB�h�>l?�sh&�43�X�_4�ԩ�N�5�l��5���������)�Q5g4',�RG~�#M^���P2Q7����]��- q��(�Q���-�n�b��c�U6v.�xǗ�����(�@�叫ϔ<J�g�y.^3£g;�)�V��d'��Y��J�⹠WL���s�����7��u!�i����<��ȋ�֠�Kp�k_�F�D#3h�|��N�8)u��p��^�ft�-�����ޏ��c	A�%�Rv�� #r�����N��$D;SE)���,K�o`��r�Ԧ��юj�9�������l�8�*,{�X����r�K���Y���> �#$�d^�<Yi�+K�)�k!k��)Ǹro�D�!��|؎ �|����b`<���A��r 4�9T��(ά6Ƈ�~����0me�ٓ{Q(�J��i�9Z��.ذM�p�L���)2Y����\6Sw���W�p�;&�0Lk�$� }�����	K��C���Qb8�7t��N@тfߐT�������r��w�	>�L�+h?g���F�k��|���˘D�#c�be�VF��։��Y���J8l�(�-�qT�I�K�bq�$!����{u��K���^\�+'϶��=/�2����bE��4��EE�#��G������f3ǧ�Z��o����nI�}:��CP�%����5�OcL��*�M�F�p�ȱj����%.�z�����p���M�[̶�w�Et�Уt�g�%,�辇2�K+-Ï� �b�(�.h�'c�\5��x?���Tx��b����>��Y��zBM�d��ƹd�لWB��Z���-���&�у8 �@��o��]�|��d����t�z��m�D����l�D	�ѣѕt�×��ٹ��I�y��ڻ��;�je�ä�B��]ן	��UD\!����PI/;䷇w�f����p;��w��\l�H8��! ��.�dEA�EQn�����`!��>m4BUIId����
%6n�B/�����ތ���|Z��/T�~B�*?� Cg�^�F�#]�j����E�}��wa��/�	��9d����CR��-/`�I
� ��몗�ۢ+_{��#L	�$�� 
�4��3�!-��P�@�+��m�?n�j�BcYu8u���>_��.��{
��"U��*�%5�T��mA���7�>f��`����aL&�`Mg��dӇu��`�A��u�q��g Z�n7Q�K� ht�z��v*E�/��.C�[ٖԘ�}׮����O����	S9e�����	�E��iO/�J���(\PG)�5�h�p�W�����Y�3:
�hf/W�&
��8�R���(����Ad^r؟/�+S �g։hK��/��[z4��>���	X�S�V̗�p�����e�އ�Af�a�u��ţc?z�P)��Ez�@��R~L���^��1��X(&L��^�N~�ȴ���O0�8Jvei7gg\\ȜË�BF��>�[}����9�WS��d=�>��$v,9B�d;�!��]׽,���9�-����c�<GNhWr�o�Y
�q���<}���U���1b��Z��w�õЩ�\�;$��mM�����Q�I@�L�7�ܡ1g��:#e[��n���c;�����[��R�aʡQy͝uS�5B�I;�5Wg��&�Т�jԎ�!&~:��P��(>8W��F���Ђ����މ�.����oMs�.i}7Z^"��FOв[Jzt�a(��A�(�����;��~�29��-�|,,�,��Q���R5�����r{�yF�! �P�9$T��<)�Kq�D֥T�Ƶn��G���&�P�(6|B r��%���!�z��QL�����Eȡ���ċ[|�{���t^���2D��׌�)��������[���I͡8�Եy��L�uɡc=Oz���",���"M�kw|�0�׽�v,겡�S�zUK� ��C���)�**^�CL_k$�*SI�s���U	h��e{oqG8�-"��T(5$��t7||�$;M��5_Ж@[a��y������9�x&fl�u�v�A)=�:��mC�(�G�s!=`�A���gA��K˼݆�AĕG�K&p�;$/�mНMƲ�,��߮o��T��Pk�с'c���:�J!˳�V�Q|��F;� D����~hH�!zf��)�;vf��a��6��ې������;��K��F��p724��^�N;�]P~)Mt��F��kԷB����{�����'�أqt~.�C!�vb�}��,.*9�
	�f~]$�Ĵ��$��Y��"�h�Ky�g/��d����Q	/��G6m����� ����9��Q����6�L2*O��9�������֗9��HL��z��N�&��(�P7JQ&�eK]�&�L��3����<�E]�<��^�gӡ��8Ga1�:����~�5�/ĴDw�@~�>=y��Y�x��i0�Lo�c}���	=��y6K*͡XkZ�zx����
#�\�	������ ��/w�ia?������-�JH)����Q�#Q�P@�.���mm�b��|���ʻV���9�L,"���L*��G#�3sf�ML�M��,���t�D���#ܭ�%�H��wh-��F�q�
��eO	��N���w[B,}��+=��O__:���+� D{����ΐYg@��� &k��D{��#2+�
�J�J������F�E���}E�
���GڜW����̫Yb�z�_E�t�z�:���36Q��U#=��,([I���q�MX?ӼO:R �9g#y�Y;Z����W�1��kFs� ����O���5Wu�����'�bq��v[*��a���,��idX�	�j��T�>�"�8��6�U��*�M�1�7�R�
U�<�eš�MѶ��!�~՗�:�~�\_��<gE�ٳ�5�%	�ns!�g�S� ��VL8:e�'��^S�	�w�Vס0A0@��;}��no�g8�	����|�����"��4zi�ɖ|��;��D��6�"8� ?��V����޼M?�esZ�O٩��u�b��P��Î�CDS�2>�	C�x��(��M8 ��ߙ���t��!'�-i'�B���8<�̡�F��󼚞Y��z��N��#1��|\�S{�S��ޟd��x#q2.���z3�ui˓�6U�`����E|y�H������!@W�?����;�O=4S)�N�,z��]���aJ�G&�G7m�Z!�M��X��H����X�3��ҋ8��¸����6�,W�K��(�,�-c:�ꙃ��+�*�)v]|�a٦�M� �tv�>�ƚ�$�a�b��X��!b�.^e&bŵ�'=��pY��(�%���c�DS��A�}��#lH�yWH(:R[[.�b���un��ցϨB�h�z(v���gq2�?o'�dZ��A���y�K2o���Mv���W-ή���g�RM��1��t���i]p�ޓ�n��t���Cd���xE)�#���%[A
R�i�N��7��.}Zz5o�-��b�T�	e��3�	h�x�TPe��.�`%��+t���#�8�S����U߃�d ��'	�_��O����
)�L.�}��|��D�wԡ?s�\���h>پ0@&QA�^���|fI}��F��օ	e)�+�ݮ�Ue,��� 6���ͱɺ��P��Q$���a$�+5"Lk T��S�5^�!.����FpP���ff��ڰ�v�&�a8�yW��,a9�3�J�'������������V�#%�W����c��z�C���#W�&�wx]~fr`�g�Q$q|�;}�����N� A�0|����ժ���Xsi�8���e�w2���Br�8�f��#ڋ�Ӵ3hH5Cl?9zF�<��!
@�R���/�,�gh���G�ْ�4+���Z4�}����s�I:G���&}V���)�֍(\(���f����W?p��Q!h�0��n�5���u��T���i���V4g��-�:��<���[gs�m�M�Fm��K�W�Q�
>�~s:)V%� ӊ��"�џ�l�֪YeZ4KQ�`7����T�}��|�Z��0?��d5�@�xB��|��y�T-X�d�zQ�ѯ9��-5���8�ju�a��~�=JN<�wxu>8�6-�|�[4�]�����o�q��7fO+=<��H��ѐa�q��*ǈ���&$�'4����.�|��A�"p-�-��/��U���.��y��!�[�����!��Q��� lh>�S��G&�f8��#J�xc`�u��q�]���W�,?:O f��I�P�h�IV^<�[1��{�G�+�qS��!Gv_���v���v���Д�b��dӍ$��g���Dd��o�wb��/yO��$���`���	k��d8S6M����[C�A���H_k���Q��� ܻ֗�� o�)	t�V�.Yʀ.��������貒�޼+��ǼUo/]�զ�'ܺ-�|%�V��y���>������D
M��d�"2Q�β�����t�E��!�N.��7��~ ʐ�n�߯E6�M&���]��K+0u�	�b]�,9���D�$)�� �=��?v���uU��ԣ�)�е���N�S�L0�t\�o<��S``>vd�U�v<�1$l9�ܺ�׻�aXh��sZ`�E˻���I	y�R߳ ?�/��@oBҳ�$Ħr7���fϟ��W�B@�3��&{�Um�KS�{�z�M6.�O�f��������/�Y�Exh���^��H`�\u�m�xG��Tu*u^#q	�*��"\��[���\��,u=����/2z5@��k�z�	,����S*�[{F���Z��P�.W�І��\?	��gh��A��~n�����\������.M�k"�y㉭2N}:��t3��o�F0ii��rD�Yε#�V��ʙ��Ig��]k/�!�DzK���m��}[�!��7��W�#]�"�����IL�5
��b�>���Ua����)�v��)�?�h�l��d���.�[�D�	ڱf��QzSTN�{1��Zm�{���������C%9����]F��Χ�zJ|���L�pܼJ:{sF����� 'ǊT�A�zs�짲�	J<�n��#2��#ϧ_fߧ��|F?�׸��9�������g��&>�!P��8���G4ۣt�{a�2�$s��p�$?�V�"�Z`R�X�.=G�(��q�7��P��m*+O���Ҿ���2mM���מ6Jyk�x��$� jL���^��-�环�4��ۢ�M>���S[,E����:w�X�yR��+a-����]x4Źj�Aǋ��ؒ���V5�:��Yrkh�3��h�����x[���t��	�<�p��mYP�z����lt�92���b�n9�,���-��\TiY�H/{���Tr�c�aƐa�e�"�`�9�mǐ�-�e$�B��g�j��;�3�LA��=�ME0uiF
@v)�r����u���!�O���f��̉�'�WpfE<wR8��u���]�z���Z�5�6��ħ 1��	v;bk���
�2�$Y�{�������LB��mP��ḙ��f3@|*��� gs�~K҃Z��V�z�x�yv.w���>-�RvD����Fc�F>�~y1f�u���x®&�*��4O:�2�#�C��tqV�z�U%����w��H��d��Xd��1�ˡrk�{vs�������:�F�ݹ� �����Cd٩�+�N	��+E���v��@0�Xw�Q@>�`L	5F1�2d��-�$��ٔS����x����c���b\ՎrVq#���$�%��y�)"J,�u��B���߱�N���jB?v�O�U߷��Yș_�v�2��H4�/��w?D|!�bC!=�=|y�642���P�tocX��sJ��
v���3Yǭz�q��E#T,�X����'9w`퍛��=�ؓ����o������|Q� 2w��)[L+�z���k8B�a:K���z� b⢡f�̼������܁ne"B�FI�,\/���sg ��	y����I���ly��ǘi��_��;e�l��6�J���DRCH�<�Tl�<�o����gU�1'��d�S�+uj�AW�'��n���
܏ð���Z���G,�D��]}j��������,�|Z��m�N�Zң�?{"5\w����j<����݄ǳ��:��K���5y�(A�vZب�S$��!G�%m���9��4���ƪ��B�J��H�[�?&}{T�3ǆR��>�=僌{���J��im.���)���K��#g+�<�ȫ~�L{�O�l^��������g��m��v��I��y�zPyA���� ����ݚ����^���)�p�ʳb�_W�{π�E�&+hͫ���1��]mJ��~�}����%���
�}��پ�ߘ[,8S/��e�6|cQF�N^����XA��.3o��'�Vx�E�ge���]P�ړN�P`���	(�0*�����. ��u%�Q̢U�{���\U�4V�^�Oo8g%��7@@ ��)��]�ZH�u�Ѹ��?Yn��=�Gi6w}R�����$Vg�o��8M8���$b�����Td�v�'g��4½�x�>����k��EW����
Y��@��������YiC����!x��墯�û�|����&.l`�\C$���NR���'ӝ�jo��	w!{��ұ�`� ���w9}�}����)D.��?eL����)�Wm���gV��j������w���^I�O��}�ب���A�9v��5���fUN���P���)m��|wz��|N�OϭG��HN�����m��1BC�b��_� h��#���˪{I[<�\�/c�}W��Dv5\�4��m���Gۯ�ɸz�D6���"D�v9��!ٗv�M���Q��K��e�o<S0�>�܈���|[1%\�=8�O�D,���)��v1-<F��G�����&"g����Tk3����h�Z�ZH@j?����2�Ǜ���6�I� ��|�XJX�l�H>�����,��P:�%�8H�MT������ ���.Կ����	"�7��W���)֔H�4�CG3���*��b:����Z�/���<D�Jt7��a�2�_�Ϳ5_B�y��"Y��,�J�6G�4�1Bm�U2����'咑�);�&�+�B`��n"�#�9D�j�W=���I����C~m�K:��R]�d��L�#��&��R���������-�0x�rqi��j������{6n7S]�5��Y�aF �ګ��`e���v�B���+Q!v*��Ȣ�I�siݢ5P�!��;��(8"�t��~*sy���tU�6�g��Q~���?����M_�.��MÝ	h7���_X]nI�u��n��T	XP8��ڀ��&��++��V���$�� ������[]�45���y��>-����BI�/�����
5����-3��sa1�xH�1N�űew+�a��L���iȝ۝���*�.����2���?g4�0
y��mWHrƆp���4�'-��S#3�9��}1�&K�M�_:#��G�@P�a�ׂ�j��]3���ֱ1kl%?�;!����$'��)T���unI���r՜�؀��»��Q�r�jO���'I���ʟ�c�uV�!��h�%�5Ks�FcR	(Vs~��F�?Vj�TxH���X��>�����$p�I�S9��L��@�J��nu�|��#��R�BOH�B��&V����n��Bΰ�	�JRre �u�yvA����������<Z�p��?��w�v,3B=R�C����o�R�����V!�� =�c��J�)c/L�nPN�`-W.&�	��5p]1;���ݡ�KK�����gπ��]L�.�@$��Z��nګ����i�Y��<�W�Yo=;+-Zf2=U�$�ojX��@9;ZQdC�+���KF�k}����\P!^Cv'�F%R�\���Rѩ{���'k��v,��l��֚�6d��9���e��*��������5C4�]b�^�shr<EaW�Wx�8x���LYA�4]��`r�4'.K9�y�|�)�H)js��ڢλ��p�xw�����	D<����"FUL���=�n``����i��r�7�T��/U�(�O���_i���f,�9��+�m\����b,���ԴuP���;ŬT?GYꦰ��6Cۢ.��Z�vg�f�שׁ4�|���]4�}��g���:��vk�����p�\V��j׊��Y\'��qj�pEa!�KJ��gV�Z�jd}m��.f�h�2O��H}�w���-��I��u����^i녈��o9�� �G�.H�f�m�V�
�_�f��_[�|>�;Gh[��I+��p���ǾA'�3�\��E�Y��Eb�d���
���1�����'a��6{�Y��������/�$v����P�ռ�@~�sv����1��gSE���$���0���·���1|����iP5���=��Ĭ�T�2׊l�����x5��A]=��<��e�p��4��r�$��=�fS�嬣&.3�܇冰�eY���{���v��|1`CA�G�uͫ6A�,�r^�Yk��[!`[6ȉ�A�T�#/��*w�ݢ�e�D�S/䗨u�~uL����-���D��8��aP�km<k�S0ep� k���F�O����8�����* �x�Zi�7	�h"q
XJ�V�U�$��p��K+�hi(�PDi��'.����ı������,����YM7L+/Xp�C����I��}��	L��+��kS8a.�qg�)�
Ђ3���RyH��0۲?.��k#+���j}�q��f+^����U�3��'
�������S#7%ޱ3�ƁP�E-����?C�vn� F!�G��Sp"��X��k�o�;V(��J�˾g�g�Ԯ�
����ߏ�}�6G,�v���F�wI�S�I������QpV/@�r�9���u��	'�kئ�r�Ë���&��(��+7�(�Z�Y	C.Y(a^��(}�~(���E���#���	Cc*��b 3���C�C��J�9/���Ky�΀N���(N=�p�����1`l%����:R�Ϻ4`9�z���V�M@�_hy�3Y��ƈ8����Y%���#�sE�,WQ�q4���*�{����k36��es]u�f{���.Ue��R&���L�Qnw��1.	"H�S���h�;�X��.��F+;-��qa�/M�6��R᷸��t����ų?��� ��G]AO�������ć#�Eܿ�y"wz!�{��X*��E�X�l�=������/˩�mVϿb�L!�&ū��\�g�j���X�~I�!<;�j��[�-�8J�p�ő���<)Z�Z)Si�ܡ���\����uf�}�c���T���ėS($c��w﬊�H�;��^_<
���`c
$ݽr2���_����+f���)M�_8]Qr�Ch���;��TC�@�#(���&*+XD���D�	�v[P��A9�G�@)�}~���P�p�j;�Ǧ)��h|WҖ�����c��8�F�����,�9+��}.&E@�s�R���;r�&H��S���/��S �1ؕ�[Ě��)+���v����8�BAVo���>�Qe��?���S~�˻�E���3B#銐^FAKo�K�5����_�>W����k��~G�}�h��	@���l:���_�	>!�R���}Lx��9?�����(�5S��$U9��u��@r ���,�ѳJ�?^JN��!cK�����y�c��m���*~��|�F~��6OEBi)/b��j�b���/yU�9�w�iR����T���ﰝ��\���M���L�l\�AX�ʑ�I�YM j�W㈋��J��lJ�Φ�T/��6� ����қ����&u�Q�䚯��+9�(��""r���w�*�#$`Qz©�n7qx�V�uԆ�s�ʜ#U���"��&L�ے0����HV�c��U�ݝtx�zk�
���|U�P;�ȁ���qw�2�Op��!7�Vs�U��<]A9�ϵ3TZd`���EwF��^�:��y9ͅz��4;���Wr��;9u��fD3�4Ub-GYZw�c�&�(HX��x���W�l�[�(J޻����zzbh�#�$�5|r
�WH� �|��4����gVO�/��C��W8�����Cl�P��%?=�I^�w�G$�z6Za>�����ۄ��u5!�N�w'�=;�z��z�r��IE�W����������SR�g_ ����&�tH�@5P�o�ȭd�Y�QxJ�%nE�H�N���VB���p峺��.ߖ�3ɢ����w���|ŧ��~���]7��ν���2�h-T��',_f�9w���ul� �].�ܖ�U��=�X�����86�-~ll#RFշ�nGo�,�f���xĪ����5^�A2�(��'{��nڅ�#h��A�$ɏ���~������:�S��dʲ�����G�n+aF7�wm;;�#�V��(�S�1d�����0� Du���ԭ�S�~���jE��mtr����dwx�0��o~5M��@�jC�ԁHy�Jc�_�4���cU�MǞH��װbJ�e��}��������W>�ڡ)�*I�B�*L��P�MYx�������M�Ty�#�:��_&�H����S�Б�;���������[�6��E��}���i��U/ʿ�%m:<��v���(�8�<ɐ2
J#e�蘀�K��,ib�K*N�ӆ������M�y@ݿSQ?�'̣��/+B�@;,�'��8
y��x!�|��Ͱ���+TK���8��F(�<\{�h�nŃ �����7���7>��`V��������hyg��y ��Ʒ��O����;���mX�8ݢ�ۍ�g���B)��D��퍶/�w�=x�R�%�!���F��TJ�aπ!\4�Av�#�H���3x	!�,�ZP\�=-O;�=L�/]��ٺ��s˥���vσ��dM��p�o�9�Z2r_Ә��U���:��]���j��ͧm(|yT�'B��
z�����a:��iG.*��ni(�Fh�w�K��〬f�X�J�k��";�[�L]�JK�O��-����W��[�v>F�X��@�m�|���;�)���*yN�g��#~H{kk�����r�H���zQ�������I�Xv��O���j!�{�Q���n��^�l�F�����T�ǁ2va�>*��f�k s�����5##�&ݕ�y�EF��b��p	��x-.wt�iR�`��ޜ���f_z�n�
�Q4⨳x����B�3}=��vW�6������-=������s/g����D�c��)�m��P�{(�gv )�;�_�2�6���O	 �|N�T�0�I�^�մ���3������qwrdWЦ�+�<>����Q�K����vE�ݔ�Q`�#�1vb����q�J�7��� H�@v/�T!� �N˗A=NX�'�NA��;��ik��vrM����ut�1�\� �^�A=j�{�0�ϣ�c��s	4C�h*�����b�(W=�X�D�_�@������)��4��Oߊ`�V��b��f��P�I���7_&�-��wv3&���N������On8���!y�VQl�5��/~��
ҥg5����i�6�����؅���R,�<Q�>�{��9��ka�{)t�"{�S;YP��&=E����`s�<������U���.!����^~p�3Rg���D̀z�L^�ѫ
� bځrH*�g��`��T��j�[�Y��K�|J.�*[���r>h_?��ŏ,*��&R��f���POqc���M�H��>�f\�����:x����b�J,��4w%�V�ڲv�(����p{$���#��x�	�� ��Zj���9��!N#V?������zJw��7\��A�u R���Y_ʀ�tnN���V6ʨ����!�Q$��\|�^o ;�3]��'�xU�"���I�x���а&U_V����5�Xd��t�E�G��-�dT�{Z%�W��0�ɯs��)þ���]	nF����H0��VU�=ڬ�,ã��֫\]��n���g\?	@0�)��W�i�\9e�(�� ��A��f�|��F�	�`�!�<I7z�^pR�J������՞̕�&�揢Q��,/�+$hs�`T�`�P��LsI�.F���
j�V}/l(M����N��B��p��O���%�ʪ4<U���u�5���LH�}�mP"��M|?]�7q���N����g���E8Ş�7�+�@~s�Æ���!�΁��r��i6�lv��B�u�\�g��]P}7"Iܧ��#�������d�z��hKzhM��V��!�t�@U]1�A�mՕAʄ4�=xǋ�Q���%;�E�@fҠ�7�b�
��r�վ����\M�0�-re}�?e7��}@�!q
�`��e/?��?���=(�nͮ-28'�d�iV���O�^R��1�MZ��a膤�9�8�������T%O0���Q �����V�'ǹ� '�[�q+�2�8�&�����2uA�blq�ͳOs`ὕN�L��o�ϖ����B	��.�3��z2�KX	��|��.��#s�wL��s�3�����PiLl/Ŋ /��_����
�+��~l�a7 �T�h�K}�6m]�^K�u�b�V"�_���
``O�4�/7S<��F�ͫ��	�f_l�ژ��q�1����{��kI�r�@+&z�|���g7� U�1��`貃��I�!c-�������qu�=� ,6�J<o�����N5�ȇ��&M���&�R�9f�=q����������G ��L���֠B/�5\::�>��o��`E�{�J�`���[�~REʠ�	87'�Z,>��4�5�	hp^�R���9��W�Nx��3K�z�fН_��S����9��X�60��&TU�A�1J��
�G`�L3�q��s���l|�ҏ���ŔΕVF�DDj?p%+/9�U�����5��jk���ɣw�u�+�����\�JwZ���{���F[���l�洫3�K�Nj��F'��ǀ�5S�cQ��ptߥ ��&È��P��  �a��rG��O�Er�}������F\R֎w�p��r\��L:�eT��(���D�%ݾ3�0�j}O�|����N#+|�c+ѹGtفu�a�
IM���C�>�r�',e'
?K(%�4J/�B0k�������/����b�媚=0t�Dan�46pWZD����+nj��۹�:�;��������ݏ\�5��_>�)W��'P|���[P��I�0>�LƗ.����gp��t�B!��}JְV���(�|��;�� �PrQ�U(�呺x}��	w�Kg+���J�o�O'��3+��`��G4��}��0��Տ2�g�X#t��� ��+@K�~|�O&}k�|�'y~o�-�B�N=��XK��v��h�:1�O�NLƖ5���7+���L�h�[@S��S����*b3�E�P��K�l�b��bd���+�iuZ���1~7]�ģ&cf��9.�w��j�O�oю�P��%uͿd��Z	�`e�Ծ]��EP�۬�2�΢{�l�l�A֪`?�I��9�JZ��K�_�������$��1�o���]`���sF���ٌiݽ�K(���aQ2K'�<l���"p�s^��+$ �5BӶ�����Z\���^x���� <Q-�%�;-��yԁwV����H��+����>|YQ�9o .A�6� V���G��"?#���N�AUt��[!9���"�0�W^ٺ�DI��5c�G���y<���=��w����Z}���	��H�����&�U�C�A�