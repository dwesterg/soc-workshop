��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=����A�ѻ� ��v`���Ֆr��S�=n����w	�B���p�G<�6v�^�u9�ۘ wm���Je͆}D��(�Q��f�����%'u&�
u�^���4�r�
�{%� �B�3#]�U+JW]k�^��&+&�î�q7;���c���X#���$8^��$�����l�Ftr��K=i����`�4^������
��e�4J������p���-���b�v���!���cI�n��)l���,%���a�:�*�P�R��g��@�������W�"߼�R8EU)Nz�+�D�aވc߂g��H 	��N�l�4D�����|o�	�2}r��Z�z��\z�[���6X��!�;z���,�����ļ'�@�P;�n���;�T��2׏��$D�8�����o���c}�ɿ��'���K�ukܽ=6!� ��M�����?��}N�K���|~W^�ů���͔��/6&��A���<j6�!^9������s#�5���k+5��]��'���|�)�E��u�_bx���񆞙�7�3����9�˻(�t31j����q�'oE�`���'����B{_�}�3v�@|����)���ҷ�u?�h�n\Q9�0w������E��{��l��]t䩻޺��e+�y��}Ηr[�[\����F���t��}��x�.b��=J�/\޴Q7-R�_�t�Ɯ�1�:y'�p�t�F�LU��췧��뎠��*��C�>`�~R�x�Nxr���\2���t6�"�bJ�����N�]�r�*a7����$���O�;������i吤�*D�Z_�w�#�8o4R�?9�Ȝ��l���Aߟ�5�?�<�/�Ҷ[u��tz	x��E��r�U�ߞ.YՇw!� ���Xĝ	�Y�d�����B��_�p樄��"�XD���t��o��od����۝�j�*���-�Cz0�4�-��u��<��QH���n	��&�E	|Up\1��ͭJ���=P �d�q�l����s��3�\�����y>�,��U�����A�=~�՘F(D�&�bc<���kԏ>B}A�� ��;�ej�7�8$�$0�Ś<�����o�Si����F/�s��d107V�F��;h�Go��xN#ѠpTG[�t�_<�B�Q\���!��IV��:���G8�)��2]-#����}��e�}}�^�r��|{�c53��u
J�
؊4%Ky&��U�moz�ä � m��%%-��C�%���"��;��X0�k