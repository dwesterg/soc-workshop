��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^�]�� ���6����pL��]�G�)�mfB6�q���$���]C���p����+c�n�� ���w�5�{JR�[���7'mɪ}�)P}ٴ�>X� �e�l�;�]�;�c-�G�>�."u���߯#��=��$m×�����5��[М�vM��i�\��	����DG �e���sup�6׌Ε���G&o��՚���lw�A	��n^�}-��,F��J����3�^s�p�}��
' `U�7>�����|�Z��"[��"�5<��^e�bzg�����I)ͫ��K!N��I� ���GA���8Y�+@'E�j�	`a���;���θ) �v!�΄])(���+C��J2h�_t�.�����,�S��t�֜�BF�װ��-�{CQ6�;��c����:�0xȫ}J�M_�@�u���*�I ]ns9��3�<�ǁ���u}��y��̓l�F��*�r?d�\������tǎK�ޔq�h%`�<�<�e���s�ũ	�}����?9�u�J��qW v�j�Z���<#41%�Ӣ��wj1"'�.�%9�G����l��ҏ m޶�����5��Y��ܒ��/	�F�[K�}���<�⤱#���* &3�-�ٛ�I��7��A��%-\7u�P,���C��:T�n�.h���1���j`v���V}U�__i�I��kKwQ$�C�Q�����2�h�Bd�����D$R+��O�3�����g�ʺ�2dȎh��N#�Y�{���#N�T�f��+R����R�{��6�������ךџ!���8z{퉛�*E�뒭|b�c�m2S}�q�V��ŁA����̬�/�l�2� ��ֻUe`�,�eD�h�Wv����7��%%32��&�|��?ӈ"8*�^g��$Xa	����u4H�;�tܑ�:��l7_��	{5�j�YOi�n�?U�����L�B�r�	�úP�O��\S�>��,�_���ˮ]hfj��o��t�#�)��bnd43�6���V7�~�: ���r�jϨśW�K�Xy�m����8ˢ�I�aC�V�9�bh��ܯ����{�0_+���:v���6WBʫ*��~ͷͳ��ȊT���8��u0v&���샗E�:�"�~�����@���[��R��iz�m@\6�"�H�|rmZ$W~D��b��kIH�L�㤤���l������>�)NV0������E�w>�"w\�z��bM)Y���[�*�AO١�d�)��¹�+�ٍ�)������(�}��7�-�q�Ĩ���I=\\=�|]d+|������E�A�܊��B2�g����� -Y�)CF#ʣ�`r���X�$�a�;.��ʀ=��� =�$dkݶq��2'𥀆L´�����q�͝���f-_�0��=���x�޾C�k\���w�n5в����}��ef�tv�,E�R�40�gB}	����^�?0����)��GAж���}ٱy J	%gq%�^��C��덯\v� �������� Y�h2K�*���Mɀ���a���3��3'���B*��&���P<G^�\����x����a������lF���Z�Ża*u��K�H1���4�6���I��o��9�j�K�R�'w���B5�Z�KI��W����EZ=yI�zh�24I1�H��d�oF����>8,W�o��a՘�[\�6u[�f��d^�׏o���ש�M��F,��~F`z{��W��"G~@��gH��"Q!�I����kf��q�#	�1I�"��q�Y�g��Y��LMk�ހEj(t��-d��
F�?�[W�o�y�b9��T�`ߊ���v���[�0=�$[Ե�ʍ�	� ��W�������uH|������z��h�.��ͣl��}Pf�piԧ�`��T}1�!pޛ`�4�sV�M]婸nJ�E��JbD��C���J�&4���5��3��FP�:��W�n�k~�H���5���:�H��6�H�>l�+�Z�1����l�j��ʨK�}*�e��d��!�d�ˎg�H������o ��L����o`�ꖍ��"t܏I��ZT�9gOs�]�����#�����Ơ�#'R��ma������h����orXg
����<8���\��Z^ң�{�6��48��v�'���qg�1RLw���oɢ�$hM�{;�~,XgWu��7"��	=��#1�?�P�*a�<Ҫ%{�k�h��H�� ǡ%�s��A0\���>��;��aƫ�<D� �Z$��1ZA�5���RK��c��Ct�	!�xqs4Jfy��/˅q%�8�z<MII���ϰwi��`}A�¿u�,/H��κ���T%���N�2�0�҃�{��4>�:��������von�����FN}�(v�|εf�v`�j��Sfx��<O�w�6��·���s��5U�#m���õu�V�a�[�]��0&�c�9
�;i-�#���X�v��^>�4��G=���"�8����} �hNX�G_�5X<V�t�6�v���X����3l�L,�ۦ���x"�fD�3�';�[���H���S���[��� �v�9�;����/�����,�L�����i�@mk�����<Q�h'��9c�; c<�g;����H�6�&gK�&P����<���K��Wt�r`a���F�A�g�����,l�'R��qda.��8e�����T��>A�C��6�[j��(_B5Ca�u?5��,�qť��9��Ӊ�
lO�u���J4󱢲�L���Y�iw����z|�vy{�����צ���I�;' �����Ǵ����0]x��l���������S ����s�̋���W���'����k�C�n��0�H.SV�E���r
>%9��pg���D�cF�m�(<g���ɩ5��ο�/�T�Z����>J�n�O@K\�!����%�L��1,H�`�2Y�%Wkk.j��S vڈ�K3�N��e��/k�L:��\'X8u����4^�0����2b��#��d'�D�����Tu��zI��%$:�=ZWLf�h�ԩv�������s�3�~|DnAu�~l�N��'ȼ��p���x.Cs��Pܛ$��BG)�*`$>̕��~%A���)��T�/�[�!t���b��`�C�VnCEܜϗ������0�
I���]����W��=EFDL��^�/�[􃓧K�%�E�Z�yH|�����j@�*xD���U.�{���nۦ�k0�]b�ݟ��rkvs{H
W���|8��UM֔��aq+5B�ۭч	NQڞ<�e���G�e%k�i��;�.��vĲ�(�\	'����������=O�M>_�ZDP�ˉ>�3�Ao8x�.9���/n����z����i���U�b���S�r��O��&��Ů�WQ��I$�?V�om�J�7�Ն���%a�*`�
Y^�rO5.���Z_]��D�I�*�u,��x+.�IaP��D�����d~i�0$G�yb��l����=����g�5H����b�' ��a�I�=w����~����唡�����ҫ���)�G|�p��d�B���U��b,�K�SiU�	��z���@��H��(���y�O��-��p�<�Z�-�U�%�g>�W��HB���qQ��:l�o9I!EL�6�ڞavtm��UwS��Z�<E�	��6��&�soU]ʔS�K	�����Tj[Ӗ�L�&Y��5�'UU��k���.u�$A���I��w�x)<X~Ҭ<2�on�)&����^z�,��e���N^�3���p�55	����X�v��↍�L�s4W�t��=ĹN|��4	�b��|37]IE����Du���1lF�G��wtuk+L�n0E�mK'׎/B�˪�Γ,#�͜�w;)*�.B�[r1�*K���j��<�]n�}��LP�J���>��6qQRu#�w�@KX��o�'R�����碣���P�y�����|8��-u[Υq��7׺:hܝ���)5�P�Y����u�v�6�RƩ�U�4�@�tț3�V�E�EZ�z��K�o��32�&U��������W6ӪI�_�FV�(� ���b�P���{P$��������S*~��S'9?t�I�U�`�
�a�z��D<6�[���5�ӥ;��������Y���L�eE��Զpd0����+��UM���z���2��=�]S���/_;�v2���Y�:?fΫ�c�B�M\j�hF�F�>$&�GP�R��Ճ�t�կ�pJUZUl#�S�����!�
���������76�٨3�<V�F�d
s����Ype�WQqI����iI� ��ɑF4	h��ưRIT�=)0U2W2<Ir���oNċ,��=�ei2Ӥ!����/ب��ҙ��D�W�����ҽ]����ZF�W��_1x��.�w����?��B8!d
��R.��dr�S�"��Z�˱�ՠ��y�9�SG���w'��������H 嶫g/�Rm�	%��x�+Y�g검Dr�E��BD���@θ@s��|1b�%*
jOu��?��,B���1kPf�(���ȹ]��ڴ����zGHR���R�܏�QY	�.T��kW�+�³~£V�v��	@�p�Jx�e����I!��m�tA�GI�U"+����FG��g9�� ���G��op(.���6d��S;�t�Ư�������̾�p�#�v*�ޠ�-�c��]�]� l&�V��AUGE��Ĭ������#��4=9t�����Pq� Q�R�%�!o� 6��]FԘL��҅_O�YTt>E�B'u�)�D>�����Q=�PR;�� �Cr��Ь��]�D�B��7E���E�	�z��og�Q��0����D���9��̭�_/�b彉>��.˅��V/�Z܀,N'����Se�\�9DE,��"��NvY/7e�MY��n��4vX?@�t0�������E�b6��٢:r�+��3�ۑ���P�@��k��",��?�:V�¦��� �FC��q2�<@F?���yq�A�<R0|k�~P%(o��Tb���
#76�Mc !b鮊k��D�w�K��t�����
a�> ]��L͹T�XE*�$�G�ɫs��>��p^ ,�[�P*X�����-�ւa̻=��z��n"��oE.Fsj�mK�l$ȉ�Ռ�yQ=���0����;���9.AӁ�]��~,�t�=w���ٴ�Ɔ��~�Qs�=Ҏ5�#;OX��W~A����ڄ\Y?���M��
1ߊ��%Y�����C�w	��k���hb�d���V��qhl�.ϴ����:q���T�,L_v�l�+n�ޏ�u9՟*W�ĩ�d��SW?-�
���Aƴ3�Bh@f��mO:7J/���M�--.ݲ�N&Th�0�����K�7�lMj�N�6�t��gB��-�ە�?���%�TV铆�
F���J6��m�#NpfEq��ir6�i���{l��oz�����J�A�L����g���R�p	�)��3����
�V�1=DO��nǻi�
�3\웦��q!��h�ˍ����E�/�|�8��E"��np��m�W#��qi���>���%�vO����[w�̎DB�VN9^�Բ���2�?��"*�Je�_�mL1��B��{�t���6���!�{@'J�6,�!X+��ɇݤ#~�ʽ��%�ar�$�V�rX�������VZ���?�J��n�!���]1�aX�����͹*=�~�`�����z�܆!��"� a��ժƉg�(�z��x��m_Z~ܐOOd��������cdm�,��,r���:�	Y�LT!��?��|��tC	I����[�w%B�rnוy�|��[tm�$@E�Ŋ��ڧ���P�"i
�WV�%�����>'ީ���nk���	wL�Ɇ�S���ovg�Q����Iu���w�Zņ�C�*X0�OJe��Eg�}2�(���k��p��}��I�Q('eH��'�e��Wd-�n?Gp�Z�| �>%)�Z�"�a�/��D�K��>��-x���z]K��]M�X���Q(~���5t'@�
���N�f�?�5��͗:T"�h���c���ݐ'5�f/a�=�X
���l�6xW*�HHD��^Ҟ�_����yn��1$̉ӤL��X=���������A\�QJ`��K6M�U�Q�7�5D@R��}��ْ��Kkz��V`8&��n�
�pg��C�R�ûP�E�n�o�4��'�	�Fo��C�'\,�̕t=��Ǟ<?��!�KA�������C���� ��I 3��Y�Y��}J��K��Q��E�S��8���u�,Sk�G��儍���i�\]|ե���~DpB�)Ʈ����6��1L.'뎨�oeg˫��n2�&������e��$��6�5�fGdi�Vb��/��'�E�e#�ʛ	Y�tB�r�1�l�@yDR�d��׍��nӝJp����	}�ZlL��о_ȳ#ݾRt�8�=|5~��9_�W� �Qȭ0M��ڱ�6 �8�)՘�ǳ������w�]�;:h��F���W�8��?Z��æ�r/��T�*) ��iVݸH��&� _\�c����7#L4�����G>�q��v�9�'��Ny��>0k[�7.�zOk*��0�u�����JE'�;/w��Uypw�_m�B���΍��f�6�yi��IRfr-�Ґ5!D�����9�<�̩H�-/̛ڜ�#N���b��KU�Ń���ý=��/�iE���{#����7��/V�V<Tg�\Q 0s+œ���\�k��;y���[��C������6Ǽ�����i�Y�lN�Q��HK^_߯`|9"_��D�jU��Nj������-�7'�t��=B��NS�l��.���L�U���*�>G�uy�������s����F��s���A����?�%u��Kr�Sx�����q(�1��@�'@�	N�6|8�,;k��7�]N}_{���u�L��Zt������;��y�``�)�k��"�k GO!>�,�sœ/z2����3������jn���~v�#�O���;�ԕ�_�xD��m8�8L��n�ٺ@�����]w3I1��㿴��˜+��WU�E����3��l����9ov8��*���[2. j��}-s�s3L�-�۳��ea'ñG���Mx�vz�;V
�:c��z���6�'[����Ŀr�w�st�F�+�f'��H�-��+�,-97w��.V^I3<[� b4�։�+��M>Ͻ����7+ݖ��h���7��T�m�N��)Pu�h}Z�$+t�&��E�w-Ĥn 3t���o�)�銎�=�+��4��FB�|���U��HQ1����df���-�%��n8KkIq���q=���C$ͥ��O
�¡�0�{� ���3cE�V�C�w�̸
�aLF9�\����xٍF�x𙾢x�B����(�֡�J7�ڛ5��ָ't�vK�M��
6� �I�lDi����a^p�"�����a>#��)9���<��wb��L Q���&d<��(f�V) t%}ع	Z�1,`8e����|�䄵:r.@��_$^�c��Y�q��GQ~��@kE��\1�ԥ<�+o�A����O�=��������E
��N~u�7����0�D�-IK�!���H�2��;p6��9���K����h R�PQ Q�+b�hLb����'��2e�ev"��
�m2���l�-m�D�"\TU+���NTjނ�O��.�PJ�b�����+ؤ���t� Ac�Kn�\w,�1��.> ���n=�eD���rAh@����\K�?�C8����.V�x�&��rߎ|8p��ǚ�� ��F�w�Q�eB�8��{��#hɢ*OL�i��\���7�\�l��	�-
�f�kdE�b�7���|~��ś&Wv���~�$W��C+��b�Ω��=��N��`=������{�e�!����Lp~��j=ǂ>m� ӽ�Lg]��P�SA��5�rT�꼎Iͭ��¾���~!��pJAR*�臼tW{������K�������weL�����=�̊h����`޹�w䕔��\��WvAq���Y}|���ǵwes��0�ЮxS��}+Cf^b,�f�guX[��f
H��ɬ�%�C�j&����� �����3ʈ�K+5�Q�]�n�{�O
t��#ciXx���ۼ��0{�^�hdg��4"��������\��TY�� �$��pFѭh62�A�/狀#Ub��7
G���OҾ�ܗ�aU��R���zCu󀝡�H�8���a�4Y�u@ �����u'Y;��}��\+�<�r���(HY;��V�U9�Xt�Ϧ���Q��B#�K�C����xitʍ��*_�#�t�le��w[�j��!�|
f�SQ)YH��<�tܨ�-C�A�l���X����I�g�oo�D#7> ��4���������>��փ��Ŋ�����b`��=�>�]�f7�!ыG���SƎ��	���6��Oj[��p����Ҩ_��c9��$��?����em����}�z�P�������|�yG���b�����SR�xegl�8[ظ�T��,�p�=6�g���A�҂��M��E��Z���J�Ё�_��P��%�ٵ߃iq���X"9szİ�)��n-�3���3^t��Bz� }�&�ֿ4ƽcí�����#���5�*1�ԕ��R<v�ơ2+��o�c�|ßx@��IM'�2�Wj�b{"r��yM��C���o��Q�	Ի�`�c�����k
�O���z&�s��f�_qRZ���-ď�7�$�# g�~]�`�t�b��"X���P�V|�qw������������$RLif|���Tl�vw��%f	],�S0��b�����D�_���!�@��ã��DV�-����ZQ�K#H�?��q8���'��U�_\������r�qU���L��X��޳3Zܬ`֔ٽ&D�T	t�����*u���I[&@��vn)��|�tR>.��o�I�:שxU"W&v�T�n
:��qx Vb+��(t�me���g��i���5f鴱�*FM�q������1@�?���#7׋n��S/��.�NZ�`��.@t�ↃQ���m��v>�.��yf��\"=a��Jy��bYL�aXk���N� �!Y�EF��~0[���uN�y�
�G�#���e:4hA�b8���vCK��}���B�us���$CO/��8S�gZ��|3���c"I���:H�+ g~xF
�l��A���C^1Q���2F&ͬ�j\��cӈ������R�ft��y5��Ύ����0�$��Έ�н^��ӯF��ڮ��kr �?��M�aPߋLã��J=Ԉ��
��$�%ϑH��#�/�"QN��]�g'��3����$�/ گDv�nu7C�;��kE���Z�����^�0f�0�F�K�/����T��<��{�mJ���v�7zt�qf1Vp��H�\��+�����l��L��8���u$x����?��������&�y�[�6[�66p����vͱ���n�ӫ1��g�����-�U�p�&�iF8���д�u���j���ڃ��2���ӈ���b��M���YV� �S�
���N�g���S�൮�ὃ�os� ׂ�Rg^�7�|x��I�%�<7�K\ybmY�T*1ͨ3L��N< .O
���ۈ)QF�h,���3�z r�i����0V>�PK~�Gs��f��ꑈ����4��k�t,<��ݰ6�����>]�H�t@^}�2�R9���Y��=���P�A�q=��8]4�k7��p%n3��?1�n��3Y�s(�Mw�Y~�����=p��r��npc�ͧE��9K:��P5��%m��vI"4V��Q-[��t��UW���G@e����+Q��@%"�E�����f���G�EN�*�3�	�S;�&8��-�Ҟ�ҭ�ݧ��:�D!������q9��?3
�du���;�[ D�e����N�p�~��@�1Z��V�B����;�F)4��nCL]����?�K��eڑ��Q���O���),Nu!�ӵ/"�&������L+l�P�������[]����T�~�������`��G�{���MY=iPN��)�ɨ�~��-L��4vwj��f���7���	�X޻��^ �:b��-�z~2`�0�CON$6��L��8ҟv�4�.�}������>p���7�A�UN�Ҫ�~��K�Z��n�з@��X�bz�@�x����t�z�iMlP�R�4Vĸ��S$���؊��+Y�^
�J��+�4B��ɲ�1gU�,�	P���{��(Kw�)J�N��?n��踕���:|F�s��K�v	_��U�r��6OV`��K�WAK<wԏ���^7o��[���tØ�x�*��"���w��D�Ǣ�z .kc�����K�Yg�W⯝���ޠ#,��>sv0Y�R��՜����'x��q���ǟm3|���W�Щ��Hj�@�! ��#��H�]�Fg	c�m��hs(�/`��7c�6Oڦ���Gm�
���T�p�@N��Bh��ýG�GF;�"���7�i��y�kK��ĭ��s�c��X���>z�c�L��K%�E��if�)cg�t��RfC�C��n�?GP�U��	`�)���p��܎����8�ֶ�<��y&�[�<Ga$�Kc`��uL Ma[�MaS�VD�0���0L7����2"'b����)mď.�0f�͡���䓅���⭝Kv��,��ͪ;F�+���g��Ӹ�_I8!a<�x�
%������eS�+?%������E��w���<rL����6 4T��v�-{�~�3���R����W}X|��k���^A�_%���0hג���X����_�iܓ� ��E3#JY���$ʳw<�6/W�,�[}Y���H4	���H`f�{mE��֔4�$��s,~!#1���G�CR庸y�m\2���E�ϰ�u@����V{�[��y���TЪ�5-�U�C��
|��ʦ�}�_"V�/rYֈ�s'"�"��ɵ��%����O������$�] �o���^�� �D_c)J ���q0JÀjH�7>k�p�l��!���{�9�,�����"�|�H��/h��L�n6�p%�5&�;,f|���/a�g_9�E�:o�3_T�g�0h�V�t���C�
�?z�v��#��,�0�ꦽ�&F���+�?}�p�ʍd��1!�u�/��z��>�y[J��~f:�cj�v��qwk�bp��m���u�����JdX*sv�%���)?t�U���U���]�.���T\�'�]e��}�IB�Ea�,�"n�@�e`YO$HnW��M�hYW����������m��eX�t`����S��t��C��0�D.Cƽ|�	kF�&΢u�U�@kztnX�j^u3�&���&���չu����xڗ�
�������j�PI4�~�IX��I`�����	_��#��մ��yN��[(��<I�v��C�M<BW�ĝ-��PGu��i[�O|���g��K�����u4��m�W�`����� E���.B;��J��@
NJ<�v��bAp��]8��UP-���%��μM�����e��d��@���%�X�+\��J="���*��a:����̖�rZ0��I��U}��7��\ �CB1��HM�|@!��Σ�� ��Ap��*(}	̚`r�'N(��^5|��|ɲuГ�J��A,�#�J�Gcy��*�@{&��$�I����cg3ǹ���Y�r(F7�¾��<�O�P{"̉��lܨ�l/�TȂ~�W]�t^;�0��S���Su��Yk2),
�c��2۞2��u 7��&��r�'hGE�����u���ET�1��A�h�%���/���}��-^;��}������V�愚bŞ�3(�`�J�َZ�C��g����wq�+:���i��q��J�9}��3{���M( ��e��U1��~�6�k53/n�A1m3�Qܣ�4��r��4wo�l�,�E�؞����`�X{{���En�	�2���p(�ΰʣi$��*����*K&-.�Z��r]�Y���BE^5
�ߜ�V�����qj����*�P*��OE�qҕ{��쿝�[ ��+���r"Qze��n/�E�'�L�e3 1��ȸxυjG���7�������y�*���;��i;��0
�q����/���<?ckO�]���ߟ�_[�^ �OCԛ�PF���srٳ<-�����Z¥%�ܹ��Qw�\��bƁ�a㙗,#7E/�H�vl�B��-�M�Bw��Z}�䚾y�6U[:�͘��6w>�}����]H�d��
Uڽ�	~U4afWTw~���5?�E�hU�6;�ϖ�u�;#~_x�7���L��E|�UaY?����),�����²H��G�H�̑2���p<Gx�د�W�On��Kf/��	���=HG�(`��i��bܒ�Κ|V\��;�B�(��=�cݻn�d����=�\�?N!F,3Kt�������0��:-�������6戴�2�?�+֙4��NM׮ �Qd��BT�ڿb�=�a���f9ڙ@�)+4i� yx{��F����"3� ^p1Q�SW
��)v��TgT�LT�-������&�*��f^ehG����k�J.������Q��w��a��]�*Y8d�G>[�N[儖��E����R�XB��E��Bw���9��r�Q�%ݺ���n>��C
`OQ�4�x��/�E�����!�ˌ��J�,���< �*mY�
c+%E;c�~״��Gn�0��K��^Ug����p��e O�p7���P��8���y%q*���_���"�`��8�	�c�P!ԙM�>O�">�R����!,91�v��6XD�<���=B(ᨙ[���и~��]I*�Ct*K{i��YA���&�Y���6�!����߰,��bI�Y��rfg66�m��?�.�W�i��,6�����:B��|3�ۓ�Դn�J.L�OѬbX���EXq��\���=T��Q���hJ�㵘=�R����RA�r��n����Mr�ㄑ�߲��-��<������qJY��%|3=Y�v���K���1�m�
�)��w����.�i�_�s��	~����	�0ܘ
ҝ�(N,��"Z��V��&�+?����>��ʃ�R� Lx���=���GD.;�&\QLb�J�+�瘫�-"&��}\\�/�~��
���}�/�ڷ �hR���6���{lS����c�ɾ8|<UԞ��IT��;Fژ��fɝD����л�q9$�-�-L8�/^����Mp���;kx�x~�H�`�~l��	�����,���.�cB)�DBF_ߡ?����b��M�� �gp����^�r ~-%�"���F��R��Q���q9KJ]�V�/|)�U����?�ׄ���O$ks��|k�M�{�p��}F�*�=�"��p̋4I��K���X�D�ovIY������+r �8NOEy�>�X�*�|)�骜�aO��
��âڠ#I���х~����� d���e��/s�e�#`������C)g�e�Z0́�0gx�8�{!��w��Cw���rPvT�J���l��Z�k��D@�?~e�6z�W� �1�WE�$�NE�y�MDU/�Ȝ�]��!��RE�D�d�}��^�Q��U��1���D�c	%�E�9�Ȕ�k�:�$�УO���m��u���Ґ�Q����	`��rx�vW��y�HW&惬��7�cT����Q�G�����i��
p���?��;@�����N\	S�rV=`� �"{62,��>	Z��Oꖥs��fp	F�%ܩ	��k�}��a$�h�+�z�&N��l�K$�Z��!�횅C�9ڧ8;g��/����x~���dMrd�X�&C�˺��Jjyk��V�X�,�R!��B&g�G˔�h��Q�%��@�x�<0[��Zٛ�H�H���˩�6�Q���"j̯7�_��%:�uN���u`�@~Q�~���Վ\U�J��xfSK��R%}�D��+�鄤"Z��ߎ��L�4��I�7��F�h��Q��A!�F�s���Lj�f\��M�!���O�`M55�c���99J׬�B����8�ǽ}^:cD��ͱ��SfZ�c܄�#OѾk�>�+|�N.�I�m32���Ɯ%tR�;����Q��txԔ�3��#&ˢC>����\ؤC<����@�:��ѭ �.��+�'`���!\�GX��n݉z���خD<����g���h����[x4hZ�z5
�˕�(h�/�U*�Z�.��/��s��6{?���j�9I'�c�b`��L��ŕ���N�������.���g ��wG33�]P[�7�bP婽K��Շr8E��?�C�m�z:5UM8���Wo;����u�?a~�6(�8p8�Y�bLN\Hc^!or�-�C���|X3)Cf���!*[:q�R�h��	
,������u{���ο��I͛�*X���a�NܨM�_U.�6ı�jvU<Ј�2�����h5)Xpp&s���viL_k��N�'����D����{R��Z��Վ�]!e�Xb�n��"� -{�G55�ɟ��?_L̜8-�P�ș)�()��M��wW'%��@�fj�2MNבc�a�f�75&���g	�*Ĵ@P�K�w���0���,t&\�*��b#�pW�=�J��Nה0|��%P|*t�g�6����T�&�*�/���?��Q���*z��̙ҦA�#2�fR�}���ATP���j���| 8a����%� ��~椫M����5	k���J���a�Yr��yH���ǣ������Ń{Zi�)��Io����b�|G�Ӫ_���$�Q�]8��Ipӄ�5����,��zPH>Z���&��dv��ήlUUH�u�uV�����lR���tdL掱r�0�������;lg��KC}��WEM�x���\I�6Oؿ>%�,��ӌ�[8��G�V��'A)B �?U���lL%��[��,tF���ҝ{ B0v�'�Qt���xK`L���c������?�z��~(� h�����mC�|�i����ȚM��)���,���*Nb��"�Q��y�)}��g��._a��#U�h�ԖE����j]�j���z��S+qڢ
��T�k�$���bx�I3YY��h>�o(��G�r<�rW�:~��T�-G��!9��F�?���)� �3�5��m��h��x�G&���mh���F���յ �zo4�	S8����:b(Ro:�#0�ѩ��(����E�ǁ�7D	�4�S��f?�=�Z%+!J�cH����g�/�}��i�d�o4���n|ET���ߎD�V6y���Z7�^f��Mo.���0ON��G|�茔xJ[�K�ٙ:��CMtp5�h-���3�G�1-�s�_��͗�W�wM]Y�P�)��Ē�B�'b1�Xv?�_��>m���]pl&ܻ{Q��l�]��>��/Y�M�BE�8��*8N�_o�u�ݙA�٦�@����*/Q`�m�{�T_v�C������I�Q��C�)�W��$�=<ʩf��9>��bַKT3r��1!#9�M^�^�7���1��&f#=8��B7��fD"qw#:��	�Y���`m$�~~E�Ee��?���R	!�����$�HQo��o���I��uxD^�ɍ���Ŝ_A>��A���|ӕtt@|��ޮ~��м�`_������L�&J����h��|"�3���:Vm�Ewwa#��3��Mj�Kk��o�]=��Q]�F0��s]��Ms����ᬬ�����S(�~�9oY�@��
���hN���F�	�:�t�a��-���{����;�i�K��X�b�k5c9�h�H�K��ҏv�b0dow�v�L�ۯI�,� �|��;�2>�6ۖ��&�҄-�9Y�ך�i��~�N2�O��w:;�o�e�0|�u��y�������5<5���0�ES������h9  `�Gԛ"h!,�뚘�r	���$�}y��[�u�N*��:�7��ܹԁ��/�ƛ�[+�j��1�:ˁϫ��9K��Vյǈ��U�F�˱�n��ژZnJ�1<��Y�ؓ��
>Ҽ�ZD"YcA]� ?����;2s�)~Ă�`��m��B�}�$��"�����а��B����(%}��?4�|8���W�
M��w_폍"�V+7g��K{=
�ꦺc��O
Hz��V��0(FU������S���To:�������2�2)�x�/�t�|��!����e�
�z�s�d�Ҥ�fkU��À�bX�V���5�p��ﻋWwo���]�+A#��à3���1Ə�j�;}b/�`���9�[��j�Dzr���ʻ��A��H�H/7��hS�ۖ�r���P�9f H݁p�A-α�`rt�N��g>��\d+�H�(�~��^uJ2��t&�åC6�͞;�FWn�k`�>�QM�������: ��m݈d����x�@ K������4�z�+��Q<�:_c:; Q���56�K�ㅞ#k�Xt�J�-�L��x*�(�\An�pC*��x���rɮJ��U�?�p�<��������i��F��b����ͅH7i�.�1"IaIt\�)��-���nE%�/G�+ͽ2b�3 d��A���s�$�C�ԊLWt�2g�r�<�r+p�0���@*�M[-�'6w�X(!5���#e0