��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf���B{��_�=2j��`�C�������7��aj�QTV=T`��k4&-���p������]���fj_,ُ�� 3���"a�b.V-�I|S�}:�I*=
g����vD��N��*^]�lDY��R�p�;�U�9?�0�:�ǝ����\[���;��Z����(��:�E^�&By��H�Η)�4k(T,f���F,K���J�V���#`ftc���e(�'�w�@`:���b�0^~9����e6����Q���x�u��ׇ]1Sp�d���gZÂ�����M�Xkf{�
{Pң�(64E ��s|g���lw��c�苪a)ߊ�@{$����R�_·���?
	��*[�iQ�����S�����{0̥f�7S��#�~��7T��L�ux*&0/ϥt"s�.�܊�PS�&X�)��Ե+��Z�����y6����*��DG��,�:_?X���C������և�%��X���4f���@��J�i
Ľ@!�0 oS�E��?Z9���v���͡\�E:�i�D��1	A��G@7�X}d�Y���Ҿ�[F��	_	oyv�Np��P盢)��-��[B{O1�Hu6!9�x���B/�1+etme?Dp�r�h596����y#{��b(Σ{�=�R��pڜV�TR�L=����߫�4�z����W�80d�9��R��ˇ���}�;qV9�{f`[j���]0x�k�1��ż�D��`qo���|���y�,xbH; n��Q~�HF�)zS�̴k�E�����*�h��SH�uE����Nq�stA�QxU�ER�=�Hjl��p��,鼄W����nm�Q��9���⪩eRƜ�ؑ��RšL'���D��#��і�����Xy���uko!�݂��ЖKK&��]�)�T��!%h�^!RF�1Mu����+"pp�k/8�+_��C���Rq�O�E`��g�-��P��gD�mu��k+b��"�)�Oѩ����Q�<����wiN�*�h��Aw������a�mO=
!�7����8KꕢI��۪��輹R�S%�}�H�.���Tێ����5������#���}��,&+��4}k�Ί��!b�ח~M�E>M&��p����a��ft��60���6!�v�Ӹ���K���-L���\���a�f������`;��]Yȇ����8���P�"��}�#\���O;/�����# 	��NX�3W0���*�$<�]$4���������kqϘ���N�E��lH�k/�J�H�Tâh�Mu���K���'��_���CbIԐR=��f$}Y*?ꗻ4����PѴ�!;¢�j�i�����������@߶ABwJ=A	�^�UOI ��ü�E��'߃��)(��3�z,`ه��h����ZŚͲ8��򲡇9�dX6�K]�� ��nthEQ#z���?��O�HR( .La��+�<&������]�[����cJEb�?V"Z<��I���a�	�W!�,��d%"q��ҁ�6cs~�}�t��9�:X<����?����'Ĭz}І��w�NmYm��}�q��}���א9��[�L��IWfc����opB�%Ƥ!�n:}W�����g@S�'��Bgw��t�>���p<��z���ퟛ��=�6\&��V��2�T���@a_��|��O�%b����)R
�qĄvX�w�\f)���%� B��v�������TP ��B]���,�lg��/S8 ;����[!a�C��� �C7�a�Ҧ*Я6�rȯ�3J�f�M��P�S��/�ƥ�s�#��'���X�2i[���K�{j8N�Gܥ���I�s�ϼq8*��,�C�]}��%�N>7�s�P��nm��ͨ�^����uY�h���g�K�o�~�
�0��Na�����>A��{~�j�<��Y�!_)�=���g+�)r��+y���*����|