��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t��"�>m���wr�5�@����X��'��-(�#W�$�p�.3/����R4Z7�k�N�5*����D�����.��.�UK������y�s����c�p{Y>a��$��*�+(�����������x$qƈ͆j�\���i�q��]"�F�8ò<bL6�d�
��-�d��������?�H�[�O�`��{�=P�	�(tC����kL
>A���0��F��ȝ��e1�W�8�q��4��$(��bf�M%�q
A�����-��:�`4S)bv�<���H�58��2�hS�5�t��U�m��Jfإ+�an�1��Y/k�?�'��4n$,N��"��=������������������r����;g��t��[/�/\��G�Ң L��o�C��pI[L��s�&��_#���)/��.�;s!��$ ��e�d2�K��F�/6}���{�k�~���]^a���4�fn�'o�&]��6������:����Fl�W���/2m�S�<���F!�uG��p�P���B2�[���Y �nM �S��,}�w�U��k@����y�FВcZ�r��9-���AzsS�\��bh+a==S��r�D��HMKh�	ȂruҧǨ�r%fc��ne&�}�]Q�M2"
�Tű�����<�k;e�H�n�)5�$����<�3������/{	y;eZG}}�����i�E��)Z���+��z4b�<ܩbB����&����hE��ڒ�&+�p�O���HR}������s������B���K$e�}9o '�yi�Q�%t(��Z����r�z�5e���=TVYv�-�3���S���k"���³�
�'��c�9xQU�#�ߏ�)� �#�i?xP,�i�[s�&8r�����/�����B�J=��7Db� �@W�-�찅3	f�^��A���w�{(�g���8��.�4��~�)���c4k�*	�qB�	2���2�+ĭzʭ�#��0��RZ�I���r���ة�2)����n�;����om�75�l@K��a��~o��{h#�B,W���5����\��sF]rD�PaÏ�`��	�]�:NU?���O����G�f���#����{���m"��G�"�Ş9�}�[�.���P�:�
H�`�@�����M����s=4O������vUF�c���9�6,!�|������X�Sy�;���@�\j��6 lx�|0��;t2����p�#bv�8l���ןT�LJ��^ż�{A�(�E0�9ts����s#�I���a�F5*�|�wcx�9! o~P��\N[��bV�q^҃��3�8��r�b̛��ؽt����U� -�5���oղ �+ʇ?[�(�^f��Q�[)�.�3��&�Y{���P[��:{j˘�
X�nE�hNT�)Ty�ɣ⑍��P]���Ūub����<��%Ynu�)^xAa[r�O_N ��š6n(5���T@6Aqϋ�%�L��\h͗\go���28{4>7�1Gu���Hd���:��1T����`!�קjC�$�����La)�2״!9��tّ�H֌���z!�:u	� ,
�nc���:@�}�2��toG>���v�_�t�V]�nT��KX�+YS��Gf:��^�v��\\��������|_h���<�ƼM���)e��
ML�c�cځ"��{ޟ�"4X���������1gÙ�zc�O�%P����<EM�>b��N����3m�UEU�~�=[m��@�{�;ܩ`Mk�ܟ�?uo��B������p�b�b6�x/�w�kb��H�Eg�FA&���7�g���ӿ�ٙ���ݣ����D8�#��J�'ڧ˕�W
����:�t-Ȍ$[���A\�ě^D)������u~�9D�k��S���@�B^&Q-��Ds��������!7��p<�I�T��Y�ݰ_��3��|T���,{�:E�Z]������L�,�`f^�\G�P6�TpOB3��o�ˇ_V\u䏪�a.���㵝I�0<O�X��3vG)�D���隝q����^4hb�8�;D+�3�yB`o,pcO?kjs�������:�x�ߔu�����癗[4W��E\t����+ �y��X��y���	�Ҹ�U��[%I�
�#7�bj�S�{>���)�����tJOxN4��� ~1z�0�b�ń��c���Җ�Pîh�v����?�����2��;����Eq�L.�M����z,��Lo]����l�\f��\��t�<oP٪��d��Sn��
#�$���<
r~���0��T�ΖU ~����t�=2(���T����k��m�~� ��C��Z�G���0���
��O�`h�1��&
�|�Ő���a`y�s�S��\e���a�Q �z�m�s��ٮҠ�8@Pm7�C�W��2���peek�6!gBQ�y(9��34ⱄ'�V�R�є~R�j�	�>�#Ubt8:�Y7�gE!�7O"\��<���*�&;��] N|�@_��GxY�b��[ܶ�����0%
d�l!�jgXuFUP������3�.��1�k�U�L�+��P�9�ˢ���0�L壔uGЕ�Y���ti��>4���Oo�]�1ـ������l..�����xH�/�B��܃z�L�@��լ`���m+�G>7���lbKq���Sٯ��H<^)\���������
��	���������;��ТM�YM�RP��j����-�t���������{�γ��ŭ�[�NXߗ(���b�,�8��s�!�B�A�O�"|�|�8�D�*�%i�J����W�d'},Y�}� ����E��ր$5�F8�� �]#�>/Ny�X��d�}�YBA��>��Z8bYb��w9�wA�G��G�,+�ݾy�ۚ�t�#�둻ÙzJ���Y��;���'ap>�O�C����6`���V
M��PH�(�e��t��P�!� �2�i�bt�{z�?�g�N6�v�B8;ޭ��q  Ỏ�X2�6��3;�3��v�8qz��\�E���֠`8/d��Щ�����"�p�& �s�i��E��~�%�fP��L@�Rί�R���ͼXK D�F-任���sEe&5�.����1Ԅ��(k�E�{���؟�,B�ԅ�k%e%�:���Q[�R�P� 냇�-�8�z�s�5r��Ͽ�����J'� .?#,8�'��*���ٯ⮩؜�{BN���~X�UB.ҥ��6�Ǆ�lZaRr��5��T	9c�<�N�4<���r���S搎�=C;�m�{��j���^�u�:��yW�����'�s+�kk�V��%�EO{����u>s�
]�zr�<<'=��J;�Q p�Pd��YS|6	#L�w�������q���y��U�./[(�l������Y\? �R9�m�W�2V4��*�&��lX+㜹Z��NZ�rkU�{[��O��X���ݜ�R>@D0%{rr��q��j6�%S"��l�؈OX�ېR����?�
a�xH`S���CU�,��Z�C���!)��e�n��b�4��5c4ݦ5���ƣ�������<O�zl�W�j�xa�^M<�w:��rԴ\Nzʀ�]n��ԭy�v��&��d�q��F�5��S�W�)��o1���i�#�s�I
:^�r�t��R�lRU����[��v��>)v�t��=�ڦ�}I��,3���l�o].υ?m��5X!e_�<ƽ4����S`bV��Aq߆���]Џ�aW���,�1$�E_����QÆ	H=���S��n-�=Q�ZB�W�֝V`�u���%>��.a�Y{��(]�Iw��./A�n�C����+'��ִ�MTȶ�qc��*A���aõ-�&�<��Vఘe�#:�|
pFt��2�W�1W�g�$�|�I��3�f�d�C�o.�ǥi���z�umN�b���`H'�d ��K�Z�^mS��)��l��D?nxn��Kh�R|S�$�
DI���g��5GgT0;s�����<�9�S�LXkKܛ�$:��+6q���0��A	�����&̸4ڃ@s�y�����/]L���Z��yW��3�g�涮.��{��#�k���MK[��i�=h�H�{�ۺO���D.E�q/��W=Q�յ5�?�����f/�b7��C��Xi��0b�m?�=Y��}�^�!���l:�_7����q6L�F<��e�ԇ��,�Ը[c'���^@K��4W�{��"ǿį6�[�;m`N�y�_�u܍��=�\X�G�GUIh���w[mRi���Ηbn����ʤyc�B�8�|x<�%X����J�SMR���l��4a��Z¼�����{��ʞ����F���=^6Y���%������NOʮo�����#����b���PZ��G׀���L�v+Bcp젩{��+m�Gm�4y�L�з��{��X�YuR��[�P�� M1W�'��*���D����Eu�`�N�@�����3E��Xn���+�vRku�L�b��菵Pl�(�_���"�S6�[��n���J�*�&����]����4{��nA��t]�r�<밲|��.>�n��C~b���O3��L��2���T��J殳�`���q'��ռ~� �����P,�@!\q� ��i'�a;0R��-n���� ['��Xx����RdH��&�뱸� aNE1*%�gp�KOo�Wy
rd��
g7�>�ٍ�t��Ⱥ�!�XAa,�������H��TT�57�_���Q�+��	���B=A�)�,q�=��q�n�ٺc���5P� *ѡh�Xy �.dˋJ
���-
ޠ�w��1B�a���?\��\7� !���.���8Q�˂.��J<
7�ر;��j�ҭT7h�Sr1���C�DMc�&:^�vw!�q��#1��^�϶�?�����U����l�S7,��3	��:�wN���BGR9�	�#@�$h0e+b_�Y&E����Oe�Fw����7,�l���X3��|����Z4��4�;��2��j��;$!R	V�Y�m �i�����!�u�*��P�)]�B�{uv�]��� v��Dd V񠹀
fٙN�h'#9���}x�r��hMhT�4d��";T����f��4�8�G�jZY��5�; �m_,<T:y�"�R9ڹ������/��7����$��LU͋d?�_|�O�	&��͖�ox��|7�0.��}U<�wM���5��y�s�e����o�I�6��F�j9K��ɔ�����B�8�תK?/��7�˞R]��I�����4��bq���rL����|�9B�c�����]������%�Q���M��/�����D�I�̿�z����5ݢ9XkS!��8�x�	뙀b�O=|~�R�ac[,s=`ުW�S_Nj��g�P��߬=��.kRj|S�
[>?�Tj)�m/��@w��H�HQ���--*�z=�Y`�nǅ�$J��d�6�^0���ܳ��w�G��ڕ7:xs�5�6#L�v�����6r�G���~��)���?������,�N����*y?��x�ncµv�?��X�<��*+�,�<���_�j���^�E�<"�{A����8�tָ��Ћ�.��8v�>��l�7���{�ګ�2Z�!r��D�Q���h}�&Ppńe�,}��
�����R�0�R�)|��{M��?&�5��X�Q�3>���Ik�%v� ��KU��'���U3��+�c�g��R`� P?��&P�#�� ��}��	�h�F������v�Z�%��*�:.�����yX�`�3�_x�=��,���2�+����AQ,���Upݻ�G�ʥ���|�1�'T��?dx�kA���<��;�t�4i����Z�]ඳe��.�����#E *�3�H �E�VC���)N*<�R��lk�F77O|�P6�r�gޖ��� \�=��Mm�+q:@��j.� �Ʈe%Y�t���5l������hL��?����	��#$��/��*��9�����sf����қ�5��� �E0I�~H�j�/U�華���-��O4�f����ɪ�N���P���Ҳn�31o,�����������æR���%�/C���l��J�l1_���Ί��0��
���nM��u� f��~ҝ�ƈ��704ՠ7DK�9�e�T6iL`h
;���L�	��A�tJC1W���&e��~�tz-���{�f�A'rV�Ȋ�㴪g����ć�yZ@�/Ro	M�F���c�M��θ����#ӣխ TY�/7�`��������L�.B�����A�Gs�T�<��;��E@ٓq>�P��ڄ�_��< ��6��g�I�o?�	���qX#1�K�y��5�D�X���/p���9���pa�fx�7F�IT�A'���6�J��X����3�=Y_��/s����w��K�{R�}��H���|�6��ڲ6��PH9�ߟMD��.q�O�20]����d�zS��"�j�KI �*�ߠx��s�Hލk�=T��.�M�6/6���}|ȹ�$+e9?/U��|�!_����5@'H(1�4xz]>1��j�	�͆�Sy�%EQ}>`��"�\k����FO�01��!�f/�3��6�l�cL�������_�ys$�����}��ã/4f��
�9
�x�mJz|�{��-e�"�A�l3]|�2�xs�x���S���^�t�0ov{��4o��َeЙ�7P0Fгn�%�H�����	#6�Z. ���*0@�x�zP$P�\H�V� ����A��qGT��q������5V��y�G�����#e ~�3��g��n�]
� �G��N�	h"9�'�]Seq�.���ݾ�S�D�*@Y�I_83�s��6��Ғ�a�J95���B쌱����H_o��c��r�}�$�%4�"L�V�,7��n�@�ۦ��t>��P1H��ͅ�w\~4�Л6��m�MR�U����v����Yn$��m&*cN����I��S*��h&��|>�֎<9��E<�����#�VӠ�TW�xW���-�}�g�L*N���s
�a�>�3�~P E� C-��PtB&��`}
�J�F��G�`��s�^ٺke.L\?�?:���$�g� 4E`{�ϗ���({���0$�y����A8#�2��.&����������U�NbɃ��#�w�c���L�G�@�M|�z@�9I
�0��D#��Am��^�]����݈ڋ�k��/��y�G%|s�]�ėzFJ��J`_:�����������*�h1:�v�ݺ|oH0����T<�/�:�������[j�W��j��"�1���ן����c���Npo�+Z$�*�o\��{��{	N�?�� ��wkqHr�����Fd�ٜ/C�A	��BR~-kbhl���ߞ�^�i'�V��t
ʕנ3y.�qZq]SM�= ��U(	Tm���3�l1��Ŏ�K�������$�9Ba>��:{�_�䠀��t���Ws�^��|TU4'6�ƺ1b��v�Ƃ�h�J�$�g�9�+9���z���������;M�O���r:��Ob�{�xym~��<N&�jܘ�J��Z��/B�L~�:v-g�"ؗ��^k
��	h���O���d�gy}~R�ߒji�/�^�La�)#��$v�֜K���)F�go���� �=���"@���m�!%7�P�vA<M��f���J�v���/hQ�j�J�`п�z8Ԉ/w7����G�}N�$ Vt���ܥ_
��
|m0���,ς=�I�m�j����*Z\�s?�:��+dᓼ���<�܍9���$��3������|-�y�q�v�ՄD��ٛ��*J7�}�{��v�(�J�m�"#P&�0\�ur��2���|���.��S��x�꼩ʷ�Vp��`2� �U��_vXܰ����"�^$�{�C!<�U*ò�gm�z;P�	D�: �DV�M땶8�ƋA{�$��+��*���6��uy�u�f�;.����cn�{!tSyk�v��`�6s�5oXI&���s:�ewhj��h+��Q�P����E�\�l]����`����𛭜L-�il���=�V76�Մ������J6� �8�݇)i����WL�zj!��-%�8��u҂3K�h���
JVO��#������0;?NW�(��#���//<۠@	�����AE$c̮��ƃ��0o�RQ�[}Ƽ[ގr�w�ؖ <]�%pd
d7�c�09EA8}��厮5W�s,���.":�op>�_�Xf�݂�����`ײ����h7�H,ͼ�x/��=a����&f0}Q�%�ՎE2�-/_Z3T���=#6=����DJhc�@IW�����Ai����k1�)ýX�ᮤ����@���3Y���$�,mq�p�v��Ƨf	��� �q]B��&V�#�Q���J�
-�^�d�b���Բ=�.=��6�_Kz���M/I�$��Hp��+''J⓺rnEq�a��@�jv�2�-����M���[�͈�qq�Ύ��A9g����5n���y7�i���V�Wu*����k��TY���TGQЏ�T��DTB[�q̽��wigk� �*5����$����F�f��j�~N_}�#'��\�۩�f��x;c_���f3WS��:���y]��p�"���Z���8%�m�&���k�'t�{}wIo���u�!�-�y��X��ߓ�G���ؐ�Ђe�|'_k!l�?%��49m�3BM19Ԁ�#ԥ A�Թh���"�aĹ�y���R
��X'���M�������}~7���9b��D�?����`��-ǭUf9�Q��QpݘW0�l�P���sV|��+��F�Gjt�k�}~���u��_Ӛ4G��t���9e��bwp�1��a|:���| �ѕ�a&���=�'C��bn��(�e�l����,)��h�&C_�-����k}�]I�-O�{��9 c������ԙI��CjJT�eY���$�J5S)(�t�d�Dz3:c_9�H��*|ըL�d=`knK�<��]��8 �z���D9ŰSdC�\�� H����O�z�7�CU�/U"��qwȽ_:��J�,�n�}���4`����g��T��zEXRa����d'O��`�;��x����#.�������N���Y5QV�/Hr�_z-Q�I7Y�ڵh�S�牶'3�pa� ��[V%3��%�����ǩ�~cri�顠����q)�p�N��Mu�{�^��H�4u�홇�X��Br�D��L�TgeG�1� ��ZS�t����c�ʽ�5�&N��A��|ѾAY��8�	 �����Zu��?)u��M�M�Qsd��ᵶ�����@�s�wid�����.�((qj�T��\6�-�	�Us���&f]��Wm1�Ł�f��;�7l���MoD�;�QoH�i���P�Hn��J~������<�A��D�j�E&�8q}� n�W�ny�5��L�L}t���M��yP���'�>�T�7�f�I���[
Ǝ�)
������D?L�Ds�y�z��!���d����܇�5ۑ�u���lu�/���X�_�^>���j�fNz+*nڀ���d���}���9���i����	9`�L�.�{o���U?�ܿ�%4��"ز�÷oR��QDЗ�s�u�ӗ���9������j�ۼ�Q��C
�,�՜(v�����\�_	���PM�NF�!ʠw��&��.�b)}�|��a߹�ޢ�#'����&d�A�)����&f�W��@YN��ի�p �,��M�"Q���B�g(��N/�P�:t\GT��6y(�h=8`GZ$LRq���,"���ų��=o�v�7���/�(��C/��I�q�f׹@�<�G���Bl�̔E��0���Vv%��B��_�9�a�k`dC.E�H_�~�I��!��8�|�S�3݋��MI)�2AG%��p֞��ɒ2Ys>�x�%x�7�n�jm��)���,K"Զw��p������ t,�	#�F��U#��h��l/h�Lx7i���ì*�1����;�.�"C�~ �����<w�7�aD���U����á�8 `%�y�Cb�Cy7�nsD��m���Y�C_�g�+u�|S*�Dh�ʉ:��z�Ş�5e������S~�dAt�ٷ(��S5��d���f����ڑ$E6�U�e�1}�Py�魎�G��4�O|X!g#3��,���9��Ӿ�a��p��Җ�A]���.�_���K�G���t�#��"U�9\���_M`ѼړQ��7F��~�r��s�#�c��f!q��֛�[\���s$7ɫ�@]+�۰�'I0k��4�v�;g��Hz�D�����<�q�Ò��"�οu�:�B�u��kv�k̰����`�v7�X��+�#a�Hd��X�b��c:FX��N���w��@�U �åW���8�~�RֿY[�I>�s���ܼ ���/�� 1�+�����#XO��|��j�AbB�������	S)���s�GJ��mg�k�)(~�j�H�C�`P��ʒ>6w��_�p�<&:��b
o�?����jeh��<Q�������9���ss��ha�^��,2�`�������Ql8JbМ���'#��`LÏ�0[d0�*n�Q�Mh2p^�����_)��J�DpCI�\fc��nr��O�_��Է�D�]�ڱׅ�,b�����O�r$�$�}�'�۟�Tr��W�B,-��L�/�uk�QØ�:�IB���L]*�wE���.?F1 �%ê+;s4��%#�̲[���װ��O!��6e �V� >���Xi�%�A��|nE��j+p~{C����d6�kR���ZU���{c^�p�fy�� ��H��/�����a(c;�����'��P�J)�p�:+JԾ3�SMq�?R��g�8���䮬v<�GRz�T�	���쮪�(,�0��?��O��Qޢg�}��n?7UKa�`�X�Y�Tϼ�q�׼~��qZۅv�_m�q�N񞪋ҏq�C�7܌��J���?�k�P�H׋I���^L�0�=�RQy������7
H@9*k��J����Ar���I0��n4(�}����3��N����M�����-U�g<�5���CpF3���.���] �x��_�����O�i�-�)��QRMe��c[��`09x�E�bLQ֑��}~>�:�SN�p�$I�{d5����+^�{镹A����y�(�0f���=-��9�7��Š�>�؀�G����B3/E@(;�@�~��ys������ׯ�BU9��A��1)�7����	��\�`�+2Z�lX�	,:��c�5����T:��y��Q��J��x��#��'�y�`����CO�`%W��8m>QS�k��I��q�q�Ư cG�#$a'�+Ec�s$�8=����u�Y���wa�L Q��+����"؇�����}��MR��D�+���ٹX$M�e�_�� `V��!\E}K'+&!��מ�r��F(�qU�_���Qg�)���l�ꆖæ�BO(�VK�+_�KO�w=o�14�'���`�b�#ʴ��3����� J`Aϙ�R'UtC,��̂; �&m���>��VhP�W4�p���GO22����N����^�@�J�Lc���7�g���WH�}��A�k6��hX�4��+����.X8a��ʥ��'y��  �};�wo~9n�6�f�R��rz-�a4lp$>��C���(Grp�LT�A-��#h2o��'�8NHzR��$���"�zŒc�#��d�5�1�GWbo3���Q�>�M<E��Z;��b.7�53%\:v�� �⇦�hb���T��H�똑2uR[Q�,(�D6u�IO�ӶG��/����Җ\�����D���;J�����T ��#r|%�!0�P'+����w9i�m��h�_��t. ��'H���Iq���T��������89Z��O�Yb�]l�'A%P��|�S2�`��U�s:*%Sa\W	�o� �U�����Ǒ ڶ�}S�DhԄ�^ �_ǈ�^��Ѻ'}*���'�}�`e���C��vRH(��֚�C�_���K_�oWt���]b�Īg��r�^(��^�b(�s���V��R��>���Ĥ���7�B���*��&����5�E���Q�dΈ������/�r���9#�*�'a�?��F���o}{[�VX(��`l�Z{w��
0P1�N"�v�߽�H5���;v�~�>�����)�s��E6T_���Dh󑬜�i�����T������⧲Qi�e�w_�C�5�-\�t��n8�f��eȔX"���'�O?i*���]��x:�ȳis���'������S�|/�s��s����n���>�
ލ{cT�)i��s;�p��Ⱦ�S<�̚��hk����d�VH�&�m���=~],,Fsf��م�����f�����H�O�.�<"ZhCΐh�5�@%�+降+u�0��睾}8����&�)x���Ŷ/������ͫ�OZPl)v��"��`}��/FբC�fB0��E%��/H�S���yf�ǥ�%X`�9��T>上AФ3!0���t'Uޒ|��z���0��f�����Q%*�x1WQQ��L����
�&h_s��Z��\�s�B_�6�%%S��I���%>���j4�z
	ս�K|z�i�;�U�}3�(�A�?����?+ ���Պb����J[��v�a"�O��]�<�d$ĝ�>�#�2��\M8_������LR���(��f�)>��ۋJ�*d4�è��u0�"Q�{�� /�7�e����ZV��/�i�,o��qY��k����&tpwU�?�Z�>���?]>�B����}�+��וЂR�0���
A$�k(6mLO
�Ӎ��l�ak�ǱUEv�����$,  �7��܌�L�DVd�G�1�l��5VL{Ht|��c�0I�-����\� ���*̔�:~~����=k�>�w���G��SNw&��JFi��	�Q�V���
u����r�7���f�o�3-�΋��si/e��+�� roC�����8鰞=qF��|Ҥ����7�q�!�?��V}P�_m�%��Mļq!��uk���:M�|����w�`���Yb^���و����4��l��"
�ݜRGm'�=�ː��4��jc0��zKq�	.��o�:�D��)?���!��)Cӂ�d	�۹;4���#;�69���_0��ul�0.���wgmx(�hU�z��&��~[eTy �|�q۔�K��8� ���"�"ϣN�)V���P�GGJ�R����3]yD���C*�����1&�c�a
fs�b3�Ϣ0=[���~�(�~��	r��{�� st\�u�ϔ=mf��6�BI�8��aGól���*�hW!Ⱁ�Z�=pd��MC�=���	r�����pˍ@ApN�I3v���)K80^L���#�tr��\����T�y��A��Z4$��{���Y��>Q9f �������)�U�;�iB�4k9�����z�Eq�yM:��v'�4��(.�8��C����y<I�q_�0�_����PEl� �֤L�(��r��
�T�j�-%]�����6����v&j��h��%�lϥ�N#g�~Z�#P�36(}�v��^ol�p��w�q&���d�K��4���ܗ-EČ��+A�g��|rf��28UyCp�Ɛ>�deW#!�V����LL��~7�������]���m;  �� �xNLV>��#�yG���M�W��^�m�e?�@u�M��|8�"��ְLS�ʩiKLCb-_4�-�su�g��$�����ћ7(��j��:��!I-�ޒ�f��1$V�Fh�2���Jw��E��<��hW���6���/ϱ��
Ҽ VG�y�R�����Œ���|3���s��P�k �%��Scv��4(�-kOD4�2���E,�d�OO��~�����^���~X��I��!�a�����+�U���<�w .9�Sܟ�2��K�(Cd��o�����Y�I��w�֓��_r�;��#�Y$T���y�ROx0�]�����	O��� ��	-[�������7���*)����F�0Qb�1.�rS3��bM�1�<\��3��cn��g�:�fr���M�u�����V4#�B/Ԫ�P4�k�]ݲr�_ȭ-�G����_J�����N��Lk����.Mm��b� ��:-�����G�W�m��Y�b&�
��5�.'�	P�8���+6K^~-�����R}d�h��� w��j�V�<"JR�(Q������L�l�e%����ae��̆��>�<Q}�0PfH�_-�K����DG���o�"�\]��Kq�k	��M֮��I��#F�U�����]M���Op�
%)*ю����
����e����y̗@yY��N�X����p�1�s�R�Z5�zL5Iv���ຫ��vX^k7�B��ȯc�d�Kڻ30�����;�{�c�MQ�!�6�uyUX��y9x�>$�*,��>�*�{��H�Y4�No���y�9��o�mHFV+Ѷ��jɚq0z@Yi�=��=N)GL�Α�gR��S��oGtk,�킶�bD۠�/������_ �:����Zr�������i����#4�z!�;X��J^�3%�<b���0�F��2����Q- N�m)��s���7:<�	<x��~$�d/�*���̨�24� f�C�u΅��Q��-�9o�YM���A��noAQ��x�j=҉�s䤾�̯nb[��,�F!n�o���M1�o�Ki9��|�c��|��O;�})Dؼ�!�͒7T�x:M�B�uӞ��]��d�Y紆��X^����QnJ�*ك�ĺ@��W�*�2�b$.�HW��e��i��>_=֊.�#�5(���#�vx�B������L"����|O*R� �[B]LpJ�N&d�sGn,��V&�ӏ���6H�Ήu!;����ʅ��x�ٜ:��Ju�SY��,�K�v������;e���s�l؈6�Zɘ0����'A�ⶉײ忪D�����
��3,�n�✼ݻ���(�����M;�?�-<�`�t�B٤Y�:\�򒂋6��
�L��yR���9?J*�A�Ҭ��c��|��+�����C��|�<���u�T����ާ�/y��P5{���Z��WLKW��ok�� �c..��:w�2�V�������9���R���m��@ܛꯨ���S�!�ǒJ5��gmGv�uXs�~�y�u�D���k �ӟ���1p�T�'�'q*�]^���=;�ʱ������@P_6<�+�]'b^� )Y7�APƙ�</ӓ��7� V�[!�c"�h�'0�>��~X��l����28<:�K>kU�+�kN)wBԓ�y�^��ng�H�%8����yo/�����do��`��"xzu�q �.��
���^1F�Su>+�\�G5ԥ͝��nϬ���X�/L�|�}]�6[r�9��]��]͘���y���H�G5�l�Y��_^�^ ����;����e�g!�'�C��BkLT��x.����乳�*2�iqљ��CJ�
uD�躁�,q���I��?�Q���$1i��|9�����FK�{;y)�С	��8�%�%�^E%�:�]W��~�[� 7�c%v���r�v�*�8�� 7�� 7,�F����-�{u@X�=7�zc��
�]�)�p
�`��7ȶ}�`3�E�eKG7N�P��+ȿ����ץh;���Ü���SQ�5��?���S�S֟Jfƛ�J�l|���6�ώg��J�^ɵ���y J^���S��"ȃ+�hq���I�0p�k-ݏ7�Bs�����
nT�py����҄�A�#"��v�u�HX!^N`aN;���4)��nN��'���yF3�(F&��EŢn�GM��g�0ɿ�x��g�=�0Hv��0�[�إPXw!����������R}���[	�J��GZ��p�&Zc*=��7�F���� �q� ��T_��=@�-8@N~��T�T�5qo��5�ai�1�����Zg۠�l�b�i��NUS�T�����#Xcf�����[9J\�<J_5 ��P���¯1x�Ԗ\��o��f�p�f���쭮]i�6a�^EH��9s�`je�R��ј�"*�C����,X���X�nA��pu���`��XI�x�}"�^��m��mLnM�$������ :��`�\��!�Y^O�lR��*�2�u*P�b���~%��{Q�sT�PvDw���k�g1^1@5l�9S�o��ViC���"�\σ	�Ъ1rp�{��9.A�J>�ܦ�j��(�u�3p�%�^�����&(u+���O�w|��8՝�<#�'m��Ɲ�������:�401��!�dD�g�Szh���x�/��g�:8{�b� ����[ũ/c㢶���e��Jy�`���Q�Rp��<F�T(	dNG��Bh���ҿ 
���3\7>vL��tᮎ�5�E���!���+Zh��j-3�U�J�KӶp�A|{_�P��`�ϡ�m��ֳ���ak�b�8�� ��Nu�4�wp�U:�Hy-y͙�dRld��03%:�W���Ԃ�$�|��q�B��޶�o���YDC*��pf��E���ޒN�A�^Z�ӧ���!
Q)GKm<����$������'�5�)5��	��(@{?\�;)�3��O:�u�bQ��ԥq�S�>�����rH��S�Pݢ3���" �I�(��Fm[@$>!�_���j0} ��m�H=@�`���:�;dMol�/,��{�12�����6��uB�������ˀ0�����_ڹj<�IG#=���R�z��!|�nr�q�����=����Ūڟ��".��u,�m���2A��Q3���IV�2��p���N�|�k���;R<���
�����vFd�S(�=��G���.�)���F����ǜ\�dmδ�%/�0׮N�^;����骕%lW����8��E��H�>f"K�[Nn�~��Y,�~�&ZCd�e��9
Ie�T��#0�����CfC���J�|\�4%����O�MU�zY�1o/YB�c��	�m!���Up�Q
CS@����\�$����묜'�3}��[Z���;��W���S-��v.�|M}UB�m`��յ2W/�����wW��lx��^��WCH��ٳ�a��:w`FE����tRN^�ꕻ������s��v�t�c��`I&X#���0�X�lnG9A�8N�j��i�]3s�����E�6�Ϝ�@���$�M�r����C���|���&��9���8p"r�%�EJ�V��e�A���rjl��L!���7Š��٭�P�}틿�Q	���`���wy�w��K#�3+��?q�Ƒ�W�͈��Å��	�(/=�ٳ�B�T�eqڲ����`oW��`/&�a��������nx��������I�ae�2G�G �u�^�x���v�k��]ou.3CQ�i�?	����`�q�rC�RR6���]���7"��`� �ȧ�g<- }(��Q��^�)�����pH[�_p=�g}/ًeKs��T��\|3�O�+��_˞����6��T�G�ǾÖ�Q��MH�K���`�	�<g(آ�	Y)<����P.L
����7iK$KB�V��"���â�_�fAc����Z����.�5iz�r5�.Kx#�6������=NCE�l�SR��𾒭q&M��ҹ�v����\���۩Qأ���}�i�4ꐀ(�*h}�]ə�������f�Sf�Qβ=�t���UGc���.T`�~���!���8?�"Qx���L$]l6�B*�AD�B��� pQ	���s!��b����R#U�q��qX&����i��c���||ɳxG�>L�J<n�)B�4���h��?�ژ��a&_�^&�_�٠��>��� YR��à���[�e���Њa�&&H"�9��*��u�y��)�����S�ni�sU�C��Sh{�F�쪁2��^3��pQt��5Z�����*��@Y����8IK�ef�A8�u����M|^������, ��T��� O5:욑�z}q�w^�a��9U�c�r�&Ӣ�Н92	�5�/JY۲ځ;�+L>���3��iĢ���Vݺ��Iy+�ii�Gw`�)ǰ�3wx���Zv�����,3m��R�y�0'����w}�M!�����-XK�o���%�F�>�%T���-@�oA�m�M�K�P0���4�2����_w�&��3�ﬃ��!?�~�����)����xV�+�@��vbɸ;�iv5df���@n����Ӎ��')�ߏ�͎�6Es4Q#	U��i��L�-�]]��^s���Z!�!�Q�H9}����>B�m�0��כp%?��b���c���V����Hn	[�ͮ���F��FӶ4���@���z�r|�x�Dp���>��Z�����+O�G($&�e����2}E7L�8ތ�[q�%䥲�%�0�@�����Sys�w@3d��]�؇GV6����i,�f�%F��Q�
_q}F�U�ɚC�z^ٛ�{"cz�y���-p�Կ��	�&4L�[�}1
� �5F���
���+(�Vn��A�Dxc�k�pI� ��PW�}��gb�yF��W���p���g�f���M	7�^�b�ܸ��|��7Us�g����f��J+�]�!{��ӀW�m߬�-�M(�.*!�Ϡ�#}�n���*�|�K�?�j����h;�Lx�&���=[��,�Q��L��cĒ�|�ʷ�������щ�&����Cj�����Jʻ��9#A��B܍��u����������Nl\g���a����gL���c�^���sb�W��4�$5�s�ܷ�����������s�m��L_I%��Z���YU�y�df�;��X�Z�U���aGD\�H�N���򢉹 GE5S��78U���G�ť�mbe�;����Շ����E��ZX�jP�F_��H!kj%�����Kt6�a�-y�UC�������bE=���%S��ï�H����)q���YCܰ�bY���o�l�k���/O�zOW�tt�̌)����=��|�:�ϭ}��L�>�F��wX�!|�� ���D���c�r�x�.F.j���b�)Z��������Ҷ����0:����Պ�X��`� ~J�A���_w����m��n�PH*W:��'�g-3�$�
�t1XT�I���20��ۮs��Q���[�{o��\2v���ko󼳭���B�z���gg蕮��1�VG��׼�~���lv�o�Ʒ; �h�/�>dSkѬ�T��`1F���gh:�*}���{��ު?b�Os2�p�ZS�#���K���%
|l`���]΁�9�2:��k��łt���M��sZ��F�X�X�q�\�.`BՔ��Z��M5����e%^���ȓ����+X�#��������,e�y�#�\��4R���_�v�����
�e��o�gم�\���J2�w��Y�ۗ[X-��]��2صf�TS��,�8���}컋�T�:�$��H.�*�����'CNK���mlןa"Ӆl�&r �h�
�R#;DJ�{j��z,1��ֺ�F����f�\�^��9�NfiP�ղ���6O�����NCfS3 �oZ��QA��}B ����Kc�E����\�����O��}?^xD(4W��: �b����l���0~�.�3.�.�[��|,���������/:7�)�.�s����r�NS4��w=�j�m6���C�
[lLt0�e@7'�� ��� ����X�Jse�H8�;��Iz�� )ZMB�4�,~��h� �S��#��'��q$�,�o�j�[�$���hx�<.��]ͫ�A_Dk����ٮ�E��n-P�����I�}�*?�e@��j,8��J��E�9���6!U}d���h!,l�'@Z�S��܂��+�x�M��O %j�a���@���Lo�7h�^�w���~>E����yQ	o�؀��xO��{)Q�[=�x��yQ3�Q�:�?����,�!jy
E�=+���pŒ�^(HK Ǎ[�#�J�M��E9'Zt74�7�R|��u,��(N�Ԑ���7M�#3�M��Vu�a3�a�N�z��)222��Hc4N-9؉V�y\���5C�G�^�@�N�#I�q;+4�n� �#���s{�l�G�Ww���"|�����/7b�y�+˕�v�~>)�{���~S�����6*��g���!g�TwDڏ73`���x�W���(	�(����9:SU��������l���ax!Ґ�x��"Xܐ�i�yaڲI��Z�n�$�ƴ���2>��k%#�� N #;���J'?� ����s1��0�G�!�!z���%Ux��=�4���-&6_:d��Z@�4U���b��F��GVu��wѱ�e���k��BgI�I*�3���&�=*L;�c��+#�"i�;bw!j�}� �n&�Ȟn��^�0�3��sFvlrs/��T�*�1ᇞQ�au���?u��j9_��$�e&/��%�j�0�6�=��l���5�0zDU��$���ɺn��j�1ʚ�:��)¯�\]c}�g���zm4l>6n� 鋄�����Ų����n�)���u�|�?
پ��0ƭY,���[T��ƛs�m3�������&<�R���m\*����_5�9�E6}���s0�Jҭ��v�Eظd�SEX��.���㽏'��:��������2����8�V�]٨�����N@\*1��h뾊-���@{*�mr+�#i�{K+���4	t�*�9A��	~�z���o�<e�v&�L맋�2@��{�����vn�l���SD?{�k�Ja�to�[��Z*���2*:E�S�����8 0I�^R53���F���'�
X�\M�ᡙ,�����H�~v�8��S?v�v����Kd�Ax�~[�g{W��é �q�2-�Ju��a��+�_�^���w�w0�󼷈�����3�Ek3H��b��a���PS5��p�v|Q3���'
��6I���ܞw^˪p"M�<�٘0C��y�d�o�^q^}1������k*�|�¥�5q2a#b�6�=di��CE���݀����)�U���B]���G��[qĤ�g�B��'��0�j�7�~������7��%�H]~sո�6�w�"w�қ�������I��Zь�{s�
~� $��
�9��~/녺-�q��D~�����2e�0F��h��͡��1�m�qF�a��O��H/(�f:l�����#;2>,K����dp�Fbܒ�B�4dc~�lK��{p�K�����lĚ������f�P��1y���tkK���̃
�}�S�I�N1���{�/(|ra|*?p�UG�t|/��&m|tC��C&�33�?.�0ʤ�XH8o�x����� r�@�4� �j=��~e*ʠZ�yFYs S!8�I�J��c� ����ڗ��e
�f S̜�P�k�H�}�,�n����P�=�h7��X���ɯ��B���m�ۀ��)Е\P��B�������9{�C��y��k�)�(w�t�y=Ml�F L�\3!!�w�$Uu]K�$������')�hR~�Gy�rFW���J8u����K+&K�>��TRjŨEO.�{�Q|oX+xp_��75��t���@�(�#��CQ�,|��*7�D�*9�/���O��.�W�WS����� �.U�����@� �c�D-�ϵ����G�g� �8>p��2��%�ޠ�\2ŭ�m���V�����u�3����܃Ռ��w����]cJ�4K�OKf��������H�U��d�#�	����o�0Me�`�,C��3 Q�Jp�D�e���<��e�6Bl?�G�I��L�;y.1�>���'��M	�R�_P<�y�Zo�H :.������x���Oެ��1Z�G�a9�or$Ȏ����'.N
�R^���Y%�%V��w\H�yݴ:^�ᓍ�z ��zv�����z���g�OV�8�>n�|�o<*:�IH��)�O�6�?,���j���P�U*�b�H�(��7�!=G�ާ�q3���@��/�$v��7�{�AnaK�	�H�9P*��]iBQ����Uo]�SEB����[�h1ܟ)x̒x5	k	��U��B{�K]�>�N���F"�|�;q���ڪӦ/zE��[�Լ9��H�NV-���P+�?����.X@��˸�kٓ[��@R땣�{�(炆e����cc�I������3�[�(I��ʬ�x�h&����|X`�A�0�"c�IOX�z��EU�6/k��C�ϳ+tr#��ޏ歷�6�TJI���;.X�:Ux��� KhP��J�d������w����\��K�&J�~��@���׮���(�r]��&Wk����;�6�T.gξD_TD\����/)��$K��'��b�2����r�~��5��}v��IY�,i�ΘI�f���a��#�k��+���կ�M5)��9��:��Z/��E�PB�@�B1��t�i�c97�a
p���X��-�NLBD��C6wA$����DO�EtK+3"Ă�����X�ԏ���N�g�:ٴv�=��6R�"�7[��t�6��&���[u�t�l.��D���>v��� 
K]�pdca�8�T
����c2|�/���Y���g��P��58Gz�K�D�-�B�m1����V*��i��bX5]]���-A�`E��o6ދ�
�~����E��t/�Y�t�L(�H�L�ք��m%�q���WZ�%=�Ԋ���rR���.G���V4|@�� �.�6H��1v[{DH���e���j����+��wR�qY{�,4�t'騩 ����$˛dd�OFiQB9�L$�r�Q�9����hkay�짰��H���zD.��@ 9H�~�PV���/�tӒ{A���s���!)J/a�Ԍ
K�{�$Y96��j�p���0���T���fe͚9��ݬj�;���5
 b�E�ٶ�>����m��a['-�9�n�`���aR{F�	���v@#�C"Q����a��|		w�gh��u��?�D,";���VX6cU_���=6��_��@���H�Z~�F�Gر��Ty&�Ks�CwK��:��N/�	xW�I�9��O�k'�j\��
�Sv}#�@������b�qRD�VS�".�#��<�����f�!�X�'vg�ۤ�#�{B8�3U��@N�<�B.%8�ދ|+��B�e�?�z~��u�-nz����o�婂_�U�ַ�C��AO�tl�f�,���������g�/��]?R����t�؜���2���w�:����%�2�r<��01��\(��٢,2[��q���,m[�Ke�)�ml#F?�S觽�%�`��z�>HQt/��g*;L�$EN��`[P��\���;��l�[�:J�ÈE}�{��� ���ۢ�ڏ���^���P&�I�{�?�D�Ԅj	b����!a*`ۡ�Ut7��辻�&������ 
�P���'�q*SD5{O�8�o������0���!�Y;���Җ����W�f�oV���$�eg�Z�:�#1ɷ�9¼�9�$����ʋ�9�@7���>^?�`p��-�oK��܎S-s�c��B��{��� $,���5�i�����k��qfIi�<��n�L������U�w|F��ב��o����\52����{a]��n�=h��+�/��l��,2����iT�L5����Ң�V��~.����z� �*�u���pt�����
,q�V��R���S��^^�ץ'�W��7�~��دR�%�V�N������'� ��d1�be:�g�!�g�qE?{�1��؅��_���^�ѐci���u�t�k3�A/IQe�9�tk������A�{-���$n
��X�Ъ=k�+���_+BP 4�	u�O
ABuD�5z�"��q��`����у�?�S@yDtn�q�?���}Ȼ/Ӑ���Ј�GdO��l�EQ�R�&��{1�T�����5�{3siQv6
�7DUd�Xoo���d�����T�aD�F�T5���_�39�tE�7��[�7����>��<]=�% ���,0\�L�>�!మ�i=���������]Q2��u42\�ږ�V�i�ǟ/=A��Vۓh����}�䴙� �� ۼ�]Ac���^{!�#�|���l�}$4~8�tॢ9	᭤��I���*[�fV�:�.��g�;c���OWfMg�q@������Eyހ�e'��>��&������i"��v0��7N¯O���
c|R�#IW�N���v���1DǾ"xĠ��S����Q��Ů v77.�DDQ�re\��
U�@�8ќ9j��i-{��)"��茐�.|0u�]0��"(�NR��f���YNs^E5翬���<_���g��!.���������H�T\�4���խ�z�̩~Р(]j^%�^ ��|�� �Hr(q o�Ҩ��؆=u��������z�d��0��Jy~9��g����w^�9.N��
�{��4ְY��&�������=M=+ё����D�g�raJ;���S��s�b�?_�e[vE�]�	R���ON��Ufܒ��C���Y���ޞ���ZA�i��c!������MXz��� ܺ�V_���M\�a�wU�%�L�O�;�YKh,ܧ����H�x;u�_��p_�ws��)C{� ���� 'i������KYP�[��{:��-� u����[�op�1�Tk�|k����ѯ<���������?�x�=t8h�Ǝ��(����EݼD%!d�"=�ٔk��d�V�`tb��Ѕ��a��큷*˕���k�E�����x&���,浐u�:��$��Uv�4�����/[�xǣ�Q���:c��Ʃ���A�N�1Aim:'��!�rq�-!����vW<�.b �����M�^��R�0��Hi}-@-�������k�&(��m}�ԡF�|sI��)����7�f71�1���S�?���k���MA�@,	w?��z��!T�I|O�.2InA����Rư�T��M/����r嗵Qj�ܶ�-��U����N$|Dq\���#�Yu�Xš"�\�o#Vu�O������v�Duً�G1�[%/�Y��|�s��j��F����g2L���g��<kؽ�rr�I�o�1�CؾRÃ_���y�C�3(P�]���;���Ō�e�a� ��ӋA]
"�n!�w\�V���Z=t��ݙ��{�j/۴a�|<@��Y,�y0��T;M���Ƨ~��m棑O���&�>[���j'j�\7���2���.{1S�?�}�	��ve��:(�Ω�|7��WC@���ɩ���t��W��(����!�c�|���uL�����d���#J����'kN�J���p|BkS'
���\Ǿ�3!!� D:�I�w^�d�M5o�:��*����1{�9%i��S��~.�Cu�&[Tv3�۽ֺ[2�aD���ȕִ&��>4��Qcq�}u
�)k�����_��R�C��ug��@:�GP-�q���V�m�Bt�}�����JM��1f���T1N|�yc���۟�@D���޻�2�P�=L�Y��0�`QރD��7���Y��/�tzov[D�:=��b�wg�jbq�a�����N���D{�'Udx��&�@�Q��.� w,)�{�%��,�w��4kϛ�4�.�]4�QFd��`���������|��u���o�3 ��-XB��������w4�<+FR�n�0(��w�.�؃\����Gi�׊�D> ⭷���ԛ�C�!�>k?���[�����˽#���V��e�89[�,0NФ'�,�X{&�z����^��I(�oo�+;Ι���TgB���� �b��2yH%F���y�8��.������PP&Y/���T� �V���p��݉�,��Զ�<�9�`�F�j:�yM��=�� ��	�wR�>W3"��J)1�A���)P�o�@H��~~�M4�n��f�d��Xa*�A�@��X�\D���(UĶ~�e�r�a�KI���r�Zꖭn�Dq^4��غ��)�$-t:�l��s�Y�o�]gI��C�10�IŲ��SYŎq�;|kg���i��ޙ��V�@���Y��'O�x��?���
�Ghx,pN�W@�w�" ُ̀+��	,�ƨ�~O���#�ԋ��9yY%,����P5!z1�a 쀲�
3�<��-F��D�@Y���6��_ui�8W�a���&xg�Km̮�5F�t�R��K�N�2�:P(��J��� ����os�0�1;�3����zJ��T،b�Ι��4�R1�:�7��Ҵ���� ;�~�%�D��l=��J"�,�{_��.��c3ژ�Q�!x~�1k��Kל�?�pפ��~L"VO���L��t͟�H������m��j�M��|�t*�Ѭ8t����B'`wp]�+Q��5L��O��a�>��)�Y}�`��Q�3�n
8��ި�FO�_��	�Ҁ�=�5J���������ar��87�
 K��b����}�*c:e�ս�O��$0%耜UY����j�]^{�FO>W6`��H�������g�!�o�Vh��3�W�&�{�̽����+js*�W�����%��sq�yU�$KB��V�dE�ڭ�H�֐GY^I[�i��o��S�ms�V��P̀ڌ�y�\Nn�*���}��>��0�x�XQ�G������OG��x��-�`��45����M��Ȧ!�+�N{��ïz6߆�Wp�a��`>F?��ph0���Պ��� �w��	-Kb�.����LZ�'4�T��W*M�~zҏ���XDN���R-1���^����K&���բ8N.�|u���&�3G�H4�@ƒ��$���ڙ�{��gP��17������OX�әY��e��鱘���-at3��*h�E��`���>�G%�9���ח�$d^�O�̌n)�rMp��ͫ�]�\jk�]��)R�|���X�L3��l�� ������nzT�����B�A���	O�g�$�\Y
�+�f��͢YDy���wb�2:sÈ��X@���gi @5��,B��	r��h��=����o��y�0H䍭��Q;�[`�E{1�EI"�"HA�jV�T�����,�
�窔����CG���?�)<�V�'��ͨ7����JL�F�0PL�>�d��
zp��e������<kw�~�2��7�zL�:˄��ਖ+��;_o�p�p��1���İ��O�(e9rǣ6
?7!���&���~%$��"��Z�9��D��3��M����1ǻ_;�C$�8o��sF���~�m8����9���~�N�D-���x<!�a�@�DY�(>�\���&��.�{a�8 Z��c%���)�^<qm���*�ģG�lmm���j�;] �e�k�)R4�&����VXe	��|�#��@����d/�&3��-c�� �
Y�I��ѫg��r�����+�/�IO�`F>g�'�͠ f���`�j��T"x���j�c$��v����j�
�B������!�9��N(b�:��.�=5��stbk�p�ogˌ�.�aP�	���o���շ�^UԊN
�n��k}����\����B�ql�j�M.�h�?͚$]���H�%]�t,�0�v���ln���M����P:3�W⑌����Cq}j��ὢ�o�{I(�2�"zR#"%	w��Uǰ7�;��~���	��L�;�e�T�h���9z�'�n�]�t�����>�R+,�S�=�5���nT���z�������Y�9�g"y����(q)T���I*[U1���Xl^�1ׇͅ������ٶy�dN^n��/�C�lR��D�E��j��a��/�����6:�4�W�9�$��cq;gʲs�񯉫�t�TAm"J;�W3���XLӟb�R��K�Q,�%��t�60��~j"pBT���n�t}��z�[Y�W �V�u��9����x��^���h4���G~6c�ix��Q��SNܱ�ko:V=xu��*mʰ��ވ;��덼�g.�;=�&�b�#4ϔI�c�C)0e������zb�K�UZ;��10����>�����	���}m(!�,����iǲ7m���0V�؅v����4�W?5��e5�i��\"'����/PCα��n��^�=��;�`��D���~�.�ؘ���8�����hs��vFQ�}�P\K;���<~��e�J��]��(�z���\G���f��a�]�/�0r�ZNh�D�!o����7���;+�# Z<��������Jl$����À%��C����5{X�@��R0<ed���P��D=[a���H�#P"]@� n,��e#����Q���b���?�Q*�{wl�9�e��af\ըh��R�r�53��%�9���9
i4Lu�K���ȓ���"�e�����,�5�d�H��7v�G�GSߥD�W���ݱ�T���	�B���䴖_����F�S`�ls �р�A������!�_%a�8P��e�/�׈��a�Ÿⵧ�̠k����]�D��]C�8��=L�#�	G�d���,h��m�aWڱ{ڈk�v$"��8��hz�d�4�1�Ň��r~��BT
8�uf*jH��LK|2�����mĕ���ُ�D)Rj�l_f?2�4.@��#�_��~���w����PF7=[n0qNA.�ЬÍ*H�+ɦ�J�߬HG�>#$����}����;K�q�Z��|�)�cO�Z������)?��=�H�Q�\�Z��R)��#{��`�܊��\
ݣ�.���ý�[o9�O�
<|�D�nU``�����cgѱo�{����F�n욉�i��z����_WNe>ф�HIz�x����a���my!42f_F�C����"�H�(��g����O�,�=	������L*Oy�-j��[1�����vUh48#�p��`����&�`LP����`_����~6 5<
��H94���ҿ��P�ǯ��L���h����ν*$���{��S"����E�&��UWJ	1S�m�V�a��͉�՚��U�*��-Ri�G�!-�&{�yt�����K�j4|���9mъ\��2��ڵT�N���=�|��Dk����)N<ޚ=�=�§.=;��گ��o�g���N�
@��B,
9�#�a�u
)�d)�w~r��t^s	����2����V�B��Dn�*ʒ�x�*�3�r�,g#SXxFe�M�[,��� I4S�{,��d}|%�g�U.����7m;�qQ����VUe�����z�aoJTǉ�SϮ����P/�*����A8Z��iZ��vj��"�D�}��8� C�v�U�o�|���2H�J�H�t��-T�2ES�.��g�cJ�J���fH]��{�[�x����>D�Cۆajl�^��-���V ���#�S2 x��ˏ7<�P�IuP"aj��L�v-� ��8� ���.�8+4?7��I����_}��˚��f���9z H��e���^����?j-ZR��'ܰK�����~�|�{J������K�iO�:Bl�F1^�Б�����b����i�� ��.}�G��b�)�@ݬʉ�L��A��v|I�ʱ�e	��E��JQn��q�p�It��e{(��0�P:<�mM��8���k�=58�R'2p�t�{��B��J?�/0Tv�R�:�����IU
�&���r݀�����T���j�0��c�\�� �����D���m�#,I�S٦����o��!�������R�ב0ͬk���~M�M.ً}��0�K��Z!kfHX�+.�p��7�}�Vn�t��b�vh�%î{P�/�t��^X>�Rw]o[��u�a�$İ��=�Y�_��W$d!v�o#���d"�1�U��?��/��\����DPq��1T5�Ux�d���6�*���{����s����)��tq=<���]��?�{�a���L|�F&��U1�]=�pu|����A+���>�tvJ�l�W����u����|�G�޵�z��&N���F�Jh�����<��z���vZ��dF��=���<T�z!W����ʵ���| (igƵۡc§�;@�2�p����<��6�N�纏#kU���L#�5��7�*�b�	��a)j����'�Lwm5�T�r�E:�7+ޤ�Q�7Pcq*j:�4s"�+"n���1�c��8�<�]�x����*�	�E�Z�d���˺��{bl-.q|Vc��҈Q�r4.�p��ɒ�bt@�=Qs�G	xk��g��L���1�Oa?�D@e0�4\�`(4�����#�F��H	����qG�\��	꽝<�4�b�OC�
��XE�Z� x�� ��UFH�2*�[[��sj_j�5��Q�_)�ƵrM�}tx���K�og�۴�����iF2�
����ĈN9�(�G���@�r6�~�)�鏟vIK��U�cM?�+7�A��\�Z�s��Џ��(�I�d��X���`�^M�Bo+h�6.�j����mU�u��5�3��Z������2���{��uj����A4p��(���Z�rdai�&�b-�6���A�?�e���ڶ�j0݃3���W��-�Ѱ՘�o��N��_����kt���F�����dM���Z�lT�z���Z{�f��J�Sn��6�]w��ĺz��,,�9t��p�οC��́\QJ$�W&���r�Ƹ
���_��H�x^�^)��!��E�S1(
;D]o�}ki�d̝�'EH���k�%�V��' u}k ��(��.�ʚz:Iz��%|�����]�,m����˥YTk���衖�K"��7$��1�"i���{��:���Q�)<P
��?Jv�9	D����Xn�K�Le�P�qADl��oo�L�Xb��'�!�M}�^�Q�X�*��
� �<Ƃ��(��6K�=����������m����0/���c/xʃ�x)r��ޡ$b|����wv69y�}���.5lW��ܻz��
¡_TM�6)k�?�������z��=�vR��s���tե �Ja��N�ԏ�&�"�/��ý�(U�<]��s N.!��@����a�U$������ܸ��S��e��_l�z^*"X��g��f%��m<�Y�����{�k[?�"�1�G���k7��vw�,i��������fO�m�ņ��ݔ�
V��%�r	s1�T�,Jk�WP�2F?����>
C����ii|������7��%>��U-��	@���~/�s�WOE#+"焋��hk��M�9NL�6�R����%-nو�e�̌MqI+�oO��݇�K��@�����ԏ	1`鬖,.O��ƏzG�1d���@�椁�3Z��[L:�.F.�`�c�<�)��Z0� V�7m�iN��>,��%$��� ���a����UfL�j=V	��|��Q�
��p���og���^ �?�s�Rb����bF{_��& Xؙ5�Tߔ���pB�����G�}(	Lǃ���r����ª1�^���"�,�c�H8�Ѩ8�lF�+�()���S��9��)X�7��,~��8��h�Hc�`�a�Q@N�M>�ȅQ��6�M���7��k��X�d	�a�YO�?kj��î�L� o��k�S?�F�O|ɲu���ղ�p(M�V��-���#)Q�P��}��M�΍h,�1,���W�Z����ٔC�@��i@JN�][nGV1~��B�ht�`�>�]f��o.������͠��+�#����4����]�\��&T^�g�o���$u���Y���c�N��m��M�0����Tq���+�'|��?��E��Y��-<� �Y7�65S1@S1r��ġ��g��H���JV8�� �s�^ZBX��^��Ң@2��o^ �r���hPLM����b%�iH�EJ�.ڲ7�k|�1Y��-�_��ѭ�}i����a&�vTKhߛJ�"j|�,�s���Ҡs��O��$=��`M"�7i����dkV�M�߻�k�X|�z�'S�w=���%p�;�xv�,P������:}��tT@)���J_F�Lt��[����͜l��q��}���9LL�Z��̧X�s�T�*�Ю^���x�n��nxeN����=�#��=�ׅd�h�I����i=k4�B���'kS��{6���� ����������^�-�Ɣb��h��˙��R[<�4Be� ��j��T����-zh��2�)M�����k�j6�.�n!sa�9�>m-(á�]�@���LYl�y���,hz�ߡ��"C��d�f��.����&C�A ��e-x�az8S�߮����|�����l��l������5�àzN8��z�X_5Ǔly�=�X���c$G�`B8v���rf�J�&��	7��)��[ڏTOzE���in�����P�H���uHـ�����ur�Jr "L��M(*�Y��QGzA�y-�����'["�ؒ���#i{�p����M2\��>�	��Z�N�ƨ�BXKғL+�Lg�褅?���$���*����� %衵��J���v; qᐾ�z�)p��"��]�z����i�Y}h$v��W]���o;|ЇE��d����o2\�r<�.�rpe9�r���"�?^ͥ���aR���9�;<gv\��u֭��H�[�lW/2m_Q��>�����l������u��V���}�t=:fN���9ki��U.���adS���d�C5�i�S��ٝf�e��_��G��W^r6X�.Xh���U�w�l��f�%�g���>���H����Ju���k
b��]/L'B��M���ゐ\Ƽ/���ev�P3�7�/��'[�6�V�"3^UE�Q��-���m�������{����gn �@H=,"a� �\*���VkBut`]��>��/�ch"?x�t�Q�V����O��Va��������w�@�ً�]#߂��{_`��`wj���a:n�����"��:?�7I��� ^F�_��/8Z�/?��H�+��<��|�%�B��q����N[�]۬?M�Gh�4���5�_A>KcO�j��D�����Ĭ���
�=��e ų�˱-x��k�G)]\�|4:u3B��v�D�S�1o�g��N���.���9�[<�}"�1\B���LD[W�>��D�e�_U���X����1���.d��ojIz~�@��.x�$0 t[�V*���\�.Ae�
�G�ػ�1�̏<2(]$�%��Y`G[�ܿϵ)T���������V�_L�)0��*���,�n�bY�&L��W�=��+�Su����^�'��\W �]��)p��=�L���4���%�[v�+�4�B��H�P��
o%�Ϙ>�Y)BB&�����do��sA`]�=�4Q���]u�V���赏��^���	��­�U0g�=�� 6QC
��U�r4Q�/�������)������ӯ�\U	[��u?޼�9��:�߭Hn��!`���`*"D���n,{�����m�Mae�x��w7ް[��U^?jOc���=}�D�'5탿R�?F����W�
�W{:��M�I����ꢍ"5h.��T(@���gz�V�CN&>�u[b�૦�<��/l���q�ѹF��I��6&+ML�&�`�f<f�yTҕ�t�h���t�$&P�ŤV;e=:��S6��uIos�(��-������Z!R7@5�+Y`����UH����7�ߛ��Z���*КK4w�ߓ��0�(���s��<p�k4v2}���`-i��}=iT��>�����/�%Y���F�=*�dUa���Q��x/�nb0k�ѥ	��c-�ۭ�^��슉��W�����8\e�9��ֽ�4h��zROh^��x�Ko���N���gBk���7��m0��<z�[rX΅z�>?\hg� �/L�`�0Y��tU�E��2�~n�����1Te�0K<g�����.g�|�s��du�`�֍�-�%��^����VS$�h�H,JT̈�jdĺJ�9�����՟��Pk�f)+�����~����"�3�I h���l@˯C�	0�$��������`��P��aU�r��W��ty��m��ی4�+� LT$����
cJ�TFO������5���K�t������t�IՀdz)dW�M�I
	qsfn�a |���õ�r?���5�i���ji��������ԍ�J��ur;�k Z���p�r�9�x���j>����';1�㖻�Ҙ�/<Ψ��ᕦ�[�4��Ol�iߐ]�Ï��5R=�����
���.u�#
�-�R�`$cg����L���"z��5<3y���T� 3��Z?��T�p�)W�]��NE�t�H�e�ϟ�E���zg~��[���s��C�~��̀]u,@2f�N��	*��TH#��=Gؐ�f���Tr�pꅯ��7�ĳog���%�	����p��5W~��!R�����ܤ�9~#ܔ��Rʐ��>i|	�M����fEV�n�"�
׫2�Fǆ�"O�	��B�V�{��2��k�`6t2s���J��E�,��Āe=�cMp�{��]��d�O�pR�n{������;Ό�l��v,��`�Y��ե+��!F.n�Xd�&�E��뭓<�Y�Z�f��v���j>|ߺ��Lui-g��|>? �x��bm퐬ns��"�R;��L�Ά�K<���y��#��tZ������Ds2th3�3�Ex\�UJ�^��!I�$!C��<;�ΪlD0QI@qsa��!�=ac/Ɏ��ή��}O��#:�Ui�5*)� #vԽ�YQ{
�ȱR+�:@sC�w����C�	�cQJt��B8
���E�� �(��!h�Ř�M�|j�H����rv�Hw�#�2� �*�\7��VMO.��0V��s�W��b���$IИ���<_�	8	�Rm�6.�[;�ַ�<�8��
BU�Ң�´&�.%�����B���O3�uAvY�K�E��u��a��i��.ې�F)6[R>���9����}$���k"��94Lܼ &�K���e���Y�#����!}`<J���\��Y����}�����[S�����h �z�摨9<�b�pJy{�����r�,i]�̯��
����iMєx�}O������s��9�T �����s��w�%�dg�Y���&_m�)ް�2���BwE�
S�k��%IA����8L]������j��X��7[H$�XU�]�Ɣ���
j섯(�J��'J�����$���*��c70�k���*bYcN	&��m���=ph�F��"�̕&��p���w�7���Ci�eG�w�?.#K���l�Y�4�ĥη,���`nQIv��F��3t]�y�h���u�ʂ=Yh�f�=�x/�J�R!Fa^2�0�C!`γ&�f'!�����(�ս1�{���WW/��Fu�0%g%�a�#�ݷ��_��{	�}x�H�8��� �CS恴Ԇ���_���%��ꌯ�oXo�yAW��^ B��%*��*T�$���%z��A����,4�hz�v�c��'��]�M�9.�L�][��ϜU|~/";�2��L�㚦F����[^p�7��J�fC?��_�0��(�S�)��Q
*d�CY>�$ݦ�4�6����B#>FE���GE����3���_��j9���6c	yWr.��;�����q�i�_�t~��$�M<\/����Z��ϟE������|�E=��f�N����o�m�~�b��8�ae�P���,��E�2�G�l�N�M�,�J=��,�݊�p����#;m�pƚ�}�nm��i;���SSD��S��-�y��~r�>?樢�Xj�I��Gf�L��E�Z�Ok���}
<�������ǁg����P��Tت�0��p��F�W2	�˰�'�ކ�ͭ؈�ݺAo{�SA���Rq���N��ͯG���9&�YK%E3��Ŋx�	H�G�%�����$@ �!���[�E�(�bTE޻������rK��º�xO�~i�7=S�P�[�n�$��7u�k����<���~Kt�.�qpF
M�̎�.y�+���3�W�v�lONms�E�(�H祁W픠MQ�G(�&�Q"-q�����l��`��ݬz�P�j9�S���z1Ţ��\�	��jQ�8��Y`�������
B�D~����%�����k�[ͼ��h�)�bT���-��jgݶϰ�Wk�v��$�<��~�Q�mcz1��jGc��ӛ*L��n����i�`�}Wĳaf�FD �~/�q7�4�	 �i�ǜ�g��o�J��B�-�zV���0:"�
g�C߹{���Nj	0:[��T���Je?{
y�xu�[��h��׳I�c?8�Q�%Q2��=�Uj\���[��ХVM)򎂫R���d�.m軵<J}"�V�7�sA��eK�R ��c�g�$����wx�@�L����<%�FdV<�1?a*� n���Y
�"���2�?+����dP�>�6=�w3�w��"���phq83,�ss/8.bf懷��tۛ���Hs���l�?��K���#�gߔ��&e78�b�O�%���!���Fڃq�!0��˚ӤtGf���K+A̭��jčW�j��k��A'2��o	�U�Y���W�Z���lo]��#әP~���-T�b �:�y�jd�]���`��zp���}���?�ټ���q�B(��1[���M�_Wi�U�a�\��384�zb	u�g���[S��`�i�CK.����ǅ��<����B�tv��ϧ/�w� �r�����%9��0Z�7�r}f�#7�qv�3R��[妐o�X�Uؿ��_���� �����2�s�����O�R̈����l/]#��M���-Ӧ�n�̶):�+t�!l����0*���jd��3�����W����C��T�{z�t}Hn����]T:�j�a�����mF(A.��o��,��ZJsY��O15"���fq�b�|1>�Ue`�Bq�/r:�2� ��D!cz:�3j���ߍ���	5�j�H�����z�h�#�I?��?Y�(� ����Ŗ0�;T�_���b�|��"3��;��Y�e3�M��m����!QyS��*F�T2�x�}\�߿��w]z���2��,S���:�n<���gZ>{>�ܻT-[�r��z�b��b��,�W�I��j�}���n�m�B�c뵪QN�qcW�NJ0ne�m�F]�*
�#o��`�?~6�����gm�MEWMF�W��"!�@Mn�7#W	Xbd@޵��L������4��JSZ�V'Usg�Z|�䦩��	��Ѻ�O@���
j�4���yR�� [e�W�V��xwEJ���	��ZZ�Pܫ���T������uB�2/X��oo�@�WWg�^= �Ul�~J����@���S(͹2jy��s|=��=nuʹ��Pe�|����+������3��p��]C���R%�b�q�:���G`�`���h��/a'��T�#�k�՛ȭ`���8��x�\̧X�������`�ɏ��B+�`bs�`��S�=gJ&\����w�[�K�\�ܧ�� ���5���3|��cr@n/佤dmX@�l@ii��eU�'YM�����BR��1�Vn�n�{�%�π��Gu�����������R���q��%�_?�<-S/+x~O�/�~?�˙؏K�F�Ā�JoB��@3�u������(��:Id��t�N7��hʶW����&���ۉ���p[f�RMU�T��ʲ��`�.�݇�å�6`�i��e9�oj�����V���E�,h+}n�q����mX�(F}*��z���O���s��)�3�lc��{�y��L�N��XQ�6�b���]���Q���PD�������}H���(�?h�{wl��.����Pd�9���l���@B��	��g���R<�0��2b�[��Y"�)�cYJ����;8�.ur$�槺F���[�1_ �i��[�����x ;Gź���7����꿧Pe��S�� l�-�#���_��uk���h����HC���W�=�T-M�p��rZ��I!ns�G��%'0�Q�B��~p�W�}�B Ef�Q�F�jL���9�QBQ/��d��dJb-!Ӷ�@$Bo]J�� g覒@�*��\h��C��b�H�߼J��q;�}I�b)n��*x�%1`|g�Yo��zZ��h�e�Mep�Y�/����$�$nm��:g��՗JMD���mS1FK�z5�n��� ��.UT0܈>�>/�A�]*�[W\C�K����_֐�۹K"����Ǆ�����k�R�y7�rKܬQ����t��Ӳ�bg�d厣<��/�p������:o0������Mg���@3r_q�F��:Ed�eƇ���"��������@��/���f���������#L��T�P����-?�V��=cl~>PH=�oi�`L
���ۣ�����7-��gB��.d{O������x3z_�F1�d	{7��P������K4��/���F5W��z��j�l�C��I�P�O�c�;���hw�#�!��k�\"���6�ν��/�Ѱ�w!����F�)}w`U�b�Ƈf�Z�#}�a���y�_*E-<
�it�@�Prk/d1�[ÔTr�'��>'�U
�`��CG�>Y�V]�z<�����%M��Z�0|<�"K�]���]�c������ջ�����i�_�A��Z��E)�v�h��6˞vX1�+t+|�j=;bf�<7�"9���(|m5|�V�BР�r%壥e�%���',-ĩ^i�Hv�%)��̉��`E�	� @��W��@��K��l�o���ðT��o�W�0T�bʧ����ś��c�ʧ,�*��;DD�s��W��1���y�A%w���2}�M�Sb��A���P���6O4N��S+TZ�:B��+ H ��^�P�[��=ZTb0����ۛ����
�6�͡UC����D�92k�J^o���KÆ��? ��1^�ҡ&g!���T�0�WoIzF���Du+�:}k��m�N�F�=�=�Jb9��Y�rm �k��!(O��(0n:�_t.���W�Ӯ+�r��ح~@��W�RuWs��1��R(Nu�TQdO�1c�4!��c�G���9�FU����=���d��Lq�F���8^���h؏���=�TyN���/+���蒠���B
�� hlzod}�-���il�n���P}A���u<����6�� ( �2<�`��˺!���I��m׷�*fSX�l����`"c����F7�N	@�W�8��xק)�167����,��m|��ѐ�	�&(4EC�N���G��ugb�^���m)����jt�����o+"|'�[�8�#3�+.��88��x��
pK��_XP
<W��f��>v;D�76d�<��{�o�o�v����W�?�[���:����+舖�2���ލzs�/'�ԹN��D<ݰ�B�����ys�p��t3��u�$-�&��%]�ʐ��ɳ��Ps����90��6�x؝��g��K�(�rZ]y�oi�K�t8xi��,�͛k��k?��$��x���Y|���ߵZD�@W	��v�Vէ�A{[�
����5A���RZ�cX����B�)�w�Z���/N�������ϭJJ��c���&�9��zh��<%��Q-y��__S�Q���S�Hm�*uy�%_���iF�'���@]1Vå�jQV����5�W�@\a�dR�ڔ�0:[cfhTfk�$�s�;�"i9����J��)��J,$�,�E�R��*\z��(B)�<��r�B8��	�2�����Sk��YH;���i�<VӉ���s�ژ���U㘡���ɛ�U$�V0�`;��	��,����~�b�W�j|Os�GE��05�A^��i�o�#�Q�.�75f��׊��`AŠ���k��&O��4��|�O{CnK���,�|�k�MBW{������n-�R�m�,�<a?��k��Ӿa�!=	v�=�:����y�*�P>�����ج\��h��h�a�&���_�π+����D�^Ԑ��I��ɷ�vR��36��4�7�)��	q�o@켤������T@l�_�XK~n�wB*��-�����F��_��q�U3����M^���m�;�[�b�7z�����	����qK�*�=Χ��]A��c<��đ�U���Ct+�m�*�~�ݸ|-!L)&�}7�8F�$�.�N�[r��T�Ӎe�膞à��8ys
�S��]��1v�͔薂��A�u5k��B���6S�9�.���<��akLb���v ��=��%��'(Tr/F�d����%�۸�йV�9�Q���x[E}��|��H�\�x�"��0�M�;WOwt��<U�9�8-�A*�,0�.�R��۲��В�=ԟ��B���A� �P&���ѐ�y�"~��@--Q�7�Dc�q�c��ޫw���������\`~p����&Y}8b����(���Q���ك��[~����da(`[#W��c���|�2����U�?j\��θ��c�*�ҙ�ʥ[��,�~S��&Xur�����/����m"�ؚ/t�������}Q�b�9&2���T�E��< ;7xb��hI�{�S{GB������$��/��:�\�(S��!�Z!�����N3��-���Ι��:d�.��avz	��>��Ъw��[������y�'�w�aܴ<�-�?�J�~?���{ݷ�6UJ�����a���E�Ze'�[��8��n�������T)y���؄W4�_�|��X[�5�LC]�	�n�;��^�6I\da��J�u .3��k;D<�ی&�2;���Ξ�FlR�lUF�ll��
QmtA)IG��d"%Kž0lޘ�yP�_�������P�,2��!��z>� ��E�e���?�䧁�p�s/e�
��)\���\Ǭ�pE�>#�a�()i��
]�Q����zc��aCS��d�!�/����X����.��_�`��N#I(W&��C���'���
�iF��c0\�>$�w�����E�	z���-��s�����M�����4����>����:�S��'#�O ���@\xc),Zg��N��)ڧY���.y Q?�s������
<D�)g|����겪� E��.�E�+'��bGa>G[�!|�̨3�m���κ	�oca�CoBn�G��:�b$40��(b���nA�Sr��p���eN"
�.i����'E���qtOX,{iq�+O�:�n�:�r���j��:l<�Gu>�K���=T.	+���kߝY��"�@ϟ{j��,�>���EG�9�~�4Qi���q�x�u�Z��d(#�V �p;�V�8������O�1m\.�ef w�n|�c<󋬴?Q��S;��P������W���PV�(�n�|���B���^/6����h���K%TKY�M1z�sק��?�G�5�+d��0N`�Ӻ��S��:�4{��(����3��|���[Q��������!���GKƚדѭg�<X�c��\o<)��ʏ���d���Qg��Ls	�Ƶ�Dw�Wn�á:Sm�R�ν9� M�aU���$O�XU�p��XQ^T\����ѧO���s+�bM)�`�P,���>�?���E�k���a�m�n
�o)��xP����
Lv2�ŕ�=}C�"�:O��G��5a��,��Z���,(g��v��N��AN�߄6P>Lm��u�T��s��P|��	�(���<��(|�D�iT��9�̀5�[���W���#ń��S���V5�J>fj�^�"�F��~�&q��]BL��8�؟=������^�2���Ww�T�`��wo��CC�9s�O��aw،u�G��U�.��X�

�j���D0��� �q���C��B����B�U�ѓ�d^�B<Wb6��Ab��C[k��Y����i�F��+��b�E��Tn���I�gb
 V�胼QڬQㅿ�߲h-�����z��V�D΍�ս���;��*EP!�-�4y� �D%�C;�
]d��yov:x<J�ݯ3�J���+�R�:}\��x"�$�9�$E�����潧N+e���qJ�qz\v��)q�b9]w|C����҄!�d���@�j��YS��	hC�v����zo�ޖ!�a�;����>��<���%D���֍e�;l(�����#@8���T�Ê��3#�ߍ�	���OԻ�ia���Y}�g��Tj'���`ax�4{�~�K�q�4�2�Gm�����B���Η���`���o�O������&�j�`�ܱ<5��Ԫ��4�~w�Q����f��h�B����Q�[t��4&��Y0��/�0<i�9�~A�:QL�/N ���h�bB4g�\_��#[�����/s4�g�����i�,��&6C.pte]`B��T�i�8E�2K�l������?��=�e`B�e�?��Q����(��y�s<��El��HuЗS��rG�S���n�k�p��Z5��a���Te�	�3�f6���o�Q�fEh C�A �M��HAOPm�?�$s��Ҋ��w���:��LA;���Y�`��JhP���Q�,��z���tWW��{�%��+	y�T~5 5�9�ND�b����h5̄�1�V6VoȌ���6V��vD�mL쎥x�#�c^�ci�>�0t�N�Sn��)����u����K|E7TK�)��F>�t�H�~�L��C��g�WLx�xM;�l�ZԴ�6�T88Is��'<b!E3WE�̌���mNk�\_� ,����iBb/����j{��6E���vf/!�7"�<���\?Q�`���������ˬ��#H����=8���4j��k��(q L۔M��<�$w[
Hvw���'��3�m��U-Pq���s��nf��NVW�^� ��!`9i}����8I^"eE�?v�4��a�N?�f����������U�}�'܉�b��1쟎���y�{5L|�z9�p��/x��d"���v��.����R,����n���4BB���qP���r�lL�A�� n�c��[Z�)��B��B�>��"����u	􊛏S��|Ѐd�%�:���Lj꤆�(��u�W�q�Ti��l<��܀R�nˣ��`��@�)�κ8���r8�6uUj�g�&VI��
ׂ���& �Q�c���,%�4�J|ߒ�3fa
'�ܫ#Qg�TS�H5?g<�D�����M%����y��>�!Б4����G5��Q�˻��&XlԄ�;�$(������5z�� ��Ͱ�Š��ǡvP�4��<\}.�,���{,�����?�F��ܻ�%~�"�~������vm^9 �w����M����;�E���	c� �Mh���T�t��|j+��`�)�B^�B��!c,���-ݚ�o���XU��d��bA�"��E�l�wT�)�3�EW����;S���CZ&�鳙#�V��PX�4}7x�<��5����h�/����wi�'���24u����
�����7��~�d��$
�8����W�����J�̫g����O�aV�D�S'���Hq��E,ق��|G��[{��/*��/�P\����J�����/ա� �x��)�e�lK}���'��DUt.#S�A���{����Y�����F_0i��h!W$N����*���"9P5嗦�����`%�g����+�i���l.I|�{��%q�V��y�zx�f&�����Ā�W�?�kI�8)�3O�w�+	���)ռՊ�o`�KK�6���v�vC=�M�>�Zí�ஶ�<����ԼW��H�˳�]=�Ic��gH�g���hb
n����D�}˙f-��;q������[K7*�7$>:�pb�;^l��f����W#���(�.2��-��,l�<��"��Ol^��g�B{㪖��n��:ŧ�r��Fȯ����-D�imLJ�"'~Y:O$��L��:�9LfA��#l�xk]!�/<,Nz7LC�ಢ�!�S����/n�`��á���I��.cV�� 0ɯ5� 4?�O����U��J�V}�\�ds��Δu	��o/S�#��kz\2z3 �zNA�S
�re��m�,UdI��PTb��$n���oW�r�����u3>�(�?�fͼ�S�H�V�l ���\]�\����-�V��#.�T��J�=h�=;^$��Y�v��O�[����52��ƻ?��~�&�D��s�6��4�V�AV�IE	�
�Ws����:3�����jrI$��`k��ٮw�����@�y�p���R"�?��aJE�������^��Pm���W�Icϕ���"���Yg�k3�T�Zy}(}��܋>�"@Ǫsn�ͥ����	��#��˥����r#�I#�n)������jx��%������Ǒ��S{��(��_��&GM�:�<��aGse�jc5ݪd91�j#y��.CJ&R�����Q��s��O9P�C�P[ݒo�KZ%	��َ+�)b1������8cAa���8�rF�W�{�he��َh_�� ���s�M��؃c���)aļ�j��T�NCi�w	�3��̳�邡�y���l�9!��S��`�DN��8��(<���h�jh ������k~��)1�)^}ݑ���S���J���� �^Dw�(�E?�(v�]����ZH"�Y��㎀��g�(�7��̇Ә��#Me]ʆ� @��ŷۛ�^a]̌2&2����E柜#b��ۃ�ؒ:��ن���3>2���m�FӔ�X��[��z�lO�g$�*�o�Z"bŔ�5�hnt���F��<�F��1R�����y�;�hxm��9H�{R�>����%��dQ����k���w��2-({<[$�l��*=qK����Z�9��o���.15-%?Q�`��1ku~�c��ӑt�zZo}��}6���.p!�7x��Q@��6�MM✈�4esvBJ; &�n�H��ږ�X<(�����bqB�S�Px�p��u#�h��ŬAJ�I� ���K��U��P�=u.��w�h�S_���)�x������l8h��+q��J��K��6�ɭ�������L��<?Ͳ_����3�5&��,�^v\�S�%���m4��˕��d��;��|��E�n��7;9y�l���*2h�I䄭?�&�o��͇5��ϛ�~�0q�������(��5hA�-!��+ބ��e�I��6g9	��H3����u�b��m쳅��AǷ�`[�"q�9��ވ��Xto!h��<u��X(��<��M����!Ec�"�Ivp�}���=���}�Y�[�!��Gr�NM��_5L=�J�_|Z��6����+���]t|1S`\�-�~LU�ߗ�'�@��������b6[��zULq�F5a����rv8۷�o�t�kn0�[�]E�ƚ��8.{D���������`<�!Z}j��_a��@��Y^�${g�;E�ϋ�ޚ���?\u��cқ3(p�\�'(O��c�k.U(řczetS/w��ʹ��V*�i���F�
�I�pUY�VZ�{{���:��å�k?12N։0�4����뙿�;Y�RG��G�[�\�r�1˟w���^0	��x.U�P�f�}L�6k�_֋p����j+kO~M��^��:g*c�~:���kU��c��	�D��$vm���\x�ޤ`�P�˔n��WBG���)��9��%uWÎ���
+�y6����l�]��5�]ef��ok�Szf�S&�W��&�)�_����c��?�C�� ����pL=���ݏ�Eߕ���Ŏ �2�;*�����<��o�k�O·*�U,���0�>�F�/f!~:�/�\2��8�LOi�c����N�_�ْ��	M@�E/�HJ{o�D����V&ˑ�6F/B�밋Il��{R��D2����Ԅ\�R��C�O\��������0�jkC�������+�=,�	*@&T�%�;z��$�&c�T0�}k �����Lt�甆�U��|�""Vq��ۛ�"��¡Q�x`B��8��E��P���Oi�Qd��",�،ӗ5b���}v�ʹ�-٣ X/l 0�ۿ����<օ�ȼn�4�Q#NB��G(����ޑ��O*q��ZO%�m����|,~�+��c@�ޜ?M٬g5g�z��O��>�\H���g��{���v����oP����Q�}bi��|9,}���)�M�dx�e(�>+u |�̛���ʲ�����2Y4?Y�P�=�]�T �Y��I�X�3L�}�#�%��`��~YɧP��iv�Ӭ\��H�λ�"�I��U�M,>�S�=���TRb׫��4�UN*w�$���Nt6��T��J�䚜U7����67����1��6 cN�^�bu\u���KJ��C:��0 �?6�i�{�T���RûI/Ԃ������j�Ɏ��p�d�N�����t`��w<�������/B��c�?
�IEޏL�{���%��n�ۤ�ó{ٝƹ�u��_�Lگ%w+$��Х3c�=�i٠*K��_ �ItUQ�a�9��؞��H�R?�[�5���>�k��|�߳�
�H��c�r�-��i�߆IzD����<!׫p�B.�M=(�O�	�L`��������x�13:u �Mo��c���鮯�V����M���9�2A+�R�����F�5�����_�}�4��5l���ߝ���dZ:<��7�]>�0��ß���g�_�zx���>��G(�T�ȕ�ɞ��g��L+\�@��~�uM9V@���@GG��Vt��D�6i�ghOK�l��5p�M��w=驢���T�ٿ�Gb��DEM�.�Һϊ�v�M0O��͙[l1���0	�P�9��4*6"u��\�h���~"�Gړm��<��&�����Q֔�Rj[ZG����:��'��yz�v���ȁE���1�����>���1;&�kH��O���O���{�p3?�e��U�����`�/��aa��B֖=�J���I���,o#��h�'_2B*2��I�g�0�����2Z�'co/�q+���?�B5�2iJ�ɩ��V�?��o��N�h_$T��m����O2%�?`�s,�~R4�Ǿ�HR��14�]�ϼTۖ��܀ݧ]���In��O�:�yR���&l���;k��*�%ϥuz�� Xj�u�x����G�?�Ƿ�6�˖�i��h���Ӗ�H�bt�Tt���� pI��d�+&(ޓ���_;��38[�"A��$\���D�PkmG�5U�zRRus�:O\ǥ�#��~E�����*g2��˅ 4��Z�t&my�ޓ�6$�y��������%�6P?W�z��lT!�=������O��9� ;LX!��.�^�	��G�R��&|��~�ݟ	*�X�"ɲ��al��Aì�ݟ��h����9g�ٞ)_����{�a��ދ����if�>H��շVŐj��%����.��)���%�N�����0�_�h�#�&U4Ӿk��[=�>��0�ibG�ɰ�F�p�P�,�e�����)<L���
�d"�Opj"�u�I��	����O\����e�Bv ��o(V�-�
Vr��-�i#�G�lJ�P�.)բ}�5�nF319n��<yB��g���z�s2��s�A���֐&�k��R��"΁�h� G�����nn3���
1A
J7��;Ւ�-Ҙqo|��D����[c��	��=������*�B�6
n%�(V����F���x�륵O)�v���↛�����cn�K��c*��$�=�VQݘgH�/����؇43���EP.�8ǈecg��K�bP�
��l/�2��O�I�5�
N3�{��!)
��5L=�hbS�Ol3��W�P� �dY����ٵ@Nm�IE��˪e��@�n�а3�H������j��x}�p�E~)����p(T޿6��'�F��'���~���n
�1_�������əCv7a\���-�H�]�
�2G<
1P׊oR�c������(�{�<�SSY1���-�"��)[,�?���ls����ʈ���UEY�ӥf[ ־㿵ҷ�#�+[o��ț��G| �/�_n��/��Zk��c�U&�����������(��+���f��R�=t��4�H''Θ�
9� ���5��:]j��9=��6̵XR��������چ�;H�d� �t��A��"�����X~Gh=@�����?�}W�pB��`�b]�S
����s8��i�*'�;�qD�c��1	�ok��UAձ]e�m �����*�/� ^��	��&�
K�CF��X�)m��P�:�Gmv�`1��J�KN�UPY�R�H50�u��ָ�/�m@�K"N,xDx"�7l�i��RBr��^(D{���{9=��k!)O��X�NOj�͝��v�˸]�Wߙ����뇹�����[�g���T�`sr�b�7�P�F>)ŏ�T�ZQ��
H�0en}� ��!V�|����t����?ݴ��-�:���-�$��</VTO��"I4ˆ˂�jǿ$rSȶ�d�e/V)Z���e�^�f�1:���u����şE�DY�F�?,*���7�E��!�3�8'�?�U9+��P+C�1�5���ZB�3���Ćj��ID�I��,?S��|����ڱ#6��rZI'F$���V��*r��<_�a����οlRā��˄v9��^)���,��w\��I�.I��=j3cyx�žۿ������[]�s��hEJ�'�@k!��a�>�+�=��lk�6�Y�)�ʋ���M�ץI~��)7�?}WyOBeQPU���(�e��O�7}e"�H��Zy`a�95*�.��>!��ץ�l�����)�*4�� V����<�v]�l���KN��G��O�n�$}ū���g^n���@ӣݍ�b��ǅ]ȐD�_e>M5��X���W{6:+�\���`��<F�p٠w8��췚�Q�IU��!�`��^�<�u����j,�/5O���
we~g��\"��­~d)��b��S>ڐ�;���p!Zd��s��A],.j��e� -�X1��
=˖�6׹s2�Y��@��FU�˜������c�>�:i�/9����c\�sȂ��B]E���.�\��b���.�t��%j�+u�&j�������3��:����^��ח�g�#:m/����^.��D���ձ�ӊ�^�#�?��!r1X��mA&��8N@�#GM(S�?�A�Ix�~M��:�q�[O8Mc�p��~�jȁZ_ͳ� ��< �Х���r�y��5�*AC��)����0i)A�'o�8
�"�
��:��wL�N"{K:�:w
tܧ�:��$�G�x��3��;?����1i�����Fb0�zF��8��C,� ��wZ(�9�	�
b�"���G@��;�0���A���E�)�M~�v�@#ć ���:\�-� �S���z�
��45�Ȕ1XI����!����ɐ�1v�A�Gwg@���!S4��HE��|��ң����B^:�����e�F�hH�����"tI�Q�ǅ� ��G�Fu��[Y�z���8��g��G�l������A���3Y㟎��-h(4nۢ��-"���3���k�O�񜇞U�yړ��|Lgej��c�,����W�<�q"���)r�L� 2g���2�w`Ǽ�W�O�����Y�Y�{�RVMמ���[4�I����τ�v����p�{P��ӫ����,f`ّ���Ev���S��c�.*漤zլ�� ���N��0�aœ}H� ?����Ǧ(0���@&[��cĄ����6q��\ &ʗ�m�)��R�[�yW�p�5�?���\�cG�&O���������k�򁷅P�Y�}M�J�v�Ȗc�]��Rx&���	����b�@x_�||r��є�_r;l@��\��+�a_8=g��K��\u�����Fp*�j�첕�v��t|3<0��!S*�R�˞�x*�S�Od ��q�Cb�QV.����~U��%�����>'kl��}�)IZr/�PTK��Mxayo\&Z�r��;��Pi�;#:y	��<O�r�u4Pc���ș)�F�	z��w�X�qzBC	Z��3-�jމv�Q;g���}|�ƺ`۝ݻ��F���x=�O��OG��?���s^�R���ʁ&��<�. �!���
�G0`m� )%�lc{C���$TM�9�}y�<Jc�JI�����9 <*�i�Y�_'
�m�1�'K��������#���oȦ�����v��ܰDѩ���&���:	2�ek�4qf�C�Io�t�k����^�PK�em��4%��*Y��o�C�N-���{�����#m�ffW�9V8z6	/R�hJ�RO�t�А�2�����2)>{����~��xB�4`�
�I�K���3<E����*Hyo����5���9X�n���ul|-�B����Xo47m=�i��	9���G� Q?�Y��r*�S�[O���J��Q�����{�Hn���@oL��ߧz+��
�?M�;nuj�	`_(�S�, q�!y�6D%1O�}%#Xѣ�oE&�n����L��@�y�p����#
=�IK��-2mH���h<�m��y�B?�e�$��y�
�Sk$�|D�ƫO���\�Uٕ��tj����_Ͼ7��m�E�3��5����[eك���6M!��;�Z9�α��#\�
9�� �h��ܽԓ댪>ɔE��ipsE���2>w7��)F��Hi����Ja�J��PS��T���K��t�D��I`I�ғ^j%&}R;�[{�V!��3:����f@ᇉS�a����Ҝ��Y� /F�\�~�Őq`��"�h0� �1�FΩW���w�MJ,?~�������"�V�(��,Oۡ�	��$�<BL�.���V�+��_�~��l0&�Cy��7Ht$��_��E/�-P2�_�̷(nǱ�� ZS��Aց�Wo��vڱI,�L�Gt��f�<aP������!��װ�&��	Z�<�
U;��su��B�R��C�y)m$�9�>�ۄ�0�Ģ#��G��/�� �~
j�0�Ydd�F!=5>Y�K�l���O� ��V�Q��g"��&FD��d�P� 9�w����81��f�;rn����W�c����;&�՞2��N��B�i��-l��h<'8a��1s����9�]����Xy��'�{33U�V��n�dj��l��hg���;�;Y�A�:��\���y���fGwRd`�Ej���ב�K��YC��3���kU�<IRxG��3���B��ؖ���1��.�rrN|%��υ�2*��V��+�K/~ƖΈ7qBWc6��'����Cw'����(�?w|�o�+^�?v�Z��6�KN���-�=��B�����S�K�m�l�&<�P4���q*p��	�h�F8Wٓ���G �����r�H��cD����1u��H�&(��]
na�������m�1�)�=�����bO��� �}�G�;YZ$|�x � �S ��b�`OD:��{J!��҂�㭙��*	8��~:�J8�2%�J�V@��sˎ�U/�	5�-�cSا9�WEFpDN6Sl���Y����=]b��q�G�x�M%-�k� G�1�՛���G���hp}p}C��� ��!k-��S�d�	V �L%|*����*O��0��wC��G��3m�Y��Pjs�O����@�+f�/�m7�6�)�9}*1��;ׁ������J���?T��o�M�<�.��&���-=�Z�e����9r�����-�*G`���$BT�&�$��<�eseC��u[���4Jv�]|��K�	�j��+��;���r��uO*`bn<�w�D_8\5!�]^�r1�J�k��c��C�m�)�>}�~
#�\�G���}@�C�����^c!R&&����F�a�2�PY�<j�
*g)��+�RRYte�hG��wʴ%O�>
�G_����4H�iM�o[�����g�A��q��L��eID��~���Y1�$q�||F]P�	���m9�K��m��s�
^��Jg���h���9"J��M0�pzi0�;��������m�T�`�oN��b���zF���5j�\cy�����]��6��cx^sW�Ey.XU\3;B!��J�o5�mO�/g������\Gj��J1�?�hk���|�}�;�J�7-d�����<�E�8����y����R��FgE��=�d�~��U��$�����T�ܷ���Ō�g����g�v4Q�|���0�J���d�WT~|�[�[�N��Տ�*���e�.�%�/D��?F��nPN��ԠK�6���l<gwhP���a�w�&�K"&%$��Xj�\�yR�q��'���V�̑rX��X�������O^�W]7	�×.��a8��(�ݥ\<��s=�P����MP�*~~���u�C&�� ��뽇���V���Y�\]���d�z�h14�ǵ(|F��,2��	n-R�[v`�7秪�m�����F��< b,؜/e0v{�5)�A�jTe�y���x����q�6�R��nӺb
�gX��M�!��<
�.!)PL�Ƣ�r}j2�eC�<(_���&�V�����P��Ńo3E����1Z���*��M���G��o:2�٫b�*�������z?ц��]17>�(C�i�.���A�ue&��sz�5�R~���T{{k6�;��<�sO�p�%�����J#�?RD���cm}r�R�l�(��l}���1s�o�T��L���M���)쩪�wcd3s��:��K ����VJ>]q��𚒈��n���ҼX�S��U��)\^S��[��JO��*�|��������O#۝��p?�y�zc�I��u�ԛq\����r_�b��0f��ѷ�ݲϴ|K���-�aX<�v���9�]��Q$X�R�ae�B�c�Z0q�8f�p���-���n�}�����I`>O��C2/̓��wW>�̈́��
�EJF���%������Ω%��U�q�f�[�?�;�	�WEc�.�x*H�xn�W�WgG����.Ѥ�3�wh��fѡ�4Z�F/0n�ZB�������v�R������F�N^���ϟ���3�����v��n���e>�#���q��9J��o��'5/k�V���J
e�*���⧂bN�ך'�>�Is�%A�`�(F,LA���}V�R��\�:��CkX�uץ���D'wy�����JS�z��*����M�g�j��� sg(i�O�{��aC��2H�}BCJg�b��$ڗf������~��=N��fOkQ�����[�^¹�sžH'�#P1m��29QV�Η[���t2��>�g�g�b�À�:NeX����]��s3�׿��w� �[a��N}���b.J0�X�._Z���;���\loY�m�9t8�<�zy�l��MҲ�D�R?������*a����?�@�ޤ����ᮃ�%�<F\��8Q�S˕���K��}��1�h:����`il�\ᕵ�1G�za`���HL�P�!�]�֝��ݟ���X�1�v��oeK\k�e��
��;8�'�&���ǂ�){�f�R�\�1یQ���ŉ�M8��X�v�X��%ЍO���0\ӿ�׹���k؊�<v�0@7M��L��S��X�A����W"��Z�&yp��Φ)F�e�j�`PQ.���p>HN\�P�><��2ض`��N2܁`@��C	��V��Ed~�Z-��В*���W�{�=yn���%��eE=��� }�=��7qb�1�W� Lu1���b�c�%(�n���v��}�NJXu_-6��zM���X���������E�f�H��ҫ���r �8��!���MƋ��W�W[��a��a-�TL�����yO7���<�MRI7� >�tp�&4�&�_l]|�胪u��#F%Hz�hj.�Ӥ�+�z��1�_���G�
 �g�S��LL�/�%{[LHw��
&�r��R2�6)��#�R��حS����;i���-��@B��qs
��;H��y�K]��N׋m3Fӎun`2usF=�/��ɕX����O��������[��
����;��ָn��J�ܟ���69uyk6�mzm���v-C�x�q��U��9�W�/+��}L���F!tlG�"(
3�T[uQƳ����U�#=-�(�6���;v@�ß��6��3����qJz����y�b�'�͋E�M!i��2}�Z����ЬC�hl�`p�G��^�R�����(����O�ԱR�y�����he�y�|f�WՕ��O�U!�̗�rPzN��a4t�]z������`��3i�kL�Rȯ@>8eT�Z9�#��bě����  5%�����Ӳ��!�����7/��9(�Gܺ�-w��u���̊��x�����UHbdퟸ���G>5}�,��y<�a��z�`h��<�6��������d1�:�f_���x��w�Ŝ���Q�������t�e�h▽���>ѷ#�>衙�LK-ms�ݛ��8t���+�`�h�ԡ%^�.x4z+'}�[��7���L�8h��QI�����W�[���݃��y�R<��u/F��eM����À������k/�RLbHGLY�
�}`ȣ�&��+��D��k��K�i�;��$�/GH�`q:V�e�X61bu��Ā�z�ap�y�t?�!l�ޣ��j�'������ՠ>�w��r|@�aO<�e�l���t���O�W�T�$�A�
!B�\��,�6��ou��cj�&Z/W�q�Hu�m��;��%��=䪇r�% :L~���ڒ?�Y�W�:p�6�b��WZ�_K{��r��D�HG=oZ-r��!���m����4�.}��󍧺�pm��w���K�D�i�c�'�>���r(���Jc��,[������wb��,���O�S~y�L;�ͅ��J_<�B{X��G����3�Dj^$��J�����;�2�v�&A�%�s���YV�?�u�i3����#���F~��%) �D�@'�Щ�E¤��E7+?ʅ���~�����8~�$sb��x��Ԅ�B�EAi�%2�&xJr���Nq����<׉��T2ݘ����&b�����������C8�Y�B�p��"Y�����yѵT	�
k
�s��`����	 oh,���/����4xP�������[�������6tW�I�UwL�	Ƭ�����`���ȅ��^�cT����;��AOR
Њ���H44��Ek~�9Z.�x1b����5�P������0jS���UO^��#�r/��)S�tD�8�������.��|����c�����g������ }��i���Э#$v0����L� 8  ń�nM!�>3o��W%�?����PkpRp��$a8Jc?D�ւ!^H�3�o�v��<�&����a���j;="^����ȗ|{�zu�Ê.ֳ*��;G�{��(ۗ��/��5��8�S���1�8pk�U��c;�_2�p��
���.d"+�? -�ee����gFxŵ^�����+u��x~����[��a���s͘�>�vM��@˕q�1�+�A�Fc��;��Ò����t���e�7P����A@�G�om�{J�Ȩ�!����=�^�����h�[�VI+�1K@����t�����:X<��Է�zd�٬��k�W� ���v��!��q\�{��fLa` �����w�����p�!+yZ��5��We}0/-/��g{��Apzxw�,U�{i���#��64���s��J��Z�x��S��M&VU����1���U�:!?� �[}��;�x����a�C��
Z)����u����#�E�Xu���1���YL��Nݯ�*K� c�L+����;�"�[TE�<�fZ �}R�Qj���MB��- d�λ�� ��DQx�"�%�$�G_3L�J������C,"g����5������3^���VFs���O�F��v��ÿ@���-���p�~�.����[�Vf!��C��������#X�@�6O[k4*믎nD���Mz�\�����	��.Ũö�A5�TB��O�ZC�oH�{���ZC��,������u�����j�:|��=E��Nҗ���.)����4��ɮ*3�a�̘�-�r]I���1'�Y�ԞNw�yل��E�z;���(��?%|0���d��4-nNH����H�ƍx�"�͵��#=>M�q��幉�݉�e�nlZ�P��pf��`mhy�r�o��㖚�ɹ�׉�Ca{wUxlE'%MݕhbM�qD8�Y_�gI痌��&��S�>��]FK#�_���h�_�CB�Ϳs�OR)��do[�Õ����o�ޛۙ@��'�m�kM�D�Ý
�C<�L�0�pW�+2�?��+��➓�1��a�k*����˩j9t9ơhH��H�V]ה��y����:={R����F܍��_s�O�.W�}I��]��a�E�[U�{�3˿ta�?iO�U�����(<bÃ�܀����j�������ν9���s%�M�5��I]A=.����皳��z�lF��X�D�O(ŞN$;fy*���Sk.��1E����^�ה�(��n2���$-�Nn���V�ե�0z2Cfo�'~��O��}�����v1����ht��Lz�x{r*�M��IG�Pr���~��h��]����c��� �J�(;j�)Q��y��a���*M.���J@ �0SA���5w���zA7��ȴV9��S67�غz��u���D�ŽV�k
����`�J�l�#Jh�gĴ��>�Y߂q;�����l፿��y�k�@�_8�J�eg�DLF}���@;�HZ����'�+�ͳ��s���\=���'�ɽ�$$�:K��GMGv$��s\K�q�sd9!�������s�o��C���?�FVi0#l�_&gB0����A�7�r/�)#�`%ږ L�c��Kϲ�ǯP+��9sG�cZH9R�q+��Q]��ft�)lV�;��~�~	�݇s�M�ٰi��N�_a���o��~mԦ�K�����/#
�r��YF[&O��V22v2�V���rIK���$�Cm��i(7r���nd��ȃ��l�3�]���=D��%�#�3b3OE���$���n~@�	{�:Կj,z�#!s��`t�N�آ�m��K^�i`:�J,qbu3��|n� vF�;�I$;Q�1���#�D��3�v	�4'��Oos���{��+��56�-�ܦ�5�)z�HL���f��
G�����Nr|���d���yR5��+k�T���8 ٧|$��J���G���@�S��e�<�	��JLq�T��8+�f���*������@���o}���H��ufBΚ�u�|��Û#�Ih�$^��}��N��<V�H�#���;�m@�~
�xk���D��S�g{�
r��SHÕa蔅"4�K[%�
�BI���H�O�����#a ��������<���R�D�}��
@�Q�_�x���6�Js|�j+hJ�ɼ)Z�4�K{��&�^�G��Ltu>1?Ģ�� �����L>���J��x#&��S�Z�AGx�կm��Ss|HdOB]tV+S�U�v�30~o\���\�#(z5��Z�l���\�z�t1���Z̻=��;�{(���0Q����F��>�.�� h=���|�[�^��v�������*j+�q||��B�qV�1W�򞹺�DtsZ~N��j8���bU�'�V*���q��0g��uG��q(|���Z�*lr����G���ܧ��[D�i�!\U�C�sx�Rh�Mf_����#h/it� ���,�]ቾ=KG�Rs\����Z���!1c;��{#�E_ȁ���$��>#���R7 ����X7'�~y-���a"�o7�_p>*�[�7�"r��"�TԜ�5=���S��#���v#!�� 4hg�X�� ��6��T�����6�^��j����2�R���k^Ucv�DCe�2--��N̉��s��u��Ə힞��Q��w�y�Q�ٛ�'�/ܱc��|���؂	ȴ��p�!_lA����4��ۛ���D�&�@w{� �߁S���t�z�|�-�K!eV��+��
RI�D��0�ş�}|��T�yG�-��_[�����`��T��������{�m�f���w2t��������z����,�	L� �|�Q�,�H�Ŵ=!%B�@b\�@�Tn�2C�}���C��ܼH/�U`=*�|��ԮJp��Pݴ%h�v����J`� ��ުeR.�q�cQ;7%��e\������y�o���|�X�1�!�$���V0�����@P�h?��?^l��V̓nE���h��O�+�v��_��)<��.�qI���{dTp?��-�>���s����1�S/F�b��i�
���)�Ajn�D�`Lӿ��J�M���?1�V�RfhN���yC�?������'���ɞ����-�<����ѿ'c�?��,��00��PP��2u�sŮ����uN�����Toţ&��tDC�=�Z;�.q��]�#�7mf��.��H����z�i�`�sW�_[ǉ9���X6��¹~.��r74�Դ���W]8_%�6=	؅���>S}y~�-By�˕���\��X�|�{�/?{"�������cQ��n0�X�G9�(_�n����� r֎�#���Ti�z~|����`^��VTo��nCd�����-/{��#�7D�u�u�j`��w<�<F0�PtϲL^�(����d�w��:����7��:�}��7��W��\*c���<e&�i�ws���y\d7u\��7I�[�7����{1�T��%�u��s8������=OO��!�H����}J򼊌4��mA����-�8�fJ�!�S�xT��6��⇜�u�[���65�a����Y�H�"�±W۠~i�S�P���|'����7�̜�0X�-�>�ሢ�ےçb}f�;1�Ƚ@Q	�өTmا��I�75v���q�
�ۍ�$^�W�q�F���N�� _���iU�ZB
�>t��&m&�T��'(h�{nt��@��>�r��b��#�̖ r B���E*r}gu_2mN}�l�$��&O;�i�2��?x>uod��O�%#g!�4�2�6�;g~�l�X�4$�Ϡ6�]0�-��b��W�\���S�:���65�zcu��I�E�c�U=v)���x��R%��쾜��z&�"�(�褞v��S
�!%��,��|��eW���A���!�Z�j�a�a�B��y�^��Z�i?R� f��*�#�m%�q�[(����e0��sS�_ZNi��u�+z.
�/;�7�2�%V��pD>������pY^��C����7��M�0��'�y�ю�*DB�x*��إw�#��(c)�gͅz�9�+���Ax�J1V�3kcЮ���G��E�!9�-~P�^��ҍ6�E�[={79�\��?a�Jw�m_��^�GѩW��"_n��G8_�w�y"�������8�#&�,�
q�3�����[*{��YB|Ŝ�Hfj���`�Ũ b���B8�"�%�D���N�B7��s'q�8�Bw���֧-w�̜��=_�u25y���v��}�R;�:=A�͗�[��Jj�ԞW���D���+P�t�پ���n����X�JIM|�����*�l<�V��q��17|�%���ˆVt���bCh�����&B�h&�Ћz�qv������� 0���vA�}1sU�7���9O���m��g�0�
��2�	\~O9u���2��5PsT��Χ�$&O�"p�3��m3ݿQ�]�-~5�Z4ڑ�;���9��X��?�W�O}���
N̙4g�U3����:D�┏�u��QY���W�f�H,�R��o��Z�� ��Aj�J��\<c��3�v\ɧlູ�Q�\�)C�<%f
ל,��Q��F�h�r�I<S�t�kG�cN��<�,�W2�J��y[�����w�ZR�BB�j�)ڱ�5���L�D�d�cY��#6_�j�IH.�8�Gf=� ΐ��?�ѣT3����;�"m	�ɬ�h�⏏+���5v�߹y:����o�~�@w��hQ$_s3�e\S�rk��v������$��
܄#Ld�d�O+���t�� ��(��;��=�0�k�+wCYg�M�t��:���l*`���("4+��������D��1&���X_� �c����p7�ڠ��0��2��.�*U�a���ĪTl��0�����D�3�~��~z!�rk��y�*��)��O�9��)�`��6�0I��T�4�����y�]�0�{�T�9cc�6��`�-�d��C��n0��Ȑ$j��0�wKcj�i���A1�������-���&żK������9���s�F>��G����ͭ5�S�oO�r�
ه)�+�P�O�:����2�ԣ�<��SI���c��j\ؕ�㤯S�׌V�x>"ӹWV�DX�e�!��,���m������Џ"�/�R��CKD��]
U�~����,u�I�[NOT�kꂫ�zh��ѳL��uC?y�q@XW<�7jP>�r��l�!������a�A��=����1��r-F�ߩk�G�_��?L�*wLNA�����Z�р��1� ��(#[Z��n�J"�[~��.Q�Vv���(�+��ǣ���j�2y���{�O�����:A~���p�������r�y��b*�Ԯ!������(���XWn$�fj~|n��81i ~8c�Q7��>�\,G��'-�H_�5�L��1ԦL�鮒�v�E��^b�*��3pPZ�q�LHZ|g*�Do�%���c���� h5C��&$���4D&�p)A0f�M�ddO�O��0�=3P�Vs�&Fa�κI�F�`��
^��E�{��Z成@(�.�zQ�:@��a{��C���͌�rq�T�C��H<;�� *� ?\��}��V���x���ZG�3[M0�$�D�ś~�t���ȿ	�z`�	�@�w7����>0ρ�r����~��;MP��^q�4�/�\'��0m8�9O��U��-�Ǟ���\=(� ́6���ջ�,h�Oo&$yH�œ��k�s»��a@.�3�"'� �@�vS�j�S�s��&n��n��B��Z��Hq��;��T��9RX	�]c>M���3�A+X0�k�����7�+��@�����LG�&��,�2�z(��>g��Ԙ}�޳5&�&Zؔ�_�Ų���X�ֺʯ��њ���/6��F�F�*�
�(�K����������|xi�~Ve� 4��^,��n���-���8����7�96$u5�A&:)~��M�_�!�-N��)�*�Gwt�O�$Q�wTo������?S�#�:��IG�5�/6�KE��C![yb�v�\a��?����O�<���s�r��kCM����e��2����}�'<�P$����4�T���gT�{�m�7����#ݒ�l�?�vq�
Rb�goVi�B,�8�!gD���F�p�:�H���IyO0��H�l;l�t�o���	_Y�$㋊�e������?4,4��B����yPn��SL�w�R�� ����q!�V�o�A]%"������m�s����*�UN6�F��:�;	�8A���.c��f$�n�eH��=�<�.�������q�;b��������T���O��4��vOO_�oȵ�
3��|�l���$Q��
s8����0��� ˟eC��?�v�V��^;�4��j=������&�&�Y�OZ�� ����� (�2D�@7IG�H(�$&�a��f�'���D݇�O)��LJ�<6��ϓ��-,�ױ0=ܙV��	^T�Ke��a)�t��Utn|3N�s3:�$֔�@j"�;1g(���8�᮷��J4��^q��J�m�H������W���._�����:��h�SM�:���k�>-��	�qOτ���.�u�0ق����C_����x�����9�'ʺ�b����G�	����8LSp�ߺ�����'��;��c˓�1�Ǣ�y��l���6�֩7T�ƥ��	�+ZY����	�m���d$�.�#~�eW�'3O>Gӓ�5�QXj�I�l�U��e�.�=��L�f���x����5���RCo��606��B����={���SU���M�p�l�k�m����	���Z�D�/������1��>J�]�n�K��2�l�m�%9��C�u/c=w�uOjyPJ*�^�\�橛�.��S�v)X։��!�ť|9���H���l�Z��cNE���4{I���ʍ�5������|D)��ZRP��W��z�Թ��N��:>S�kJƍ�շ�Μ��d�H�BO�t�A%��4Z=�U��O��gZ�7�s�C}$:�����wGN��M=֘�h�� ���H�����6�
̗��}T����C(��<{�yG�t$��|M�26k����\�����KI��i��P����+�O �*�����G��Ԡ�LTj=��#��u~6���W���������d�.�V_��?�p��9}�E�裷Uj���^�d{�^#���(`���g2��[r���tB.H�t��i���c?C���
��j�2�u�YE��������H����,�:&D?���&�^	��ժ�� y��8�̵�BsG�Q��4�y��>1Cs��K�����GŪ%o�Z�����O�y`/M�|��sA~�,�;4����ܴ���R���&�P̐�cb:U��<P�*Bp���jzm�N�^�c� J��˖���X�}.�	���3����t�V���4%/�r��|�	��hq� K�R5����j{fެ��;B�����g��\��`���F�%P�Ef��n}*q/6��Ğ⫶����0�=V8-��`B2T~L7�u%@�?�]S:�D�������rS�TB�k���y�Lc��
!�?oVI�ҹ��P/�"xg-o�g�E��8�,�U=91�+�l��a����܊+��a䟈�9��'&s>��7e9a;�O�f�'f�l���P�n�]�T�%��$��4B�RvK�ι�>��|	��)���-�2��O���X�{9��=��wʎ�76R�Y���H�#����� a��(�<�$,�S�s��)3:��5	#]�4��W���`��x��CUoc]qB��ݙ�q]�eP�'	�#�s�x��(�\���f�pl��K��c�6�P��Q�X'~��;�<ɵ��ƙ�����E�s�b�S�
-�A���pi�w	f�C��A8��ݡ& )���r��Y¸T8���q=i��8�v����X�%�/.����B���y2K�f�Ο����� ,v{�`�����4=U�s�V�f���D�^�9Ѧv��ː8ωp2j�e�24����M�Vňj�q7�|�+i*�1I�>pEZ��MCq�$��^�?����+�B;Ғs2��;��[��G4��t���i�t����/�☟�B������~�I��j&#	��D�Pcs�?
����Ł�}8-�DJ�!�m������<�*=���Қ�����ÿ\|�*��3�6ۻ:aنy�+�"�Dr����������{O� |�:ɏR���mx�<Gp��}j���cM&BC�J`Aǆ;�f(�Bb��_{WI�@B�9D����&g��6�`F�pL�)�Jo�Jry�s }\j�dӒ�.<�>��	��t���q�V��̠�63����A�1n���A*� ��8�d����흝��BJه���"��l`"Q��%���bб ^ F�h����M͂�1��y���N�68���yb��d;A�$�
��*�c+*B障�0�4.c�럼3ҳ���>J{���3�3���u	C%y��j����v���P-���z��G&ه�Ћ[���ɡv�`=p-L1�|/*!���ߪ���0��˼ ����5�D��N=�5rI����Y[�x�͞ϯ)��;�T:��lD6F2<���:(s*m��^�.������p���z�����z>��8���5�~as�s�Z΍&1�ٴ�)�G��E_ 8d�C�+����Ø���:��U0,9��������;2�}tp� �U.L>�>"��&�A+@j��|�]� n-�x�w!_�����JXf�� F��-u\a��m��ì
��{��77�����yz"���K$��.�B�LBM1��ծv��G�Χ�������ԤT�]�՝����Ӫ�\�[�'�xI,�^E�y�{b��!5%��+5��x|�eg6��'Ӓ;��O}�r�NT9e"y�=�#���,��Kh��rDq&V`p1F�T]=X���~�Д���/h28cp�j/��ч:���X�nf�_�������PҘ(��IO&�a��z,��S�����9��  ;�&}k�la��vDlM��z���|�Ռ�2%�|nD�~f�w�j����Dm�C��sɲaa�g�w%�
����i��סB�'��
�	�[Ɉ�����y�#8T�`�J��&Fy��F5rg��P��d���\�'�Ɗ�*��8�
i!w�G��]6C�=�����ۉ�Sk�[Tr5b�*'���F&o�:&���|���|����I������b/�(��p��7�`oM|5F\{_�����A�t��#ȟ�ޤ��G+Ds��vc)f���z>�~����IL�/=p>�?8��1��Q�c�����:��L�(��ɾ��딄�i	\}���3��4
���h����o� ��*�
g hEFI�oA�BmaA!������W�m�bL2V Y��i��B{m>���)c,�Y��>��FH���
���X{�u꣎Jٚ\�8S��Oz�w��4��Q=���pEW�Ȳ��e�8�xpL�)��J�����8�f�
{�dŪkl!j�����l�j�>F������]ְ�j�E/���X��j��~hW/Mx2�Ȧ��oE�E����>[c��Hm\�]㵗�k�H��O���]��ځQL�"��(6B3Z��ŎM�9T��GR�@�P��7��1f�7�h'��T�I*��i�]@aX�0�׹0,$���{Xa ��c-�������I�n�?S;�Z+O������`/��2�7@�^����L;�˕�2�C� �t}�%���@�H�<����AFמ�\��3QQ�6p����8�$P��.�J��*F��/��`�[,��>�©�P",Q���	ھ�E(��O�����;�\����C��j�)b������g����)�[f�Y�	�BOz	�.D�uX���2�����\Z�/3��ھ� �?*�~}�f$?/o'Y8����4�j�+�9���X��~��ڨ%_*���������w�p{��Q�:p-���:��,�6B<����@�'\)�;���G �<�wY�v�ꓑ\v�fݒo����آ�g�FU�32�^u���.@��)�|�^�-�j8'-wg��bx�a��eY�����hPN�vI���C��z[s2�Ef�G�p�R����O;�����r��eJ2�a X��Զ�/Ůu[��^��r��{�nx�쭁
<��D�����'�K�ӏ�k�	K2��<���@��v�,�e���H��s�{��Zq���z<�.���1�~1�aZȹ�e�Lf�kX���[uIw��������E�4���ɀw���s�i�Ro��N9QA��|C�v�p2�&�@��o�8�Ǵ�0cnWh_9�qIh*���PߏR����C< J�T@C1�E�Қ���)�v!EkY��(�/���{,!��Pare���wt��� ��s�N�PV �B�@����	�E��r�2v�ħ��MVJ�Q������ G��}���*C�&��#�z�n��]?7߼0����LS�¸ÅD:��o����v�W�-�g~.�ӡ�W��|J]�=�1�Vx�9�f-�h����?sbq�lM�5/x�*{0�f"�,�$^>�^3����"�"�#}�1�n)�6�JTܓ<�h��\����E��&�2��r�j�;�6��;jo�:=Q�Lk�v��뤨.�{��8�W�W��(�h�lt�#C��)�hxi0�|^�\��,C+�P�)0w�l}������H1�&A�R���; �V/)Sf��5�$ �Kݹ��l̆����qg4����:ה���)I��V����
}J�v�+/�ӡ_>��&,<|PE Ѝ��tA������L1V������O�^�FQ4�|���׊η�㚛[���D[[���3���1�gW�ג&��2��������0���3��o�+s7%����i�z�T�%��68�9��[8� '�w ��GIg��nRh��N�A�`6tn3�w�Cl�Q�o��' �ߵ$��OsW��@�`��TЖ�3f�[ĳ~��)�m�"�c� �S��/i��c`��)�������y��S�*GI��V�;��G��ewM�5�<Gf(���:H�\�a[�N�*7����i�K��]��f��7��;)��߱VjRޙ����y�q'��n�͋��?���ݞ	WKιa�� �{e���?2c���~��'�.����Sn��4ߵ�4�)��@�����t�`����Y�?��5M��FP΢-����TT��u~'2�Jm.v\!Z�i�c��@�)�
G I#�ey��S�駣%�� �ѫ��F�v|�}�3�#�V�q�XR��C }�g����j�	�pm�� �ʓ9Ԇ�}���x�5��hk0�C�d�
�\+������p��Z}�]LyE�Y��Y'��l���)2ɨ.kd��7��M��˒;����,�J0z�A\�i��T���q��j]�גy�'%�S$V#w�]�C>�gC�v��r�l8�rsf��I[l�,`�ԘK$qImݶL��O��'f�{���R��hR� ���{gj�_�[��t�� �0P�m���|O� fj����kb�:��JEd���5�1��}΀���V^
l��!c�T��5��ʗ誟I�렠���I��> �.��6L(��?W��O7Y�W���ƴ���z��S5.����sPg
2� �*P�������4�)ާUz�sӇ�U������X%��khj�Qo�ހo
V��゘H,l	2tuM��s��݁\���v��l�>�ݘPw7���p�U� ��� (W(�޶�=����y����eho��љ*��&�%�D�92x���!DI�^&�x�pf�'6ϘUF_ѱ�Z���p�P3����(�t��yX�3ؗ5%rq�I q�Ժ)�#n�[��U���W�_���cɹ��!�8/g����-�z��\cʛ�1�s��;�Ū�"5����|vwT���a&�M1c�:�sQ�]A�RLq8[�X�`t�j)��=��q����|�?]�g��HHr���Ԣ@咠�H���,��G�S	�󙽼�����q<�l�ͪ�E[�Y &k��@K��|���2�u�\���)����f�u������=����/	h�����H+��lSB[5b��x��AYJ;�?ֹ(Z���)�#Sf�.�g��)q���bQ���隵G�OҢ�D��[Ԇ�M���a�n6�3:�w;߫��Ҋz�]O;f�'{sqY�#�i��ĨFiIs/�»Ύ�[�e?����=菛e�xd�Tɛ����~{�6��*SqL꙰�x�����&nW�ս�a���B�{?g@R3��Z�"n�����S17���N��BL�"(6�iC5- 7��ȴe3˴f�t��
v��s�W�*3�1;��}��
��@fl6����~|Ѩ�8�8��8�?5v�6���v�@E��	z�~
��+���X�FIp�_�|:�
E*�_��a(�@��L1�$�ӳnq�?�e��-�	�$�,��}��6Wbp=j��L|��`����F+���GH����ђ�|�Y�z�Β���2<H��LA�wj�=���ҳj˄�N��^��~����z/qfD2l,�BE6�@bw ^V��%�=���WZع��s�SI�`�)hU���	�~C|F�@���N�7R۵�L����f"@���6]�R%o�x����k�����/�e�p�G�z�.�K�%%C�U�
Ga����V:�ķ-���-�Co�żr���um����y#:Ã7j��ڧ,W�Z��q��+ �"��pQ�����`/��ʎw��N��tG�2'��T�{�Ƭx�kX}AfS�4.���~(?�N/��r}�C�)�G�Z5�%�D�y䓭Imw����8�3Z��P��o�0�2�,A/�pZXrA�V�6qcl|`�ǣ?(X�ʢ�8��M&���:���
�K ��-TOx����_@�*����0�!�p(w"b�N�r�=4o��������
$��w&��a�P�����T�2��Ǆ����@�$5��ͪ�$zY��nZ�p��	�5("?KڒB���7C�kh����k^:=�HhQ]N!�9�j� �Z�0ڌE__e�*[p��X-���l�J-��c�Q���d��L	i���ė���DP���}��y͔[6��)���w����Eb�����ɢ\�2F����F�]��:>�����3	�I��ů�q5�-�䕻�1+`������1ͳ��@֛����&��u��r�u����Q�6vr�>~Mи���!�����"R_	�����8E�����^T'+<��R���8\2�X��EǴE�R�z+�6��3�Q���6u�7?�1��E��ܪ??Nh�0n� Y�1g���r_�-a��X��T%�m̞�_*��S=O^�8+���Į��ըT8��J�`C܆aA�4�>TJ0����p�3�H|�:4M=����Ƨ��I�4E��V[e�D�#jo���pv���=�/w�e��[d��Ҟ剀O��-<�P����idn'B������8<oڡ����>�Ҕu&.7������K��l��v�O���2�J�B�/�� �k�� ��WV�V�������Ņ1X�;�W�6U�{�d��/�i,�����%Xɥ�Ǔ3�];���Äe�9�^ә�tPab,�z9�YD�f�*�!��ɥ�#�t�?9��uq[�؞#�Dh��'�e�r�|D���̠7��9	��f�ߣ7b���U�q��F�Ri^(E�:4r;ٶ�eR���������In��j|�c�׆�}�,���h�p+�u]����M̹zv����2����kӯglԴ�x]���e=y�FU�:����!Hƙ7я�E1�1�ƈ �/>��G\Ŕ?�
�7���6e�1t�r�iͿ�ϗX5CZS��_O>����NR���4.u7?��1o���� `��p�n0>��'Y�ZY�F�o2�'#7#�w�f�F���VY��,�t�W4M�O>{xH؄Y��0��Ad��]o���®�5�I�)��}Bq����БFb�K��9B��Q�&M6Yڛ����w[��<�E>���l�	��?w�ol��mFR!�p�7a0���oTa+	0�����;���E�OLEI�3"�Lt��#�{��q&�rĆ���u�U5�+���h��d�7�}��o���1���~(n���A��I�����h)K0o.�<_� o��MI89�?�"�4��w�v����T^�J�f}���p+��WTr���D-�y�(z7o"�Y�Ҋ�&;|���A�����.�s0Xi#�`jS��o��T-�#Û/`�bL/l���w��F$v��Eמ�u#c=%��۷v6�4'���:Q�%�3�*�J��-墮�5��0����Ykl��|K�R�nSN܇c�čZPSW��Sf�3j	<�t�yI#߭'6�N�\r���y�T�h�ST��Uqa^�o�E_���EvU'�����.�nءN~H:���4����ߗ#���xw�o�X����Jzԋ���~5�����4��H�껾��ar��W����@���C����
�߯�L�˦~��}���0H�����eJi�a�>q>L#��K�n><o�~U��<,�)�Yzc!V�{���G�K�:+0���ß:��1&z+���0�(����k<v��?x83�ҟPv���D��h��}8At)��D�e�䩢�����*~�!�O2���F��?����̳��V�xYr�*�^gd��M��9�P�� s�h�O�'����������~�7�x3�4�����SV@u )N�/zm"��]����/S�q��,��%�o-d��b#��d� �{������ygwQ���8���>\v���{L
�XB��t��u�����R4��V�_u�3�NF�	�YQ�G<���q����ZJ�8Q�c�o!O�m�Wi�L5�[A�LH��;���#^R1�K�S�T�$1��?3��[,;>����nU.����Fb
x
ܰj�u|��������}z{~��+V�~�q�����-�c��[��
қ3�Z)�pߎ��h�1d�9F��^�nbϻ�;�w��1�p8"#e���Ǉ�L�cO�,�a�L׾g|%����n4�>�\�u��ߛ�&9Lt��2�,����y�$J �a�5i��ݠT���6��%��������<e�	V�i�V2��J��Mj>���J�LG�w�L�'S#�V��@������g��I�(-��{7;t]�gv�����6ϲ��d����~?��}H����wm�	DȤ'�[�������V�kImS{�u�N�3, ���#&TL��^_��"�ӌs�!�H46�7�=�@���"�q�����ߙ�Y�ڶV��J�~� ː�R���Yk�-Ԥ�)!���q@gq��z�H���Si�ٔ�}����䓞����4 �Pjl��zqX����;��R��5�m�2b'�ʙ^g3eh��?2X�y&W�{W�$�8�kɘ����|RmT��UIFi�g�m��,L,֭��_DT
s�_Ȇ��{��������M���6)Ҹ��qI���-�u�e�n@�T<��x��Ŵ�E[��K4xB݄OA��E� �p����h��K��vJ7,|�l"	 ����4�pmE�=�(���@pkl�ݢ�d4�SP�`��D1�$|H����������:���?$������+k�;�>9��Տ"a��A��|a�S�;�;�y�G/
C��]����(��@����e�W������v]���'�̴qϔK�g�qs�45�W�����PK��N �I=1�$<�[�v|1����x{�hXؕ��H���FQ��X,I����XO���|�p'�E����G�Oy���`�F+)zf4���E��&_<% *1{�۶v��O��\b�$����d���dJM��҄Al0�GP�u*��O�A�v@%C�4����ص���V�1��8�A,]0�M)6}� �qƼ�D^�^���-�*�o��i�#���e�3�E��J[h( 9��8���͚��C,|���l���цK�Z邕����p'���Y�o�����>���`��Haq<7FJ��0r�d��̋��]�.y��3_L�v�� �x�繆�H.�������s煰� �3�jP�J<���W���=q���q�?��䓊��v��������Xc< Ն������/�֙�bp�8.��1P"5}���vH�Яzӗ��
�U0z=fR�`���"V�i��͢�$f��-��.k�������&��m �@�^�q�7�CcN�g`Z�r�U@��˖IjL�,)W!�dNL�-�ˍ����о��")�7��=��b B�z�O������>m�i�u�u�D����@r�&{��z\�����q�
�;ΝPlFӝeU�Z�� *�������l���n,���O����Ιkd�L�D:(?��Z�Zdł!PuU����t+/�aa������r�<*��dpSQ+?\h�|⓪���Գ[��Whϗ��z���jC`Fp���%S2Ք4�ž�2�MXB���MI:��d3i�J$�"���l/jS�I�I���m�$7�vٛ�r�8S;Q���R_���j��vN����1Y��=-ⴍ;��2����BJ�@����
������|�
�]��.��N\�W��uPV�C�$�!@sm,:M��gtmP� d��p۔Y�=�u�-:�!EyF����ϙr�oXI*��n�wcOS��@�A��A:
'u2P����l�g�`����=m�$���2)��`Oҫ�Ȧ�a�e��'8}������P�qq�
E9��wُR��T�x���`8OY�����{�Aɪ����Z���
�Q���qN�Х��<�.r�\�׵!�Nz������Y�}�[����yS�?���L�i�`��-�1Q�ˇ���f�'?�8���P�Pjy�HmU���J��P�e��с	��9B+@)r>٨��z�R��3yV�Ȇ���/��%5���U�@��y%�Z{���g��}���U����e���.�ZM�I�����2۶����|ߪv�4����}��ʉ{�D�.��Ϋ��.�c-Y�5����m*l�$�Py<�n;?C�7���1H\�׼G� _��\��ܦ=(�=k��qc��Wk+C�?�N��8�Sէ_ey�<;o5���cy�Ή̈P�(����	h�a���!}ۅZ[�	k�c�8��S���V�%�͸O1��Z#pz���;��\����°��5V�
2�	���@�|f�!(	ɽ4��$ca%�0�8�[�Rb��Jӷ��v��q�h������2g��O��*"ʍ���'��k")~���h�kƈ����*�멽I^�&oǉw���-��\�-ն�5~�V���m�n�H`�d'G2�J�X;Y�2���r⦾S���+X����hrT���2�Z���pj�&��T��l��D�]�@|,�*)�x��k�1�(ƹ�]�+�g��u(�Ŭ	�|q䕙"�v�ZuR��{ A��y	���Kl�PUzm����|���1Nq�]7�l:T�-\�#��f-�k��?#}I���i5��d3�{�.7�'z��WqĔw�L�Q�A���'M����6و�k�k{L�(��*
OxX���1N���R�r��2��}F%]I����uR�h������O�>�7~~��/�����@�Sf�l)PG�4�Е�:�]4�m����#�ޖ�h�)нd0�ܸ��6�x��L\�����92�(�5�+�����1��o�.6z��b���A�Xn������~$]���`�)
4�M'�߻=k/qU���8tN�W/�Cy�{am"K?��a{R����kQ�sڢn2���2�1��5�w�s}�ձ8�.B��k����ʞ���n��R����ǥ��DB֭k��}�������~v�"���[-Fk^����p�Q��4�SĮ��.�. �Eύ#��ݽ4/���\�����
�2�O[�������H��"��?�V��=:S�0��	�'x���1� a!�V\�eG�,^n���fcvC�Ģn���К�$o���c��6��^1�:]�������E�SK!�U��7=��$�X{58�Μ�*P�+f�>��q���)�斃?�t�%��u	i��i���e�;� ��C.Hj��K�c_d��lp��h�Ў�ؿG(f�f��u
R�5۾?*4�ծ���g��a���2��=�$�3���f��b~�h�	!�a��%{2/�č�6�#:�U���|<Is��НP�u ��a���SC��������#$฾�v�؀ �,l� �������}�Q�h<:]�a�I�D5�;���51�zK�i�a]��1L^2� ��7/V�#"*�����EG﹘��k'�̶������SFIؖT{G�,�w,������JR���� }d�ꓳ�ɗt����*�H�%���C�4�߅G;�G�(���,�=pn��q� '=P��}kʘ����#+�T��n!U�*I2}����<��D]U��v��+Ϫ8��I�Y�E�\R���eG6����j�ѻ�ڔ��=U�q����n0wG0���wN��"��҈�<�ɸ MÉ�Rbj;y��|��}�?lk>�M��1�\�{�{s�����yNؾD\r����j(Mc�Z�V�d���2����70r�c$���;c�Ui�RO�+��D˶��n,��Z�Ò�IRMp[\�ow�-�V���6�\�N��Khݸe�v�^j1#���s�;��%�"�l�R P]�/
0 TD+���e�`Wn�!O%�&�t��)�I6��ݯc�$�p��XFi��u�q��<����dF��U2iB�"��5�-�zNPW��Ҧ��F�V�NLZq'�;�7��6ڵ�F*�q�$���.�(ݡ�2��G����G+"�djQ8ND���dV����J�ȇ��!o��ɢ?&�9�#�0p�a w�S/��m|��zx�Msg�C,�P\8/��#a���Q�m�Vf�����B⥷��o��+�-�w��FT�8"�n�����������&�(uQ�9��� ��*�<򦪅	.�)��_	b	��ްz��뀹�d]��Z���r�}I Ȥ��^�����_�j�9�&6M�裦�asQi�`�G�g.�e�s�	�Hмt��5a�bT$maX���A�.r\z��.�G�|�����Y����YJ���E ��Y��w�V�%�n�*�ՊC��EXg��2`G�v�^����v��G�+�'�w��.�2j)
8P�M_�B��Mw*��dŨ��q%����u�j�����j/�^�UmA,DW���5č4�^�m9qc�a-��!�
�d�D
 ��B�Ki�u�Pj�Z���U�ו��g$�̦��� �%�E��>FJqiA�Hb/�Ƒ�q�"~ ��w4�A�(g�4��L�=�Ŝ[wO��7�=�N(�=�eCӪ9� �O�]���s/F�U�_�L�?��!	��l���o��s��M`^�_�Im�6�6r̈́ۡ�m�U�r^�ױ��(D"����1��s_����G&ͅ�Ww��g)c\�G�5O�el�޾G䛫8n��Z؍�/3�tSǚ��`�8�*�e��r�����@P��ݤ�Q���?�h_%Ք��`ƋO?58���.�ʚ:NQ5�G�}}��iIͻ� ��9��
���,J��G���������~���
��x��� ��G������\��h�����9d��Ѐ���YU�=�}�������BKh4q}�w�j_��9ζ��p��8X�*���G?��"u��UZR����p\[.!���G�ׯ_-��~�9��7��=.`lO�I���<Z&����q���m"��u̷� :R3�#�@���9�#DXt�4�@����n�g��13n���6Iu��W��������W�� +�H�PGmD�d8^%-F��_j�u��3��ն(9ѵ��38�6&�L{v9�VWj�9�4��r�;�J���EJD��,!���v��2�Z�}�إ��ҳ��IF�9�iL����FSr>)6��V��R�-ZDj�4ʹ{��k��4�.���p�4��h�=}�-��fi�Q���nU��O#����_ �$;Z��:�g+�ı��}%��k 1��8Q���9	%���_	��۹՜�:�G���c�`29ɟTC[�N45�B���\��8��9�����m���t����CSN<s2���Y���6���g�D�f����c��)F<�8��l���w㔵���V_M��Z�5�>�ưh���^��h�Bm�(6�̖�j~�!	k��mu���K��0��F���R����;K��1E�a`�I	�N9�K����[1ﭩ��?}<~��du��m�3��5{��O>������Y������;؂��ńu�X�G�Ak��-�ē��ZC[l�U�8Rˍ93s ������?�>��R�����ϔ-�蜍{��B��p�΂�Vs�q���Q��?&��Y�$R�����?�=,�mb��X/z�nG���m49{G�d~��r�o�S�D<����aw~)|��2/�m��.�T���5������-�T������~m����/U�r�#g�����>˧�ߓw��ޢ�bzʍ�Mq���*�wQ���
��o,�B��+��s�9`[M��hx:�,	��dr}�.%��:T*���~��9_Ub�	LK�1Ϣ��֌M˯Y@��/BH��H׭�W}J��?v=�Q��\��a��.l0*F���ѵh��.ա߇ah]��]�}�$P�ܚ�h뤷��C��Xơ��+-V��H@��ŵ��
5 D���=�l
$J�YԈ7-�X<ψa���~��x���(���x����i ��q|�y�|U��_��nq�%�n2]�/Qx�#�o u���\�tj�'8��a�̤��4�����.q��⣸h�z�u�N��)1����]�dw�I��Q1��T��[vCԖ�"s;2>=�]tg� %l���#���>_���o���;Ϊ�҇8SR�L�`���tf���`R.>�ξ�����-5	�Cr�E���;I�ם���a�����0�!f��6��wz�Ay��=��S�����h0�7���'�hC�����D�t_��@(w���T�w�}���{�ac� W��=�P��[fM#]fu����᠃��h`�ʢ���X|�.<�w�x���(�}H�X��)�H�~�Z$��J��Y�zS��A�v���U�O�D�{���E�A�o� k;���1����g��HR��2Z ա3)�� ��Mh,��l>��MJ�F�w s�{�S��m��ܞG4Ŵ�+���qr`�x��x�~]�_���ݖ�D,��C�O��x����ce�C��Q�b����E������P��X���1<Ka��Qx�Ǭ����]_�ג
�>�]����1����`b��&��\�l��\�EII��<ݕ��i͠;f����f�.�< ��&�_��$h��cC���+O~�Kg<��~�3�n�`-jQ�0!~[��=�����o�꣈�nQ�l2��|(�q^?6 4�u��f�a�Z���X�`?pȞ�Lt��O&b~9�u�g~f��Y��ogk�^�V�1���u�Hg!i(�DyծA�Hb� {f�еK��-&Ɋ~k�@N�����vU{Q�(θOZ�qֻ8��x���J:�]6��ܞ�&F��ڦ6��A�d��θ��<�r筿+X�>]w4Y�E�.�\8�Le�y��5GW�ۍw>�c���0;�U���-���B5��u+�p��x�6�>���f[�p��l�@u���l�)�G��e;QfTP�� 1�(�@����X7'7��żf[)U���uJO׽x�C��o�c7�~�����qE�' ����N��T��I�.&��
���IucD�]62�5�K�8%����F�}N�o�7C�4�/Y�p/��yS������L�9:3g+{ʝ���l({�y�8�}Z����v���q)K��i���i��	���ƭ��%"�Cn#��X��(��*�������ls��m`Hj�E-D#�C���"��"@9��Wx��ፌ�-m�B_����t�[��d����o�B�>V����������@a�É.��{K�qw�_��
�jv�x��̀_@����D�שP/��A����N,z&�Q�߸i:�2��L&��K��@)
�C- J�
�b�0G���$���=�-6��63��6.����,<8�J
=Ц��)Y��΂���B��o�`ɹ/��45��o	E����%�|�`�sh��\���F+�gC�S	YH���#D�ZF�A��+>+5R��O�g�Ŕ�.�s���iP����s
���ܸ�P�	���p��nS{��W��T�9�u��C;��^M9	� ]���7���Iҽ86�^�+��-p���u�#Xk"Q�&�$��|¦+�[���>�
�)��:���Y����l�������q�ϕh�t�:�7�A��އ"���*�3=2��zJ�w�` c�b����U�����Ӷː��Jƽ�5�!{��ΆG�d��Ń��lmu��Y�tQE�������f����'��� E�^7�Hqi��R?X�c-�Y#�77�T�DW+-,�G���`��џ�Ý��V�#��Ǯ���o�jI�qL񖐋7�)g��kCT܈X��#Ys�+��l���3y������` �"H��Įzd�!��MK?�g��2�ZM.�p M��D��܏��=���T����ft�D��a��'�ճ7{�O��;m����Km9�\ʐ��"��Ix,����ų�u�,��ę}�Ʀ�����5��<P0}�m���|9���z6�9�@yBgf��X�-���s�uI�J<��+DW�Q��S��{3/5�����-A�W�˳g����|�:O�\�l1o(fӆ�ءC��H`��n>�K'�(I�z�0L�0Ry�qS�n��W�0m}W����򺸈(���5�����5~+3�z�7hZ���c�9����&O.��Iz���y �0y��R��G��Ïh�L�p�3�4��aR��(rD���j���~���R7ߖPĀ��Ǚ��K,0�hR�JO| ���i�թ��4myԲFc����h:��M2'H\�1ohq��ԥ����ڔק���ΞbKhhX)u�J,�U��3g�o��Q1��р~T�`�P��!��+
�?�O[�]y��y
��C��js����|�gXE!VQ�-����P1%�ͅ���sB��`q��~�\mpDC�-�_��=1����F�Xj����,����l��Ő �����4��#V������ X>�ꦞ�&n�Y8x��W��%�$�Ç�����oyj�j7�'B&���4��B��v�Q��-~X2y��yƷaF�
�H�{�\���?+�p �����NB��,�
tz}��=�B[A!�E���[����̞v���@N}�~�o��k�d<��cI���>�a�DZ���Qw�S��ii���<Tsy�8����C�<��AzO�*Y٠�T&&��2Ԩn��.���bn��d��S��Љ<W��hy�0ʲ78��_jFS�˕BbSl!��*�ZRw���N���)7󅝪������Q �^WC��phF�r�ǁR��v���v��X-h�D06!�i8Ї:� "�Fq�p��� 2�s	��C����t�2lA�1��WX���#m#9�W���0�yu�9�҆��/#,K����۴�_��iÆm��(��� 0����,LR�L��d� �A�E���n������1�gs�-���.Vw��Sy׶�<�~����@��t-nwI��an��\�9�@e��e���_�8wfe��R4�Fy־�-.����-3Ɨ�^�j�@f��ب���Ύ��� c�t�έu!�x�S�^���m�9���+'�o��쟂�8��J�7���7[�B�C |c�_�1vZ;�iC)��B}"&
�JC�zt���6��T~x\�\3Ms�_��� ��\�����v+P�����Ll��I;�|� (O�j�}�#u�����(�����r�ُ�):���=������C#���}W%~�"#�c���δ�ZM+rJkw2�D�^˧��Vc�Xy�U�v��U>�����?�ԍ�l�͗.	�|���=Z+F���3es��Y�s��,��J鿗�I�L´�����,���	���̺KD �g�ax��`		k��hZ�E�Z���9,�m$��x��7|�>��!yj��ĄЉ�{�O[9G�IX��{�u�G�3eJ�Ed���D_�عEE��W��n]jI3��)6�U\x�\�ў �^�5S��O:�;P2��N��Ţ�;�y.|�?�s�/�콐���������c����L���*(�;�d�2:W|�m�y�ڬ��'��&�g��8��=N��k���J~p�%��c���t��+m���`����^{F΍x�t�Z˯8ێ��?�3���]#`�l��7�un�J��FtI�!r��b�FćF�L���|M�a�*����_"5L�1EQi�wΠ�A�]՝��LZ�?��V�h*��3:�ij*%G�98�"��~n�J�>�[����ô8/?�J��Փ�5���S�ۛw0�ֵ��6�Sk鎋V�A$.9KnW�5E=J��F���-��08���t=������nbi��ǧ�}�c�Y� ��L��P+eGڬ�����M\���v���K�VonMb�e"��{��p8@FOo�O���i����#!����~����.Q&KT���Mw�����<��IB>i[S��HHB��F�V����T��g$�l<J-�5-ǀ����5����vRJJ��K����$�[d����vB��+f����S�s�?M@g3#��%eQF���?m�y���4�IJ�*��e���{��f�Qt����Z{3Ev��ט^7�:ۻʼ�3���0c|� p�������,��}�4����e���Ș��b��u+��V�)�����Yj�M�~ajq;,a$٢.��;[j"UxsN[���8�8�>-S�d��Ld�I ��0������~R"-du��óI�I�����B4�-w�й�e���b��E8��m���C@	Ni�a��.���Qȷ��&��
�Y�|���:�����3�(5�?$��X���>�,x��Jt��K�Z�lp0uDB����&}9�S�����3���)��+'�_��<��
�GWd_.~��C��Q�}��j������C�7���}��+Ft�NqjZfQ:RF��#Օ^C��_I��b�S�-B�\��r��h_Q]�����!5?��{Rޮ�8���u����pk/�\E�+oMK`)ǬtO4HIc��b��i?��4�\j�;��2O<�+���aK�EN�ra�6����H�>.�]	u�~H�͒��834��O�,��#��Pg%q�z���;�#>� ٴ���PxKL+tZd�Xc���'nx����1�p��N���dNX��aZR~}x��2��H��H{_��oSBst�4ڋ�i��{c��ՈP�������p��q�[��O��O�߮��6v��eض�$�i�����3����Z:�A��)���x���..�OD=�u�#��j̑ ��Deh)����ߎ��fܭ�3͸l�4�a�����������> ��g��6�D��w��j�.8��T�D`�1�$�F��b���k��-l�I]��b��t�`c��f��w�$+�t~�R7k�	!F���9�,<�=�l�B��`*F�
������W�'��K*�C�L5!lo� �a�A'��r�i6�Q��n9ӂx��gy��L�����c \��ݼ�<+��ŋ��?_=3v��z�Q�uմ��y区���*��8e�<L��� �up<&єQ������Z����Ȭ�%��vߦ����P�Aޓ�~Z�kMuJ�S�f_�$ʈ2Ź�*���������,��4Z��v�x���0,۽[Y�H)�˘�4�u�6ˁ�%욄�9 ���Q&��;�Ea���y��dwހ�[3�	��P��D^Y�-��Q��xDv�6e��i��y���$��5c0���@��3GI:sk�!�:18}Z�v�MN��ܽ�n��|�o	����{n���r���_&la�hO��6E��np��Ȫ"9�s��T��Q�G�z:�B� )7��J�p���6����I�}��ʐ:�w�v9�W9˰n�Pd���Ҹ�Bl�΁F<���i4�b�luf����LmWw���k
0�q����ëo�Y��.�����y���:ު7��bb�|�1�g{;������K���P��m_�GW�b��wR�A���p��8&��Չ&��A7BLS�N�-Ԧ�탞=t���ʽ/zJ֎J�ƣ����IMb�q�A������Aŷ$v��)AW��԰�/F�V,|F�P�w��ET�(������jX�]�Ւg成Z��j/��Y���)�'���9�8P]���]7^��ۂ�\�Y���Ԕޯ@dn�W��	�l B����v��n�����~��*�ໜ���^,���F���y@%���1��f��9c��L�d
������1^0Щ��*ڑ��gx��g�Q62.���	\	�����qgkcf?ե�d��\�5�D�.�3�E��Ɔ;vVS�����f�-��@����V�\�{sg�H�C����gC\������`�=���sw�=v�ˤ��(<"���˄\L�<�$2N�I�	�cyQ�-��YS���E�t-����l�Kp�{O�~7f .4M~n�7/A�I�HE.6~�+X��.U���sf��*3w(zr 0%����@��x��g��W��گ:R��z���bB��9l}=������$�muO생u+���e��o��mԎfuE�o��V�pJX#U2χ���r�T*�i��,�+@g_\�ozM�e��ך�Y�wF��1���a��w(���L$<�dF%jNS��i�ZW��9$�2a���T�=%��5@���_����iW��J��Y��C7?0������qȭ=J U�
�/�'��Ց��x�����DrxlV�\EQ��@c<�IКk�a+z�N�z��� *T�TYR�@��T"1Sc��w�O�7�ˑ�z���<��޸W��S!C�)���6�Ҙ�:��5��ŷW�׷�����yӓ�JǸ��l߆94bRm�����φ�$���!���*��T���C2i����X�}���,`�ߧ`d����M��,��,m͔�o>Ls.po���Ͻ~���C�)	�n[< �� �v6�?cI)�X,!�-t-��ą�Q��?�t��@sR͋:���#a��9�^��@�&�=T/U�x���F� �'���4(S۟E�|gfD�!Q���I%Iy���S@���?_&	��f�Dx5����(��g��V�E�2A��G�@%dF|�J��8[�0�\�HW��+rO�\�dP9��9��)�v��郥�BF�dw /�{j/�enHK`QP���o0��ʎ��_�M���O"�O��ҏ_��j:�����~2�s1�'���6$����+2x���Ϧ:'QC<��x�;��C����_e@�Z���`��8m;1�]E#
2|)��)iE�� ���SJ�3oȸ�W����tPB2��G���HB��r������o�tk�&�m���2�l�,X���+?���[X뉑�1Oy=�ņ�Tύe@\pΔO�v��1�����]l��vBc�υ��f��I��.bRo�ଇţMk��5�0�V`A��w�H����������+�%�0�D���� ��)n����B��s6����i��<r��F��+�K{��X������u�J8Rgٹi�K�2?�)?+|��G�k���^�+gFԁC��M�<�B�� �88�r�E@0���� ӎߘC���s�J�GH��?W5��|!���^����'�!.Ot3v��U �g"�����y?�,���Ep��]S���a���|��{���nV�����q�OV@�����ϤR�B��w\ض�3�>re�(���0`dF)}�0���q¨ƨGv�탌��w�o�����a�,�[6�S/�����U���B���k���YͶ��0T�A�p2�����E�r鴼�� ��ԽlH��'{�$:G��I!����W�y]�V������t���E~
9�o����vUSD�~��]��Z�<�*}�JP��[� 1�vX���:��(�3�>y�c7bX�.ܰ��޶�<J�D�K���ִ��!|�(sA^��>�����C�c�����er�B���{���VDd��MR^���Pp��08�U���_ �gϒ���iz�7FNpG��PYr[�aY����&C�u��~^̆����%�&d��?��ҀGޥ�J]���v ��zD�-�;����B4-�0z�}!t7"�j?Ωt�0��j&1X(��HN��5�n���M�m��n��g�!h'[�s`n��u�̉Z��)W-�_���sٷ��M;*
nkCI}ր5&��U{%e��$��_M`i	�^���4���ؖ;��u��P�����0�ΤO�3�Dt���=^5����t�n�K�9c�����w���
g`t�B?�cݷ���"���z�E@�M����a�v޿{9����>�.�v���F�i��%����&�4�&m����6Vs���P�l��g i(8���a�j��~������t�\�|��[��Ց���L$d:d'tZ�@��X���?$l��Е �m�T|��1&��f�70�W�mM楜	��;�t'%����!���������wgx�}>��~|�����P!2�i_i��A��0�7b@���,�����v ڧ�cHO^H�6|���c��p��}l�k�V������%�Y����NV�t
�.9����[���8`@�1�fUك���:�ۚ���WO�^۠S~���)ÃSV�/����b�w��T����`t�ܥ���`��JCqy��:������S�wS�blM�����Sϖn���+�S���3�[ϐ��h8��Q9\�ױ����H �-��@��jS姨��J�y4�C�aQյ��Ȭ�Q��*�'�#�]�eZc��N�~�Tꄜԥ;��	M��p,����d�p�EQ=47�W-q���eA�;)��Ƞ34o��D�܊�y�׶#�f�e�q	���o!\���L����ʼ�N�N��� ������\�K�P����*�G�?օ�5�����b+B�<@�˛��s�'���1��w��˔>�`]j�9���A,�%w�}�R�π�����4@zo롼�u_}<�i#��B�IȄH����Y�@�bb�>�o��T�|�t�Ҵ~X���O�qR��t}
0&C~�J�n@BU�~�/�25�ƐGXo� �����/w��	����#�CK ���V,IY	��d�l�+�56�b�;�*���2a�$Z�T�;���(�]	�o�ϿZO\�A,'t[v5�x��[49���)��^�����Hu�: �[�!��/��Ϙ���i����_u�W]5�Ϙ{K�9?�*��)���BSP�c5�O� =S���d�F<�{������`�w�K�7Znf�D����	���.��*Y�=�z/}�Шnkt�Օ�f��p�����u���x��R�No���.A����2p{�y��"�V��t�%yZ�����[1SAZQ�[֞M$+by�����"��(Toj$�B���\����������Ք�]�T\����.��:����
��
BzXW��[���f�|�m� ��:�	��v���fG
�ȅ[[XQ��:/M��'f�I2�u9�S�F鍇��X*�#�m�)ZGhDH��Zy#�f4�8�t�j��vS�j�	7�.�Î��󼾻mA��YIvB�G�?(� &���L �|�����������T�=
"U]���p�;��I"�2-���ow���j3�$���K���ʠ��uF@洚����&��"(0τw�_K&NR
|�wZ�OcV�����Qk�a\
�r#9�����,��a��y���0�#�Н�n�t{�S[W���|�v�2y�;�L07�#T���QE��_��Y�^�-�]�!{Y�:h.�j�aڙ�+<���R�fp���?3q<�q��ro:�uE���5��4��|�i>xͽ,�kI}��F'��y�����
�Y ��@��qQ��(��c@�Yw�����;Ym'���m,����e�Z��Ο>:Q�e�6)+'�1�vZ]��i���P�m�y��߹ �Mou�]	͈A��apJ_��_�Ŗt8�W�����}R ;lCV�P*�f���"����"�ٴ���-�a?��r�#�՛�-��ھN�
^�8�����	ɫ��`G��ߦ�'FR�c����&E��U�?$5WQ_�t���Z�@�r�[���e�p�A�8�"��(�I�\�������BC��V��H#d�ƴcI���6s|�	|~`e/{kĖG0Uڹ-��j;���%�P����4b\ڧ��D�5)4�3w�����X�
z��5�31���]x����Z�RMu
;(H<��w�[��2)��o]k�p|��׊5���v��;qR�0^ߙ�icm�k��Z
Me����q&\_����g��&��R�Ce�l0�"A�T��� ߳�P��<�1W� �£E����0�������[3 �:��V���C^�S��!59	o����
�g�:��V�nDL*���'�/l���4��[��9' a�ɝI� ���A���LC&B�REN�(���<k�i_��$l��Md�4�u�D��=*�[���E/BH�P���x���pՠ�"���Ï�����d���c�
�7>iX��`Aȡ�j���ٛ��~��w�"�]&o���Y
����C�H�2���_m�\y��A�>P{#/��`��K�	�G�e{��e'~ �X�2�08�t @o�U�a�v}s��V�����A朦;�d҈t�hz0ւ:�k�]�+N�@��`<�v�2'�F�Bh�F߷&Dg�/�'"ϊk�G�o�,�1�Y+`b4�2���F�r��}iZ?�VQJ����a�e��������-B�ɢvN ��y#Mi��f^M��/���8�[��B�&?��P�_%��?BtG����`��,:�8_J���"|ܚ���Uݡ*��ã�&Ǔ�~��48:�a�S-{Dh)汃YCB��[w�(Վ���'��0!!#�����煤u=���+�]3o����4p���ʿ�)��B8���x�ڭ�L�����r�`_��h����%�R��8#d7'�1�R��Կ,�a���%^D�.��#{�)�j�����N e�ն?��,Ъb�:VO����|O=��w����	�Y�ڥ�5z�";� ���3<�'ܐv^��y*w�z��7k����)Y
OQ�Ӗ�2/�I��
_O��m���o�������)�ќ-�OЮF`dt��F�;Oq��ua�S]�`X:����فD^�I>8_���k�Yd��io�h��<RQ}�k6����������[�:b��@�S��B�ɉ×9Ul\��*��zb�S���l.^D��V�\��'�y�LX.��-��R6$��'�,Z98DJ#�p	�l3� "XA�z��攅S��/��_`V�4�Un��{���A㐛�
	r%�̻~]��+9�pZM��^Y6�Ŧ��k�i�#e`a$q.��M���3Wr��X����Q��ۤ�a2ڈn'�c��u�SP��������u`�ל�GTʚ��Y��^��M��f0w]����!��eY3^X���"+aCY��_/��e�ַ�$u4��l��Na��gQ��>� '&�/����A��G-ih���/zQ�K�XV��z��)���7>���U
�k��38V��YW�DO�3��=���ڣ��zɅ��F���e?�E����i��̸X�|O��%b�?�_&�&$)�B�(�l���N�j <���xxX�7l�ɂ����#��{��W����F���f�:t�� �]�~�����ԋ7�,�-w2�P,���<ӳ�l!Ԕ$]�<t�w�^��qo��o�����Đ͐�W>ݍ��x�d�~)�'Y�H;9�m"K +E��'�����:��Z��L�@g�>�KW�d�L=u~���Y�;sX��\3��0�[�DZS����L���
ǝX�>�`>�g�0��t�ԃv�)BD��lo	�8*r ����>ݎ!)�l�pЋ<�J1�����K|h�3{�>��l�V�tQ�8$:��b�iSv�Ͼ�館�7����VH��F7曳i{����kW8����l��na"5�W&N`yQ^�]�~�G$��i��Q�YI��Ք=�ŀg?��}�r�]�����t�u��ޫ1�t\7ߓj~�S@��<��:>(�0�ͪ%D
�<�%f��H�i] ��M�z�Py��B]�)���68�2�i����FΘ�*���r�)��(1���q�j��´mE}o2�Lh�����u�i���!�j��n���H�4�80�E�<tّt�!B�K��V�z�YR6��*%�[��SQ�}�������q�_��	�5�֑L���
L�ɩ4࠵��������.`f�M��;y~�X�So_�ej�E��p�+�p���,t7Y�Z���X2���nW���w�0�bh�?ͷ��u�:�{f����h�n���Ǻ�5'��&��kRI7䇇ݓ}���R�1|m��E�$��b��#�ˆ�f���Ss��c�2 ~�	�Փ�܆:A�����Ѧ�V3�5��F�z�����(��J���M'�)0�>{��^��QT����M^�݂0H��ii@����h� �1����q��g�p�G��'	ɩ�����>]���)�pc�A�#śt8��.���j�v�?,���_	�ߞ�G?�䙧�Z)�i2�^��O��nHh�K� ���&Ҋ�@\�J��9�+��zUZ<�lr��?"B~^C���E[�7b��:�E�{�k��/)�Ȍ.`�a�oDYJ�=�+������Hٳ�R3���\�]�)sm	�n^�G�֣�n%	P�d��lSn�Vv�fR� �v�X�7Nr�nͤ���؆��%Ui�+?1��&�V����)4�RG�p߲j.���#��)P h���E�]��6�xv����}�\�!�AD�pm���Ce���q�	��G��5��>!�O	���"�;�{?������-�f����_Mv��a�u����H�h���Ur��,Lz�e�O�9!yߕ��,Y	tf�D���J-�wq��F�������0�y�P��jD	ZGփ�F}`��$T�7�\7d�G�>��ZJ�lwKJ�����U���+u���gE�/�7n�D�1�(n��8����b9��96\՚8T�L��~}6�0�&
�;�=�:��x���&��\]��\����W9|)B	�7���2�I�3���:#p�z�<��,����7��4o69�^oNw�
���1�nC����%a�s��p�Y}R��Ǚ�^��Z@���ģz����7xi�~����
~���A��=�^ێ�%�Xʋ%�@��o�-Ct9�����&-eZ�i�ꗯ�%Vȅ����P}�[QҘ��ڟRI������f��Ln>�Z�m�i�S�®@H�M�~$y֑l��n�!Lю�5La'逆n��$a�5��=����E\�����;�NK�$Qe�7d�	B�rFйH���ܖ�U����0�R�PS_$I�U�}����sc�Fy���x?ףIZ�����F|9��i���c��p�ƴZ��i��O=��~�7�lSO!H*�4�]D�W�J�&`�\���U߻P�t���Í�|g}�!D���:H���p������mo+ ;�(�计6�-�侜�
.��pIq�jk��$]�0}�O	������L�ju���v�U�[4B�wgo��ӑ�J?m��Z�"����w�9PIj[�9�ЄF�Ĥ`4v���~	�Inq*H^?���S�:��#�v:�K0S#�B�:𤾕8"H.Sҫ�T�@hcЂ�bd�ԅ����A�d�e!T_��u΀y���!)	�C��({�����# �*_â�������&r1V}d�C`�8�!���A4rw�C��|O��@^�I����TbS�@��-
{��?\r�~z��LP	��<1�k�4l+]��\���-dȂ�o x5�)=���r�O^À�`kZ;�#f6��>�0��ygt]bF�=����XX[(��`�)���+�K�n���� ��+�,FƬ(nB@◰0��1��Y��[�l'Vmإ���x_u���*��{ܛM�j��C�����$t3et�㒲G��C�DG�J�������dJ��QK�R���8Y�8�<�F��`��9�����t�m%�M2� )�nb���jE��q�����*ܨH8Q�wg��`Q_ߵ�ˣ��h��<_dA�I�
p��n"~����炙��%�G����t8Ah��.ÖL
J�T?���*�'�w��Sl��y��H.wp�kԧ������:_��&���$��;cO-���& ��d��"B��:L��шh�H�S'�9*�̀?����̦1���S�SD�W׋_��d̫DJ�W��$��4�I�p��1q����u�r� �{(y��Qa�y�$��,�~,�\��4W���\|4Wk��~�w�}6`�ܲ�����ds��׎<���i�k��$��պ"��}���-P��͝.�j5�?y�T�3��m83<���ASڙ=�����#��$�^&���N.8w���5��O��\��y�zЂ��-������������n,�x�`�z�II���ڦ�-��ង��L2�D�?R!�8���Ee'8 $���BD���A��҇��tШq����v�����F�Q��{�p�)���3��l�q��{�*+���(u��B��(a�@f��z����=x�H�j��u��s� ��L,��g���9o1Kn]n�gf�r�,౫�h �C?XK�Lc���n*P-��\j&��0@����!�D���%���W�#t��	�=�#�Y���W����7�$�{�C5�~L=�w�����**ywm4O о�����ė��"`��[�Sr�nzǊ��i
��m��'_��:��>K�֦O�������M؉f�n*��1��U�����vX��'�^.]� �"�1S�M�Z�^�	�
���`l��)����L��MJ^��>�<-*�3Z��F[F����m��u7�ٍ��am���<J.�!3�;rb3��!B������6\�o~{hQ^� ���h?��)�"ay6U &vD?4�#�Ä�N���O��0!p�����s�ȩ��_�{����=���='��M� ���&�$j&� �'i&1�=�m��N?��I'�������c?��L�|����nM��C�b��/����qݕ�>�Tǅ��@QW5����QG�1t�����ٖ�F	���{9m�����p�]X��x���7*�`�g����|p����;����FW:�'&��a..`&D�n ݴ9'%�+������p���zzK�AK����Г^#�ޒK����&�q$��e��qUѳ��]��R+����Z%{C����?>_#�
�q-�0����I �E_�s�`����@�[���w��j��9��whx����{|˚����=&k���h_�󀗹ϗ�6Q�[�[ ��۬>�̣��C���D��o;���s���6}>����}�P�Nb�Ks�ِ�a�l/�4�&��{P�����Q���Df�]��^����k`�v�Q�X47����o���H�G.S�������+L�����iw���Q|�p=���p�[:��%t2����M�-Stɵn0�q�x��.]�o(��t�IK��v&�}�5�ʁ��ꚙ�VoՅ��s/�,7��#�J���nQu
x�r�j)�KZ�] ��Np�9� ˙�ʷp �0>=.��]���q嫋AQ������n{;�����7��U��*��Uf��x�t��{�����lc�~���X2��`�N��Yh$qh1���N(��l7�<:)tg�C�c���Q�I��M���s�H�~��_7Gk�0Wq9�t�?�>�;�P�(��
/��N�"�&*`�v&��R����_s�Xk)��[�Tޞ���)-I4A��� 6�t�.�%��I�5GKx?�Uy�2�v��q���?}◹�H.OjY�h?���,��<����;�94~�T��x�;7��bx�Ԩ3��EV�;��bk�:�5�>Y$I(�|ق2{WA���>� �20ު��\�1+,���Z(D���T�76��G�F�6'�{�9�O{#�&�]#;{ߖ���Ϝ��ȄI�>���_26G�]3��ǌ��=Q�y9��G�1����5��W}0��	���i�wan��D~�[�}�����gf��O�&�C��CT�f��W��.��3�O�`��u��7o�%S��]Nw�s�N�,٤��,�K��<ŰPK0�!��x�V-�����k5��F;��2w���(IY���f�>d�_���}�а\��wUX�6��R-�������������Q�D|��i/������kAI�_��>,e��f�X�f��Ct���K?G7ݸKc���#��ɷVʗp�� �L�V^/HH��9O���6���P%�k�$Q����xuB9��f���	bE��ň`����%���1DX>h���2���I�,�u�]@�N���*�o�T���a��NB����;~�����*�( �ݝ��M�rER�W��pO��9w��07�I�"��H�ն1�OC�\��ʡD ��ٷe"�fZ�Uג.�F�_��L�W���l|"2��1��ܿ^����ͥ�� R;���4o�.]>}j�Örf��lZo��]U��7�5dr79]�vv��{�)��z�;�\�N 0R������RV�*�XR8(v���w��fD�!�����=�md3Vz?��Dd��>-xs��1l,=��f�4[��V�z}=V癖�c�yW�ėE�����!>�JW�0	Ee�|p_Jq� �Rq>u�}ZZWG�)��%Z����O;,�3Cd�ϵ_���2���p�.��/�I���k��%J8�kP���� ����31"��E �M9L+KO���%�G\T&�t�v\���+k��0��Y>o��r��1MB��Um�NdAGs;��ȥ�
x8h�Ec��6 �c��lu�Gۣ����R��y@��T�5 ��XCH���Y�z:�]�EB�wM����������Fc/I�Ƿx�"f�9ֲ�T�S��@6�:�����՝(�d�y�9����~�&��~x��F �����ࣃc易�S@�������'[6p6�(����jk0�&�!�r^A&b���;��*���o{<�қ�}P�����Z��4��1�H-L�>7P����#k`c�2��pk�˃�;���)�kǛ/�Q�98�Yxbu9�"��4�q��[1�f�u�	����3e����iDRy�5���S�6���$=��նa.��T�a�j�DO��a�?t�s}D�)#���瀍������w�OP����";�佤.�6�w$\�\t��3[=W�����P3���Ιof����p��)��+P�Ŕ���W�U=K��m�Q�	/Cz�-���$l3~��*��Z�I��)��ё�p�DĂ9���6��>��I��h!%��O;�)�L��Of��	�699��=��O�!�/H5Đ�]��xX�,r3��Ї�q&1��HNy�Tt�68�S���:��ߨb�y����n������|�6I%����t(��+���$���]q�=yw��/��b7a@����β�;�Q���X����cV�ג|}��U���<<��u.uy��|q0��ױӊΐ�[k����)�C��v�a��i} [&��/	p�]_��#�z�~���*�G}P�$��Ց[@���jS!���*�(&�۹��:,8�J�l�@��L{l�4��A@Uo2��j���r�"�J}�8r ����ѡ#�"�U���
���R�Sk���:P�zr��y����/����GK�ٷp�l6�S>�+綆����3�VW��f�ۮc+W��{V��d
>�I�1��;|��e�=�����)��ߛ���~�)����F��t������������-����5W�c�b��}]^�2�,n�S�:v�[�Č W|�"=:cZ'k�A�E{?���Cn���=�#1^�u�%�5dprfr��la���h���2
as�	�*6\��]N�GI&@OoBq�h��j� �}�	4��x����VN�\L���6!ͲJ~�7UM��O#l؁9���@��M�`��	/?m�\������ڴf�q��-���Q�K Xg�Sc��آ�\M��I!�~��8:�P|[���}�Q,"��\��K��h�����]U�Q�������\�H����h��p�)9w����r��\�"�⟞�-$�����ѿ��QuLo�L���ȜP�����-�^���S�><�-�͚��ư�3��w��<������	��^�~S�`LH)�>UF��&恐�:ͫȴ;r�� )�'��ɗ�Q�PZ�u�\��ye�wn��>P��=�w�$�D7�QQ�ޣ d�R�Ī���wJ����8�}:N��qW���f�ؖ�̍m/ �ٽJ�����a� �[�
����:ȅdϥKb3�KۥA����5��՜����(�?�5l�S��W5=c������A�yn��R���8���	���	�;�!���)ܙ�����C�1+׫�����Iվ{��3sX������>�z�D��:�aLb�*d�$Z{+�?o�9��udd�n��SE�]���u�/�+��������-��,�R�4��H�$7�{�;v7ì�2dO�ٶRJ�Qj}Y�$�?��}߹��h�x9|��k~Ѡ��{��%KM@��F�i�K*t�����jq�Y�r�u*�/n( r��8�������_��A�����m��(%�K��?�v�M2�H����L�*�������h������ڙ�h�&7���2J��n��耤gu�W͂����Q��$��+*�q�(6d����A���5>*�91�xb4�8W�>�1wB�r�VK�����N���p��,*h��ơ�-sj��g:iP�	�u:����p����Gc
���!x�~��|B)@㌕�M�p�H���Ϫ�� �?󥼾�����۷��7�
�tV���I(�ڈ)���9����k�|��3b��iC3�!�ڱ�Ǝ��|EC�'�^A<�y��}����VЭYi�G~���0Y<H��J�����9�󀒯'?�w~q.a��ֳ���w�{��w��	�ڒK�|����z"�1�s��xm�� zHy��ԏOxi�.$�B�ɪ�W�����$��]�؝���Яe�)r�g�8� a($��c0#HP�6��F�����|���x�V<A�7�QL��(�BX^C�J�/cW���y�lG7����w��ɷ��O~��C���kǎ�;Q�|��3�E�R=Ѳ�I ����m/�B��^H{���۽�ytNX��+6=%�܏Y����g'<C���_��hE���_BA4Zhb.�������;Ch���	]�t�!+eSR)��|0l C|��>m���#](�/�o�e��1�����$�����"�z�2�WVXd ����S'sA�6�g_<N\���\�]>�����2S��\���D�9Hr'���Һ���D$#
�7]�R�Vb�[�1#[�|J�t�QOd�|Zn���X͉d��g7ѿd�e����J�e�x�;�aH2e�h�
,r�9��:y�H�A��6��%k�V�4O�;����n>Z�4VPg��4-�/Ĥ��|�t�c��{�+K�>C��;Y�F!�9�B&�<��k�N�)��>S�)�$
��B�c�v� }蝠p拷
�򵋞w�j��k4�䉊��z̏���۾P�8~wx���4����6e+5���GCm6TrPtŷ�
�GYe�2HY�NO�.	���� v�)d� �8x����D����w��w�R
^��c��(Z:>p}l[���ڟJ�N�����{Iw�s����S^�ܞ�4f�u¨�
j����y�X( �_�;\.ЗK:���r�H=B�wpC��z5L_��b1�_�.�g�m�4*��.�