��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���'gW;�9CaE�h�\@�+��
1D��q�H�.1`�T���4�ß�ư)2Z��>ڌ�]B�+"Y������Z:mBE�Пʎ��C3@��1~Z�!���8�m8���e������A6<�{e�q���m��}�2LPbs�=R�|P�X�ҵ_W)��[��)�U��x-|�p��O�oJ�+ði}�d����}��[[8M���z������N�D�m��o�O�"�y*TG�J��]8��Pv����ц��&>�T�����TNn�Q��Y���v��l$F��
��z���Pw���z(�hV`��qO�q�PW܋(�[�]�O*Q4��%�����I���Hc�A�':(��N��8l#�R�W�����Wx�2�˜�g��;fꠕ�����oJA��6��n@Ց!ncT�܍��e���lr������G'�ߟYw 	F�f���l�"2\Gk��UM���By×�+�0���bF]��wC��9s�q��,z�{�o���|?!o}X�f�P��@f�K�:�U?P?d ��X�b��_��H�~�b>�ճ�Xh5�R�g��4�|e����rX4fo!wÂ7����!E�����Y$L3�|M_f<ւ:(S 0/�ԑPEU]��8C����y�Dw#��V�@�#�Y���Qy���d?��W�2+������Ҍ�4�v֍�8����0��iZX��U5#���,��W��`8�U�x�<Ǖ�����'Zqx�%�6[M!¤$uVk�R.�SgA=�"�ùH�ʂ1rA�k䐦�gќ�x��l��2�Jcbv��g�O|7��4~���q1M�i���r�ǘ{y���յ�Kƨg���u/�M��M���~��E|Q>KPJ�\p�xRXN[)zB��F�/O�H�xWk�B�@��u��irsų'C��ʩ
tz9u1��! ]Z�-�3Bb��VX��|�4I@��h�:��AlVQX��%G�Z��t��{x��:J#�uA4I�~���ٸ�3.kl��QC�k���&�l�+l���E�?��+���!<e3.�z�t���PGL���+(���oU��׀#4�1[��5��d.���Y�O�'j�O��5�k���Bj�7�}�0�n�l7���˧�|�0�"�����3��.�C��vG}h�ĭ�l5F?��e�q�UL:�A�! Q�Ho���ɘXާR����1���ja5l[;$��~Gc����x�F%#'�m�s���ڱN�ݩ9����z��	�hf�ػ\��:�fquʇ�y�7b	wZ�������[�:7��5��(s&@���=���yy����j������h~�א̠�x�Z�J+�6�_�\t2�چߌou�HZ���f5AO��q�72	[���1R���\Y�!�/.by�(Ul��ar�6ik�]��}=K�=����jȷh��H��I����@]K���O����zg��gAj��~��>���RIl��9M/ۭ ��֋����Sc]�H��aɖ9�Cm§�G���az٣���({�#���U-uA謜�8���:��鴯�}��	�.��
��3�(����V�+�(�����x��c����?��Vqk�� �V	�<�2������Y5�]$���[�}!M�MY9y�B�

�`|�lW
�"�xQ6����U�
g���M�[[�g�T�*.ِ����ܬ>�U��v�<��҅�'GV�nՐV��i��j�tj�A#�K���� �a�����GϽ�M|)�3��M_h& ���~ettv�hk���ej��+k��&#����cE}�Q3s�ʻ��	�4�����.�N,k�p^�v%`)�5Gp����V��!�<�SlI ����G3*}ܗ���J����W�}��j�(�����@��K�}3������}c���ɒ�E3kiG���ɏ>���ͪ�{�r�yQu�Ya����LC*����+��@��O[)Cy��Oӥ�G+�������3P
*�yN���@�!͍�C{�Dzp�W+|^'�Q�Y�s��:�t�­�e� f>���S�=���Ӎ���'�P���K��U%/��2Ý��w�d��W~J<�(��x��4?���?�$w�	��� �S�	�\��]I�Z�����X�f2��c�ܑ�cNť7�Jo��4��G�s	�?ٷ��W��`;n�� U��@��U����\&U08���1��)���&�`%;g=�J�Lx���.,��)�4*�R~'w;���t��V�tm:��nCpm�.��ι6�ςD�0��:�)�ëdL#4��gbVM��z�|l]���I�f�BQ�u �b��mE4�θ�3�
�Û��R���v��M���;	��A�n���v�Ѓ�<�/�K+��xe��f�.��J���4���1�:p�{HT�BXO�c6As�=��8k���r tR�@���{A�]�#Pdw�G��݀[�����%�b��1nݾ� t�Te��E��	CF��	�����۵|��eg;� qg��R�4�(�JWi(DK���P)��[�aD��:"�x�o�F�gO�yJ��pͭ�|�E-���(D_&e�*8�O��o_5��)�*S�a��`_��u������oh�ݪ�&�D��W�Q��Bl ���oKۖa����q�7�O*^u�>C3o�r/��R�F1@ALF2VeĔf�9Ug0�^��^�y/�-5�W�v�w���f����_������6<��E�̈́���b{���Ԓ��;�6Ij�D+�k���C��D|������M��h��{B��nqʷO�<�]a�W����-X?�p�/�+q8�kYn+���v�_���%z�a�o��n�bֈ�h�5˞K�3��M�lw$����� �}��}�{�L���	��Y���V�!��K�$:��=���޵*�E�D�R���=�����Ƹ��7��gF�B�����zS$f9
^'H�"B��r�����d�1�� ¥ �"�{a���q�]��B)΢F_uH��+��ߖ|@��^�@u��bܾ�G��{Ti-~���N��y�JK�LUa����/�{��$*�Vc���x�I��̭@5F}خ%��']�����h�ue��R�;����ٲ�p"k~�� &�J@g���2�@�4Z�
%!�M\�����|��:��b[=��� ���¨��aoH��7a��������Ύ��~��J�kڨ�46e��.D�Wx�T$F���nX{?U��a��B<<��s��cj�wJ/��Z���5���Y������֙�ݚ^.�a��?b�i�U�S̶��9*�|���:A�2� �/��B^�<�]i,X�:���MSS^ ����G"@�b�u����[w��
�'2�%Oy���ܨ�R�����������e�s����ʅEǈd�v1��uG�p]�K5����kM\gx���.�p�KΙned��]��׶���)����4�����ӓ�u�����k��_���%�p`��%�P�e2�P��j��27���.�I�&(>�� �d|�c>����J4���B!t[#rk��S��U J��►�#}<�DiF\��r���$�������F&O]g�ѽ�x�ޯ��Q���:�Y�#dZ��r�������"G����[��+`��(��"8v}���P��[Q.<,�Ez���")���ݱ`ǬO	<��E���ƒDG��<��a����M�rA:�x�.�S�OmY�$e�B�phr ����I5���A�Q5HW���Q��4�؝G�'Rm�'�9�՜��:3(\Uk�t��FT����Qvfi0�Ů��vL>�wH������Ē�0U��A��*UV�嗶�ɐR�C�<D��/l�h�*�o�"b��='f��GtK���Gb��y!��2��(ѧh�d�G���X|Cv�"�uw+�k�4�(�Hʸ�}ӽ�;�<���c��x���U�+�X�I�U'���8���iTO.���仙d�5���)��PʕL>s�vx`rd���c9N9v�z�h�i���7<�L�{�R�i4FsP# ���ƹ'^���W��8������N�^��7�Y����|t���}����~	�OV�ӓII~:���O U�r�p !LVQ����OI��/fJ%���
� �us�J|p�?�Q�N��xY\�\�H��t�-���NE/�]�5&s<�S���ғLD*M�pQ��B�����@�
@rܮ�Pb�E�$�5�;>����p��m=�$c������� =�
����\�LU�vg�ܙ+u ���7yv��B�{tў�_w�n{3k�k_	��>����ΐ4�r�*]�3��a�3��̏�Z�V/<�7I�L+s35dUy-7��,�q�/˾Z��=����:E�T�şZ���҈��H�Uo�ߧO����d�M�sNh�yId�1�]b�,B�i�iZ]�f$t�6�~� �uX~.��)�׫��4xH�K��E��h�@P��ջ_��ɨ���'�l���'���{���T�E�N�^��pr�)�����c�VdG�����3�v���5-7?_ܽ�(�mP`Ǔ�� gT���m��������������B��C����({JΆ!�OY�F;���Q�� L��@9�9�
�n�
8�DD�<�ٗT	)�z��Q��:}��G��	�x���Jװo ["�+4���R��\V�n�Uڲۡ�	`8�>����ֲ�.���xyǆv�d#T�s����Χ��đ&���B�2���4~5D+��o�/�������"��?�'�1��6g�hG'��9,�s����W�'+ւ����+��2*{��#��2�N��ϯ�M��!��1Mס&YО ,��
 "�"�+�o-��1&	XO��)�"и<~Nn�ti͹�C��)�6��z@;nD�ʏcV��Ѯ��d�V��䶂��X�
uc��$U���]�f�5��e��� �Q�vJ(�d�AveKѷ��u�?$ĺr;��w@��*���"J1۩�H��Fm��H%�k':�U�0�����t(j[�H����%f�,���4ɦ^M�F�;�@ͽ�`��[;�9�#�dZ�+��g��rճ)�>�Z3���|���r�o�=}����cFK�����R)��>J�p�hQ0�omQ��ֹ ��V��:mjfd5���mG2�����: w_��'o�?|Bz���B@���yB0������ɇ���R�,˭e��Vރ���CiP"�K��A�)�]U��D̍|�<�1�����:y-�t��!������HE�ȟ�S�\<}��]��x.�^>�	B 
V@��=�l���S��%8i�p#栟��g��eY�[�&H]��(�]GsN�/�atٰ&׫|]3T���4<�w(w�Ŝ>��?�:��٣j_k3'��{q���[����<5m�?�G��$(�O0)�,�2S;_-���M�Ω߿�fR�EcfW�n����:ܡ��@p�\umr�L�.��8��e��w�Vp�髱��g�1G��W�˸$b���tf�aq�E� �_�6��a2�j�^�뚢~2��"^�ɍ�O<�3�H@F���&n�Lx' 葮A��7��	@�k���˥�uK��_N"�?C��_�:P�mɝ#Q�u�.R�����dA��Z�$K�ZV�X2L��4JKF�1;�f��`!-0!C���d ��2��oaUoGKf^��t���.���^����Ë��=J������6���jKL�"}�N���ۗ`~�₮�=,K�Ǆ�� �&@�.�f���>}7��Jr���P����OHDm/8�"{а;A�74�X@T%�f���Op��h}/A��({���l���*i|/�~+#]��T:�۹�%����m^��n����UNq+?��#$�{�[���+ojX!�~�oށP�0�:�� ��Xڧ��˖#�����d6�[��o��+2;<S�ە��0Bp�c��y�/��N���\�	Ml�� ��u�u&L9KV�D;�:�լ�UTMB+�2��9����
hW_�(��0�����<�Z��xP�à�J�;�=�!1�C��,��EDYL��5����	)t�E�4�e�o!���
�u6�ԑ�v��k�MI	,qW�}� ��� I]���*��Kw,2�z��0}c��Ѵn(�L*�BD�R!��\~�t�$Xav���)�����wHM������槶a�zwZ�'ʱ����V\�L�'��}s��� <~P��[|oRu�Ԅ�p���oú�u^W6��z���t�{?���OZ@�3��ʍ�Mr0��'�oо���~D�����YU��D�FP|�Ʊ,�[�0?=#���Δ>�l���\1�U��:Q}{J��
��E#�|�!pqٟbDj�9y�o�~�+j��� ��o���cHXE��+�p�?�NH��o�8��&�Y|�V����.c��������sK=+b7���T�w��;_ȹ�E6&���mlg���/P@#2,�˦�)�Ly�FG��6�#�-i�!��I�o~���J��F:?�K6x3�e�Y۶��~�c��1� �����g^�*�0B��lY�6o$BO�O��@�4JՅ��(�g�*����8�����^AI[)v��.(����}�pl��}���e��Au����	�g�	�;'����ԥ�+�1������
hp4������.�Α�ޯ[���
��5jc$D�¥�r����,��>���%��s�-�ns����T&`	IF���Of��%q���2L�f��57;��p����dJQ�`�j�9��~��am\d�S�c%�s���jS��vN|�%�Ac?��D��4������n�|s#u!6�'�"q��4Rj����?[#r�˺C�l�9��ΰ���v	%5lI�1��}w��t	hU���l����:Q�����;�]��,��t�S�h�����%����5P_��G8p(.�b;	M���o9���{�;�Ne�[�ٖ̪��=N�@�����0�;��B���v�?���@�gƳ�I&��)cKu�c��_b|��"'�mfc壨�%~��A�&��*�hC^
j>`3�s�L�r��Fr�ZZ�/�n��ݟPz���aWX��j���S�Kˉ9�>���\���	r�1����p�{��Bz����޷.���� &j%V�:�P�7��>R^t3p�k�=�N��ă}�7��?nl2���'��Ȁ7.i�ړf����[�{��h���d�M.���>�bIlUꊍLu�ב���zW�,�7��ن�$1LN�y<>�8L�:���\\��m����q�1��X�zY�Bf9bPm���AP-�N�0>	���4���o�8Z�p E�+���*����$P��Ub9ʬ+j ���V{K�MĿ^��*��M���t�|v�'J3����fs�wN^8!��uB��s�mȀA�y�S!݃�k�26�Zv�<�;~�~
{{�6D5�]@���-Ɗ�#(�0�],�u�$ ��wp8�+�ęעN��o�7�	�־�?��:3��1�/���v\��o��ƀ.!��W؆E^���N]�c(�4<w*��j�+���~-'��SR��$]����������	\�%�^���A���٭�q�S�s���߮���n'̻��iQ3��v/i�p�}dK�2��8�����J`Ƀj��+�ٔ�}jg���Ӻ4�"և${��w��J�^�Z5�LE�S�ˮ�A��]�U��(�:���-4�'��/'*�T'�_��C.��s�-����@:gQ-��;��