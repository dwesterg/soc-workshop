��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\��On�������F`��@w�;^�f�0�E=�)|�q�`��E9�1Eu2��I�rɽ>��	�Leev�G���e�}�N9'��Y#"_^c�?�&��4�9��O,3��S��|������)�p�@|:�����[�^���&��撡}钌U$��kК�J�}M#��6]���o%�("�q��k�����?��0 }~o"T��do`���	���둷�j"����/㏣�ف�ʘ�AP�1!�6@� %0Y4q��Xp��R�O��K}�Ώc�~�&nn���Z��[+�n��?	ZL��ctɀ�f��
Z�Tr�=�&	](��
�ʰu�r\�����)�߅�'�:����fTMhuX"C]�(ߞB��M��͞r��]lkh�7���	�5���B�cnp07[j��"G��6+����E���Q��r%຃[�'.��i��_�,]S$>ME�w�`�ʶ�9��X��}��S�zx�d����{?�ѢbZ�p?�����O`  R� o���ג�9SQ����/1�M�g(��P�~T�1�k[��YLcf�b|�JJ�#p�Iʓ� �&[s�H��%��CV�}+�	+F�]>�Լȷ�����:�cI�h~�2�٣0���뫊%��[z�d�Z�9�=��Z�x�1��M7S����.�\��R����/��L�}5Z�Ч�G�tA�W�a�� ��5[�I��q�XZ͌�7gel-��~�0��Q�4`�4����g��X@ֱ��SU���)~i��� B0av��U�(̳�6[���uW�
�\����?��I��jP$�y$:�%�CN�k�Ŧf�+��,v�>�뮯�C����0O�	rõ���a61|��ȀW���'�uD-Q@h�d��#�PV���4P��>��A�S�#Qvl``����Y�����a��IfL�����k	Q/�P6��gs@�<��W�O��M�GjN:����d�c4$_8�gK��R,S��jG��i>��n�-�:�K.���dp&�B~f0�vm�@���4ȵ�72�+��~����n�"�^�_��f�C9,������Ǣ<����dp��7�D����zes3 5tk/ĸ~m�}zb�hՊ�_����:�;@��B�{��8ʀ,��=�K�� 1�(3ĩ#	>8i*h5�4�3��׃D�!��(~Φ�N�U��$�$����c!<(�?�TDT��nJ�R���Ip�����
�H���
��������ʕ8�(���W̧�?�s~�1t�J�A%rJ�;+y�Z��C� �(j�G3B�Dh�I�@�X��m1w\Xˊ�a���LKU���س�!�|{VZ�!D��u܇W�(�Ѫ.�8��w=��%�j4����76O�m�N�酃����uQ)�RT�������v[&��ƚ%2 ���6T~���|��L����#�1 �R� �R�⽕��wA��U�Y�c�%Z������ ����z�y�l��e{w��Դx�
E�m�I}�Rn5�[E�A��ڍ�L�y)e\:�l�G{~t�2L����t��:�_7UNE�O�_i��$
�!ƺ�D�d+7��[��9���_�ˢ�o��b�cs�+9W��'yWn9e]2��.��������uZ�w,X��'<�r�@�I�"��	�>�;i�6��P<T��'�ؕCV=��]ƉyO��y׏��z���Q�2Y�o�@��~��d����CY1��^OJ�`˩�ճ��)��r�F�7*��]EZ'����+�F	<�E�)`�x�3b��G�'�q�������&,Λ�z��v�t֧�^D}�ؘf�;Ӝ��L0�j�J�AAEMJyk��}�>���
Nnb�,5ȫ-�����&��(�s�˜l���ci!�}��	�|L�����E��߅�<��zP�S˨������W���R�֝)�"[ Ę<)_���`��!	����>8b��9���r��}��%2L�7�`��̖�=�&�e�(N�
K��҈~?�iĆ��Vx���}�?�FF��d$,K\EWY,�aG�S���,�_/��Z��o 7��D���U�Y�ϋ��E��nN��b�\�-��}����x���f1�b>�w�)E,=�P{P@M���=��_O}{;�>�rP�<�H][r�����`S��"�ݐC�*(�F��.�i_JM���	�]�����@�!�u�k��W!�;�*�2e�j� �97x`�gV	@[o�ښd�WT{���R���?e��R���t��Ue��@gR���' `s�&�=uf�@�2h�� �����S�q��=_��xꖌa<Q��4tmɂhv��ĺF�9c���~�d&�(�VV�jR�4��2N�q
�,�l�'�g����g
e}�3R�E�O�94�9��:���z@����)��̜,��Mt���D���o>���_'j��X{��:/\�gބ��XV�eT�rà+�Ugy�u�(~[��	�`����g�����V%V,� ��)��\��ߑ�%�2,��ѩ3���У�s�d+�>�r��p� �5b2��Tۀ�"�@W��j  ��JI9�=�_�v��M���U�ʵW̹t�n9&�]��
3Ά(�ޭx5Yb�ʵ|���O�.�(#�re�������Fg |^�Ud� �	=}3���߉�.�H�A"QKi��`�c�_lp�|��@!�����YgU��z�
~I�2�ԭ�J\����̚L����l_�����4gn��xD�=���5Lúik�UB��j�1���Sq>��;xX�n��`V�+_���bD�'+�&D��~헼���.~�m�&��S�b]2���k���3��u)��T����j�<�7�_�����$���%��׆��	�:9� ����?�����'����ugk����C�,2��s�*-�
�bTBFy`��+S&3�B	�兣���t8��rF��dG�bI&im��jdy���h~u�����Y�, ��/Aݘe@zd8��^`�wy@�u��#�B�˵���g�N�DE�B�9C����q*�^Y���;���'<�@��FQ<���� S^o���j�����ߙ:���X��'��H�
�Q-���{!:��nW�OҨU-|\����M!�O����v��i���]X#��Р�sLӀL� '��Іlھ4k�����PI3�Z��"��[[�;��M.���v�v2R}oPA��� ;U���~��Ч�nmXT9=ݥs�8�q[��9�H�uZ(^�,�Z=�����o�k��˓�η�o_ܠ{�4�t��@
�`��.�u�2<pp�/��+�S�k���R�?쮑*d?���mO���l�<9�O��Qs}NQt1�w~�y�D�q�k�r��^
)D+wK���~�A�Y����u�z;��b�QڟG9��4Fy�q��D�| >16����[�8���|�y$�	(�m'q�\����6;\�ɑ�pk�n��{��Z k*�;����م�)ʹ��h��q�gs�/|,��j5�G$�v��ۺ����YЫx���C�J���q����g����-?0E��R��y�̦�B�'�53���)�X$� ��5����+��Py����w);"�'�E_v� 	�����\j�㠁��4>��A��_s�p�7爺2�0Ҫ������J�D���&r�e`�P³��#p�%n�V$'�����μ��m|� �E�z��Y	sc�*ZU�����2�\��#��͆p�{xb�:�y��JϢ���g\���t���G/1
���E�E�c�C��)z��dVryK&�����y �Zu��;mż(N�E���)~R��ua�7�=��3�i�uu �/͓lҊ{:J��9���� ^�M�~�qD�n �6�����|�*_��~���y��� ����S��U�3U>��B4׿�=���<b_9�����$ˣ]�NͱT��f��1D�c����+������`oˏ��ює�����?SDT����6ƪB����⊜���`�Eq�gKx> (�m��l���R����K��ܥ
9uK= uG<�l�hG���E�X�p��R�f3Y_O��}?����+�ک���"��V��7�J"���rԋw��u��R�+�pUh�>Q{�RF�F��B���l�ĩ�M���2�֧��k�����DF��çğCڇsNQJ���(!Wh,�$d�'��Oб(t�,��־�����8B�ɚ~+�����_*^dy��/�1Ō`�@e��,!먊��t�`�1�x��Ok�&��%�$ZĿa�{������DN��bx`�zǸ4�+"}�k�3쉂X�_��He/2%!I�`��@�~bJU�8�l^s$�I�?̙�����񺸟�2�F����.��o������������)'Й1գJx���tAQRk[�+;k��@�7�65E��8si��H3F
_Q��&���9�/Vi��L�>��w��@b7S櫸����s��U�� V>R�[�ݚ�k���|sJ�۫�4���wV�q���'�=����X5.��'C�=�:m�9�W�7�(�G<I ���6��P�w�����d�����kp|��� ��`=7鉎kY���k"�J�u���P���d0[��q�q��_�ۓ�`T껮ȇ��3k�����`�!snH�A2>5ᑱ�Y���	W2�6�ߏ�Y�����Y�[v��ڐ�_2��0JE��J�b��Ю���*�fO�����4k�g�	�Qu����Ѱ{��ޯ����z�H��0v�^d��t�����;�F�J/#>���I�;����NZ���m��oԼ�����_g�Ig��,��ɩ��)�rZ)�v+��`�"͍eV�g���	O����>e]rO�4'u�v�;$ �Q�F�d���1�]���|gmhJG��*�w	��h��ĿP퇃߰����^�nl��8�A��� Q�f@U8���={�	Cz ���Q�<����Hl�qS�J�&}����|�|��>�����en�N����q𠯸����T��O�����24�$�2�<���`>B�H;�1J�����o�Q6��$
���yԃ
4�8-���}��{�q �o^���L�v���<�����PՕ�����J�0��IG�VH�6�4C�BIgdRN�5'��5�#�M�����i3�c�0
 ���@E6�Яf�f �"ඉ�&8�<t�5��\��q2��z�����ͿE���C��p���p�����Vé)���E�� +0N��������+�M{1�[��C���"�cI�w�ۥ۶f�o���t�g�j�>3���kK<7$Y'2u���u�F� ��
f�hXS��W���@rα�(�5&��@Lk%�r�׍�x۫�F8TV(�Z����p��2����E�6�kH��=>�aY�J�?������N����^E^�C��Ђ�����]ܲ�K��G}�	�>�̪����Qnu��..�QY��Θ�y�*�n;Fx2c�HWn�sE���Z�+�� `;/<ts�	�L{�F�8����qI�s%��W�wg���]%p��K[�FMw����4>��x�8���t��_%���OH ��ʌk��?>G+��F��X)!S��hC2~�����K�>�� �;��w�kW*�z�C���oZ\7/�B��k^3�F�E�s� �(�L��x��}�*>�[M�V>n3m�Ya|�>���n�׮{�oS>�lGV�u�_4e���XBo+w�KK/�.�#�;uQd�J��y�C��Fs x�`\�\ÍTϰ�z�KxώD��ON��ۀ�Ψ7��0�����S;�
�-��'�Tm9[���\��(�m!$Y"B����'�iE��y���)�	�ϙi�Y=�@MVmt�������L���*.�#d]`�kFS�Ri��������,:��>��G���$->�~��ٟ^]ة㹾qZpg�ZDNR��1EdFL}��~�d�<�5\D���僷�N�tma8����=��4�8Q�	Ƈx-#�P�Je�>�٦WĵVz>�yTCv�r�mS56N�[C��c�w�i�����������?"��ߎ`Q��`Ċiu��bwi?L�E�K�����$�|��=���(J�Ó���he�,Ck�A�3�̭gb�BVo7���_�tu&��׬6�{���Lx�������P�K�RD������t�q�7���)��d�{��. �:I���mVX']�����m�D1U��8vޢla��ćq��e�qēϋ�0z�3���͆gR�t����~�&<��Ö'� �ߢc;{��/5�x�\�=@��$E<��(���h�G���\xV�sc$���3��kmj��ԏ�7_�x��,k�i��*�����V�$����j����?�&m�����q1��(rn8-)i������#	���:L%�l�
$�d3���"gF�D:���+Ғ�$�!�7��k�GL?rC��:ۿn"��5���d�G2m��Y]�' [=�1�g�Ui��RKc��A���"��Q�X|be��'u�!�ֱ�*j���f�_qh��E�ÞZvƎON�N zz֑?}��:;w`r.T���5d��6�RPp��wҢǢ��	�X��*8N�͏j�r* �#=�y*Ñ@i�|(5��M��RKs����J�
��-bC{�6RgO�_f�$R$h�i�
@z �T���{gC�mM��������9�y%�����"�n�.׫8��z�?،�5��Km�=	F忋X����ֵ�}�%*�>�NQ�x��	�Z��Zћk�:�GEo6w�W�of�	+r3e�_@S@�#���� :)SQM�*I)X�d;��d��҆"p7?�u'�a�dŋ+�-���A ��l�?���8�l��Zr��A���y⧑���D�B&��M��؍7#�+�M�)}���xo�}\�l	���a(�.4^~*�A��� �'�7J�Tp�g)��!�4&�%zk��-,m�+�s��F��HNvߧVg��V����f$�=yS䚩=��=�HȌ-|4&�kޠ
���^O� �-�>�k�6P��s��m%ۗ�5G�Ov��S���36�������$�Ϻ��A#�M�*��]]��۵��ə�
��V���-7F�݅^9?��D��Ă�g��`���%�I!4ӋrS��BD��o�L��mV�Yq�.E�NrW8D�r��՟L��{�9�N��n�l1q.�&�k���I+��m[��lg\�q<^{7�UF�����:j����H#duE��H�tw6q�Sb0����e�G��&^b�\����w���HP�F�o�(| ��7�&s}�(��o�F����F�!�IY���rl��Q��4;n�i�
Ǡ-���Q'%"����w�(��$��hi�B��;�Eq��	��^�N<�G�(J�Y�s/&���T~]���׫s	iw�U�]Ɇ�ʧ� ���ԩ.kh7�@