��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�G�'��"í�|�<D�\_����c�d�Asay���>�V ]Y+��=�"'�`}��Z�G5���H����.9�[ ��LZ�]�s/��a��}���mT���w[VRB��C������4/�E�^ZS''���QXV�v'q@Z0K��ٰY��>EL��}��f|�iN�����J�x7�9xYɯ�6�y�=ιG$
����q{����@Z�Vb$v�����EݴG�+����h�g�8>V��xq�����պa3F�v�_�j�S�6� �m�t\��R˾f��6�.d��*Z�x�ىx�!�Od<m~��E��;����1"���� *���-]mh1�n�t0�قdh^�>�o�5P~hm5���pw~<hn�Ͻ�PN(�cA�DTsOs�PX}1�Z\#rhLa�=P%�cU5�G��L�\��[;���W�L-�6g�`�`��D���dt�������-�>��)�����ɨ��1p���w��
e��?��� 6_�e��p���\�\�X�s�f��.�&Kuz��c^
��R�_p#q]\+�d�p�؎8�����+�3I��J
+�a2'���P|�(z.�4��+4�u��ֶԓy-dK*�UeT%�'�H�����'ƺ���Bꕁ(��Y�؍=Ǽ����hq�1�?���.��M$.�M� �� `]�����(v��8��2g���{��.��k�ӓ���{T_r��*�l��z]�cg_��"I�-����ȶ[���Y����sK��)]��O���h5�\�Qx���o��08,ݏ;��ǟb$���n���ʣ���*u��J�(�g�3}�Ms�hҎ,ph"nVA+�ߙ%�o���T)0=��tǰ�=�w4���
�	)�A/��N�_�&�8�lA�j�����t ��>51*dn���1�tw��$�ϱ3�n޸�'V/�������X�����i�čRHJ�U���]>idv���8�?ˤ�_-m��ɧ�W/�@�.��T5-�=s�B��K����˃0�kF����Q�,��[&�8�Bl)&�Wy�:.��D0~K���z��!˿�;�qQT6�{u�%.r��B�K�w7������r��S="H��� $�nV��4��z�T�џ����nmэ�CK�ˑ��Z�̗�������
c=�l�Z��M`��C=x��F؃A-�uF�Z�c[ս�D >�Z��PQ@(A���\5�`V�,�#7��Qg������胭�0�*-��[��:qW9�,g��4k/�8a���;\�bV%r��-��ݓGS�uq2��h�g���Vr�/�Oy�k�P���H��%F~e��C�4��]��_ &#��J���fj�0��˱5m`Ѯ�$Fh������Cn8���B���?�*y{��W�������c`S�چ�=}p"ݰ�.���yv���T� �
8��q-S���jA���> �)�F3���oo��K)c��b0]�^�F�9�yJѺ;�d<r�Xi+�q�C��r�e6���6��c-C!�q9���'�=ȸ}���m:ЉI����K��h����u7N��~��%{A�ق��r��z�'aY����������3l<sP.e$�X���\IiD��3bs�5៥���Db1���zX��ro;��&��լ�כ������Ka�j�:����v�J���8ֳ�5�t��.w��w�������ݔ�@�"�x�YWA�˝�g�����)��.������_Ӊ�^������ fi4@]��Ǥ�p�	�#��p�`\4�?O�U���э�	���������M	1�A�9`� �?7=G{�
	$�Vn!߃�����n
 %}���y�dԹ���E�5]n��=l��¥i)�f�f�'?���PE2�r���o�\��l��`�5n�rf���ܟ�2����ܯ�t-N�(b?�?���{]{��3E��,��Ts7�'-�qߢ�5�XJ1� 4�����p_���y+�Go�J�^�(�*��)v!d�5�&�Hv	H	g�Ouj�>��E;�*�ÄN�7�Ƭ	m�.]
��`ɂ4^ �RŁ�&�VJ��c�����*�Gh�ˍl��U��xQ+y�������FD�*B�ʭb�|�~�J~�ŷ��vk����v��H��1YḂq����w$������I��<^h���P_�ĭ��5��{��c�͏��Tf��{)�GsMC�m�N2x�:R�S"�����+�U�+ⷶ
r�'!z�Sq����䫵��Α�6>hx�ntr�%�p��{��Ȣ_D.��IX'�l�ÀΟP���08��%��X3e�Qi�1c�Hƭ0� �\��O�c���s^L�{���
e��N������k+R�͉�n��}&f]õA��R'�c�m�V��?=J��S}�+ F��+��ܒd��8q[=8hu�a����g]_�W,!gAgԵ;�l�A�|�1g.�B�/��X_��`+��U?��4���{k���g+�[�y=�%r��#2�3��S�EZ�yv�v7���N֏��"�kը�(��83�+����z�?�`�3��CQ�h;���=���:�^aW���ۨ����wZ��&;oy����R^A�x��h=W��=:���?1�4�\b��Yw��YH�}���* �)���� 3�Np:q1p
�9��'Ѭ�2k�	�p�Ͳ>�ſ=��oK�p"<��(��_S)b�2�c���fld������$Ֆ4�p�j�/*}�~���B��;�R�'W�M[�X�!�ND�*�9#�<
�v���?�_���Lh�/[;�	e�;^0�aq��_���$Q���7�)�pb�V1CI���}_�QB-�D)�͎�l�{�v��<1�ڬ1�2De;@��~d�D�$4&j��|��X_���	���A�~��>R�Ȋ���?��4
O�W�jt	{(�tl��,�a�!Vh"��"�s�^irZ	��3`����s��T�祐�貙2�m��j[jj@nq�N�.��`��k΃�3U���L|�uR�� ��"�AM7~֝�L�}��9�-=��pd}�4W �,e*t��@F�����"�����ܬ�2oN*)�O����1o���43�g"��>w���u-\ya��Xyb�zgc��;1����
[�����5c����W9�E�+Ѕ ��	�@�łǩ��!�-�v��򔊶ȠNѰ�t����v�����#��,��6z��
��p�{d\%yص����bZ䰐.9�lU�Yvhc��d�|�h~�Qd���B�#���FV�M�����QQ�O�ޏ|��̄mnQ,�g�,AY��(*!r�����ʹ_'a	|F@_ɨ�,6x����E��{y�Pa}TZUA��.�y^ �`�xq]��v\H5oZDD����:o2_����։�w��v֒DZ&y���Zy�B�V$W
�32ory����(A�6�xX�9��]��=������zؗ¼�Э��]�yM�ݔw5�*�=�~�N�"��q��[s��ʹ������Q�`Ƃ��ټǒ�m��<{>�^�}�-��TÄ$�x��н�8�_��UU @N{Vy���kע�@΀y	�k�~�ZӀ�n�����I�y�qm}���2�9�o��5�3�!S��V�`�����7�u$�IX'yA���@�y:F��8���qP�[|=F E��j���K�>���G��Vu��V�ї7OK����n�fY��uߵ
F�2Q�u���I���w,�n�)[�i��y~�>KC�k�;�6+&0��?A�{o.�P[�И���g�`�p����B�XC��g~".蠻���F敪�_�qM����J\��\�]����I��GVz�ш���D�d�t��9R�b<���C��X��c�9�)f�@�&~�\;��|�^�r�a,JX�'!�d۔�C�y�h�E�B$e�.���[]B2p��ܝ͋���u؂��H�j�<��]���V=�b�,3%�_U��)t���nHL��3�ɐ�s�O��X��СZ������D�
�Q�c�7��n��L��,^�3RM�[�e$z:|�(��r㚍�"I��-�N���� ch^��L���1�F%�m���l�N(��CV�E�>��zZz���
�gcB�H�僒Ak����w���Hv���@�:����팭a
��P¢m�(}���ꗢ�^KF9ʤZ�z`U}Z�F��IY���|���)�^�Q0ɿܼ1/æ\�e&Q�5�u-�@(�6�RM	�ɩ����ݦRL��g�1����o��E���B��4��wuX�*Ȫ�R���
Y:v����a0���:%BV:��@����=���.���0�?�kM����5��+�4��B�W2���X|!�u�OP�W��F'��>hB�e����{M����?�/��A��c���z���a/��!��%��j��q���e+�0w�)�>���V$�5�������E�l����	�0��
�]��R�R�r��k�3j���d�|�6Y9�~o>�xQ;�m�q">�|h{`d/)X�+v� ߻ҙ+�_���2�=P�b��O�spt����1����*�-U�+���o��ׇ=fe���*.t�̯|y��B��Z���y���a�[L�P�|�f�9�q��#�ܦ2��M�l����$�Rm?m�$�<Җ`�P� .ӵ�=w��]�_]��]��.���(O�f�l��F�\�u;u����gY�;:�&!�b�q{(tD�m� ��s�0�;���&�q�@}WܢrW���^�^�����=�uif��%q��=�2Y����m��̀x���(�\�S�;�F3�@+F2���8|��������_�j_����R� �h��'�&���2�ٕ��O�F�p���a/a���& �!��6�d�߲�Iw���`�0��:|S�⧛Tno���%�&��a��aQ��u��S��LJ0�3*L:5fg�Yb����W��*8�J���k�:�+^�nt��+=�2c$ eHn�Zu9%����1�𴭵����$� /W�.V	"�. #�9����Eғ z�M����R��-����9���d��4m��3���k=�n-���<�B>�)�D`s]�v�Cg,W���]	*��9w�g
I������ml����;����IR��������/�ec��{J�҇��}$�p�1&��Ȓ�dΒ�D�k�Ā.�L)?�=��%?�����\�v蹞����B�S��O@[��/%~4%c� �yXY�/@�P
*<��A�*�L0>:-���C��9{���A/�!�Lu�WABK��PV����u��OJ��)��knv��
�(";@�?�L�g�)��Uߓ�RLr^l�ZǼ����Tv��K�:��MAϒ�i�I��~���1�*ޭ�YS��If�q�u��T�q~w��B����a���
��r��W��d�h�B�观��pN��=�-3l���
��6�k��ُ�����2�n#Q<�3ڋ����&����/����(]�iN�� x`�A{��XxP��u��Ʉ��oq^���W�1ôA���}���[�Y� ���X~FW j�+��.A��+K�b9�G;�BXv9�-1;��D�'*:��I-���U:d�d���I�SsŸ�v�E!�f���֡�5B�Q~o�Ī�@��u�շWm��/ñ;�@#�ڶ��3���,���J�zG�Xр��H8s���$T����t 7�r��O��+(&,�p�
&��o4LOjۃi�(��r�N�%�Y��,����U��=�1�!��Y�4�ɠ$�$��RA	�=;��>Q�/{�byi&:�/�so��6ER�P�W+�it|23)3sO��"�M����eJ��G����`$�$�y9�뚠N���y�5�+��7^����d=:Ǧ�Q������7�\�h|�f�v�)�d�Ǫ���;���'�;��Y�͇"��x��Vp����4�VD��Am^v,��	X�a���tr����B�惋�~\"x�~�����Z�DF������;�X#�#��#j�;6t�v�֚�@�*��
���.�{��(م��v �i�s��9��%�5K���4[�3q	��I�6PF�c��
�3;aç?u0����e/�K1��y��X��L2�^\��+�^�|��1��^0�p�گ��֫%��Î��FH(�c�)��~n�B��P�Y�d��p$m%V�P&^h�A�Ʉ>�BzZr�ڍQE���̼)�����$JS�Em@w���fm�=b6�ۃ�)�>S>���W���¤��<I�BȰIC����1"p`�&�XM�i��D��V��%|BZC�<
x1�r�A�T{{c��7�&��ܭ�c&��>N~�� ��UMA��ǎ�/�n}����k�K�l]:�n�r� �.�4�~�7���-�����GC���#tk�̬����]y�\���<E%�z�Zp��� 6�X�ۘ�\�oR%�	��҅�l�ȧ��ܹ�7h��Zo����P`f�R�q���|g�{bt>�k���Ei�+��C6�s~�����`��Y.�[��������������|yƱ!�P�C��t|�Fq�Q����;�3!U���K�&#U=��Z <t�P���2�*��\'vUآ�D�n��^��Al��o$k�2���T�p�jۨ�K*ˉ�,=���ٹv���v������U-�lI>��e��Q���'[�MKA�9:���~�����#�����/&��3�e�˱Y��wc�'��5�PBbLd��ȇ����0�����,ɷL3�L�ɖ���Ύ+Oe��%�,]m�3���*��)� iw}��Ĵ)7��taE�"١ ��<��.(s���[�`'�v�w�S������7�h 29�. ��B?���V�9���<T�Ta���:��G�,�?�B^�iᲦ�N�F8g�䣪B��M��^?%C�B������ښ��=��L6��K rW8U��]d��)@�
s��g����YD��RL����J���q-�g���	"����|j;�D��[,>&��ID��-��RҢwjWtuY{4�r�e��A���i�u����8V��a�9��2�����~>�Y�oS�i��P��Gr��@��q�D���ʤ�������S��g+��t�h�/W��̹BUƿU;�"��;��&�M{u����v��t��9]x��"��������t�t�	%+�Z����WN,J�ĭ��2� s��j���|Ѐ�}��Vފs9�JO�#խ��<����2&�|.g���x��jԮ�ru��Q-�"b�(i1ԭ&��-˘�ƀ1���xe�Lَ\���P��62�ӫ'���R����'��B�h}�"���RT�4�@�㚎Ox�`f5�Ќ�ht�E�;]���s�P��4�&RT~��1�P9L��}�	�Q�B?�p+��Żz�l�%�&C�_
�P�w�����O��w�܂Ȟ��A\����m��b�Z,�˝Ug����p�r�R�()�)a;zN�w�&ۧ:!�;��%�(��T,���ڵ��cO�ચ;q�8�{\4F3E2��+���(q̲b1�`�:"����/N^��
� �����;ԓ��L=,���$���Cf05�T b��1i�wT�~�ϒhMsNe�]s\�n�0�[;�}h�ڝ G�k��q%p�2H��|���Tx�ʋJ��d%�ʭ^�M�"�V��ŷ��w��-\����a=���n��/����[<�?ѯ�6˘ ��I�q��,U$�VM�y�$h�A��-�΄K�o�]�� 5zC�dH�N����Bx���M*�M@������!o+v�����ηj�����o�G�/��`��Z�.�v�q�^9�%[�1�g���J:���i�n�u�	O� H�{��&>�c�~�W���5&cvo����:޽k�ȁ
n�*��w�cN���4���0�EE�]�F+j�������r0q�(J����_���B�̒nѵy_3�A��r��s\����A��D�m��d����82�TQ�!��]����j�r��G���[`�1!���_
|�7Vɍ:�a6A����ǰ#أ�2����6�X��Z=�%�0�L|�!&B