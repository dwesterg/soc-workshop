��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��� W�{.��h�ג^m�JK���T!��e�5r�`3���h�?8�:���y���7���
Gs�fb���0�w��t��w�v�R�ŏ�DM�&8�&�8�|����՚L�-���y�7�S���m6fݡo����@��Mӊ����%��lh�n�&:���zH��(�����O�.�SX�Ε�ʀ_�f�V�z��Z�@^���X����5 S7�@H�w%y������2���,��u��V�kh�9���������[bS���L�d�S��ž-�V��Cc��=g�K[�Q�sM̮�A�]I}��X��"jօ���oO-�?8t������'��p%��zc�m:���W�ұ���b��F!�,��a�Ш�RK�C�������n��lR���vF
��Ŷ�^�UF���-�����%�p�v@;3�]�.��f�'�eI�Z(���^�4���!¹^l	G�`������\��=���L�өI���M�\� z����@�CY�رH�n,#З'Jd��0F�t�G�-G��a!kyQ��4�Ҁț�W�QSs���hQb�*���5���:YP鬏#�}Dje�Eq�p�po��,w�%�~Ћ�!����d�3��>��?�ZG��(���(�C`o�o
��@-]�ƤU�a��Vy�:&de#�=�; e���-@Bk��S��R�*7?�D���/�~zg]B�MH��⑙;��r�h ��3�(��Kg����!�������2yB£`����CU�9H�`Φ��6
w6���bj1x�o،��]�Fڨ�ҝ�-{rw��������v�C� �B|A�D����2�4�k�	W��R\
�!V�E��X�;�.�\�rPJ�JqKq��y�䭈��T�&��G}��pT���H�/ܧC�$�8YU�>9��Y�e��g����"�YΙ�ǟ2$�z�|
9i����_��Kz�ƬJ���i�d�Wd ,����`�L�Ͱ)"��"Z��{�}伫�'V�'�!��y';��Et��d��,�u��Y����冏��P��ڬ� ~�P-��b�F?4��t�:f�SZ��x�_���7�i��XY6�Du��Ԡp���Al	��v�>O�$�{=l��"���M�k�n�ɲjm�c7�v���#�ٿ$�R�����'�x)<��[�
�e�sc�QQg�&�+�?�om��������o���k4��y`2��*"K�[+�l؈��6�QA�K�'xb�2I<]p���
(�F���eb��q���K�H���.�q�@.��+5��1�i�W"[���*��\K(��H
��l��#@��~k��_gɹ�ӿ��o�t%Q�Wx4ZEY�\P�~��-*V�<��/�V����ʺ�L#(�śJC�I����)�Ē�S=�v����Ҕ&�U�%����~t�෿o[
��Ȼ.����s��%�t�;]���g�Ys��
p�u���B鍂/�Il/�c�rko��g���'C��3O��u���_���H~�v�@r%������b���j�@�����)4BR�����;�-B��pDZ�' F%���~���%x�cn4�/S�o�|jT4��*��g����?���b�$�p3 ~�x���qa涓,5��L��h/P~�o�qV��g�A�$�.�S@�j�����٭q\O�R��J_�&)���0���H�� ��[�%�Ns��/_�DROj�64J�F:��2�XL����9t�gՍ�R��4��(�^/��S]kTht�wސ�?i�n
z仓b���[l�+ӠZj!��=Y�0�����[���EY=p+M��oz�7ɻ��J>\��m�!o�Z�O�Y�����/]���7�HW���'[2�L�ӥ9�K�:�1��ܤ0v1hx^� �(BT���	�;����@�;j��e(���M�-]�'����U�# |��<J߂&M�k���o{c��PֲJ�F�*���M�#�b��U[��#��
@m�_�o�dCb��-�V��F%�����s�݃�$���Sΰ�QU��B��MH�u��z���e�s�����3l[��?��$t$�x�9LHɆ��}��ꩁz%lt����K��/>�;���5�cӦ�������:�b�T�7��U��;�Wu����AΕ��� �h�V�W���}Al��Co�?�r�V�0M�dÕS��[{#JԲD��yz��ux*;LC�&�U��D�I[�K�X�A��.�&�B+��"��� ��h�h1�)$�0��ޓ�a �1����r���&��e�I̢Ӥ ;g&m��p�&@�˛�A���%�0�wA�ki; �W4�G�oٛ� �xP/zy�N�9j�%�ʥp�p��g2$�a�&%�t�xpb�I/e�� �$�h�2#g�ZJ>�i��4��B5�Ö�
n�aTU��w��'��ч�J��'X��F�w���8���Lee3���.,K(�M2qߵb�����Y�a.q���fB4R����n?�{s����Q :HF��؇��V p��Ku�<��K@�I�i:9R�(��T$j�B�na<)�f{/�6!DV{' ��i)��^�3�_w#?F�6�WZ�D���,��_
�_�	(�
��$ZQ|J��!(�3�y�������m ��C���;a�����"���T �d�G�Lr+�<i��K�������E�
"��j�+�$��u�p��j�!ɠge>s�sdr��� R0�ɡ:N��z�:�3x���<�W���!O$����,vs|��D��q��z��'RZ�i���G�5L�0�Fy�":����A�wԔ���9�kvbsXᓒR3��\
R��~�ߡ�����B�����)%���29b�
QJb�;���+��g��,��z�Ma��x6���W�r|M�gnTR��6��F�#�%���<����1`�U�!�6�@[��R~[����r�Z�;A^W�gJ�SP% ��6�� ɞ* �n�Ԡ(R�F� \������K'����� �W:�F��B���\"�}{�߳Jc�y�ځ{�w��)^2OE�BV
N��N���q���������
�Z����zk�]*�9co������BKY��ɒ�4/��2��)X�Sy����.գh���B�'K�sq��Z���ۥY���嘆�k+"w��|�M/�6�s�P��M�Sd(,��$��^�B�u;�_*"��{�5�����Ih�P}	+S:���g^~$��w����.k�a���֚7Toc��S�؟�>H7t���5�n�P���6M{�B�]=[�9Z�^�E���	�Rs���� �^_�t݊,�P�fȄ��1�W\z��r"AB���v�c^H�Fͦ��_�T+A�O�Į��{�P��rD����iR�)���Q~L�Gm>���Z��mY�6|�oҙ;z�`����/LZ���9�铤�
����g��>:^�8���m�,�9V��Q�,���V����v���|�"R\��d��*)7�l!��)a���9��y�I(� �zf��	ɮ}�1���(�m���Ŵ�
,q��w��Ž	�������!�kL)�Lft:鰒@�D����}�۝��+�>�EF�����o2�	'�jfsϵ+z�g�`�	4q�B���~�tw{�E��������֥�y3n%�ᙶ/Y;�\�7�jhk�����H��n�u0���ȼ& �e�^�����k(b��q�/s��N�!Q�zi(��l� B�i+�pn]`��*�F��W_�������JJ��{�i�ŉ��p� ���	�NN���bo*��KO:_�b�@Q�N����3�������z�&����/_�#4r�W2�J�u�Je>�y�K��^���ċm���XB��x���t���6�7�C������RZ.ּ�׈(�^{l�M�哩�a[��"��j�-��b,���-��O�5!���'�e�����i���/����hrxt��_�,,�=�[��^:V��Y~��G?�
�Zla�/4\����}a�����ĝbBwl��p�^p{L�l1�F�7|mc����+�ly]&dGn*D�ۻn?��Ѝ gAF'�w�q5���L]�l���~	"�"{p�r��F�؊
�������h@�s�<�,찟��F��ܿ����X����tf�;I���4�]��i�^5�_0��)��o����-�#�٪�g��d@�'��
`��?z�^
|՝�l�k4��@��Tp�
�)�	$�X�@i+��X*�4*��|̞��ri��N/��}�7PQWuμ��l��T5�g��4%C��W~��ݣ!8+9V�5����c<Ll2q`���W`������	:>$=�Bpps��Yr�~�D!}^hx�j�|2�r��Q&�xHq��u�iK���ۆz�
M�WܗO9Pv~�p���������)Q������U�ɖ8D
av��G�R.5��	;K\��/�7,���z���[����ek�m)=D�%��I�]r�fOB	#7��w EK�=�k�Y��Uq���cb	�iy�<�L�rW�w���*/3[k����P*�T�Y��k������Fܖu`�[s�Ԭ�x5� Y�%�)F�;Z\=�q6�>љ*}ߙ�.�̎���^��x5����[�+4)y�%B)�t�v��B|9�g�d*֡����X���&fHp8�[�I� .�(��w�#��JFT A|ҕ�?����+E�N}�;*����Tw��|��� 0��N�e�*-�n�E����=�w�Às�E�I˄P+:& ��q|ȁ�lhP����%���1��Wg,��^@����05[O�sW�ϟ>��*f�0Ϋ��t�4Nc�v� ����¡?\��gk{7W��o,�B M"���8u���b�X�Z=��sg�/K�N6P����|��dB���Ir��ÚOP4��T�C�{Zv��e���ffc㤁�,<`�=�|T����5�JD�7i_��Jґ�LqR"/����:e�Jr�I��}U�&C���L�)����'�qΤ��Y��#5b:ɑ�H!QW�{�ыL����e^��h���H�F#��7��l�U�=�a��V����7�-Cg�`�0����V�F�o���Z��+��%��X�8�7R�`��?��i���J�7c
-���0��=R��R���?p�T��)؛Y�y��7vx���I�"F����o�,u�R[�EG{��L��֍<�Qi����
��mnΝ�>�^(5���iǒ_���7όXk�i|��]���#���5?��T>�nP�k3��,7�8��Ġ�w���!�8W��b�ʫ�4;p3PJHF]sQ���RR;����Z��|<VJ/"�o[�1�����b�ƥ�ۺ�P5@$����VtoR����YH�#vo�|�O��Ǐ���y|�N3�G[�<҆z'�~o�l�$�d� X�?���M��Wj�n�pZ7/�n-.1�N:��K�з�R8����Ṋ��E�}���H-BE�,���m�j��ǂ��]��f�\j����7�8���1��dzaP�Zh��gY��1��$.�D���R�o���@���
��u�}���������s���Qj��mγ���"V��FR�mƺ<F)��5���S���݈����� �BKù_�ն�;��<�0��x�p׺龅џ�p)
o�ӡR3�o�����4x�%v�/W��J���ϋ^��^J���͡��S��H �#!�\�����+�W11h�h\MQ\���_��Ta+�Ct9�<��WHJ�uи��T���w�u��S��������i#_�N����Fi��E�>ٺ�#*�K���*�&��a�𜙁�,���$kYvl~����aQ(ɿ�<�w���� CSذ��r���)R����l���4�N�L;
�!�f���H����u�&P��4jQyFE-�j*��%$/������{��f �0��bAVJ�މ�%,o�UZ�%zt&�s��'%҉JM��#��Y�8Q�p�Q�E�]�@!�U���o��Ǭ�׵Ҟ����(�lg_�7I��WQ��i�f�7�l��B��ѥ��g��:��M���&#�����mY./Pܕ�t0:E�xE���cn�co/�Y51S3b��G���=���h'��h��w�������N'��N:tӖԍj�%g�D2�^��c�h�P�ږ�{��"R��U]�4�W���*�+�;z��W<���vW{G���F8��i`pT��C�%fiL�a�<���/�;��ƚX��-"��70\Yu�l�D��i�P$H��ĩ���EXY�>��9�+H=��;K�Y�[N'y�X����S�� �3���(%<�Ǫ�(q��{3���~R}ޫ�N JW]Pt�s�h���X� ����k�)���C��oZsEh��_���D_qq��'��jF&���g$=���УQU�M�� w�!k�,�l��)��l����N�i���;_1����g_��H;U���,e��[��e�ט�%���Z��P�{O�a\�/� �8,r\D��/h�H{N��$�J%,��mk_Z�H
�w7 L����b\��e����7R�?"�G�A����B���z9'�>Ѵ�"�6�#�&��h�
�ȹG��{��9�A��^& �{�Ŷ�p-�=|ԛ�rp@i�v��f��a�a���6S5W�-hS����Rr-�y)��5��	��#B�z;�R�j�����Eep}�<DpY���l��HF[�[�-���ҝѨ�ٕL�y
�ǰA�C㢨R�zK۵?6V�Nۿ�0$څI.����ՙLS�pYC�a�1�D'�~ʐ����v��w���q���I��؏R���#l�e�`�!c����l&���G<���܈���J���<M Qp�j�,�_��>M'p�z���3W�=������I@��G/�`�w쳭�ƫ�.��Lq��~6&�D3n�Ū�!��4`EC������n@����'�9..>���O�Wu���;u���Ȫj���0�eNJ�����*��/�������u<��x��n��@B�>>�A)����Í/���8�� :��_ң�!��x��S��#dBi]F��]�������\L$�ծ�R/��_�V\�/��5=k��N,��z�$	���~t�%�N��e�6�vx5���C�T�?Ӑ'6j�WX��Y�P���1Ώ��pa'~���3w^`a�+�~���K���g�H��-��4�NEbxi���zt��,Z�6��c QT°�w��Ŧ�G�G��ܐ����һ�զ��*�Ub�x�_�Kq跛�қR�oJ^F�ُ��Y�P�����-ı3��Ȳ�EjR�%aK��_�T,_a��1E/�����ow2&W���5�;��cjVKp�����ٿ��e�
�9�e�z���7�5��-W��.�B�
5�֋�|�}�El�3�m�e�fˈj�;�m,��N�te�q�T�J	qi	���8���O!ч{�w�
�Q��ѷ>�Ŀ������h2w"��~�C@:U�\Q쁉X!�WQ�IM��r
A6�&�먡�����SW��y�K܅��F��:��x��V��n��d�g�ٶ9�HI��e�.M;1.����|�띔i5�{�2����_�(t<�4�F���jq�b�-V�Ӎ7lo�������/r��~��?AO�g�w_���|h1��!88l;��n�}��Be���y��t�Bv��MR���F�ob�W�?LƘ�C��r�\�z:w���
V]��#x�l!m�㧩�9]��[F�y0���0;��-B�v�@�ZU��"�t+;��$�ؾ��y�i�a�蠤w�U����&�����	f�8��>Y����1�����O�����Д35�����v�y�#���"Z/�ꎰel�jy�n��Ӗ������a���%��&`T�'h�Wg��ty���.�I��ڦx��6�Q'�|��Z<��qt�s�>�n[}w	Y*=Ny�/^��=�.�u@ ~փ�����w�R`Z������ �˞��;����>�4]����8���;�o�[�U�}�� � �7��"��<�7���ʆW�MM�R��"2�gc������=p��,���J�Hz���d��|kL=茢vq']^+���,���<�4Q	s��vX��{�.���F`|�R���I��}q�MS.OS���(^�Ք���_���v�W`�˂e�#��@7��Ԉx�IE�l���Cw�
wP�&~�9��v��788"~��Ś�f�-�o�������?�H�,��ONҖvh�4��W�x)�l#Tw�J.{�>jsCy�fQ��i\Go�ݧ17i#��EpG:���b<Q4�o�$$���K\p܆jT[<��n�%c�6P�走����ˍ-����$>A�����L�����eZ���k&V��~3�Xb�]�EcC��X��U\�7���t,��n/�e��
�6��I�����%8���YY�&���j=�+r5H��k�gT8��2��]��s@��kVBK0�#֑�Q��z)��)r}d.*�?����^(��llK��ٯ/�G�(�A�xU���͆������8k�^S���$)3��YL籈
��*_W9����:+��O킓�<����e�a�|/wC�)�ק������-���Gs��a�J5�JR������رQ�J��:�)�EF}�����Z��pX��,����۴��Ak���>,߯��j�Q�ΪM��H�Tˎw$%��H��nP��z��͛�-)�nՔs9��=����Rڙ�F�`c� )�YgG���������!��in(/00�Cd�9�N�j��9wob�ut����՜L���Hs�Cρ��Aa~pʋ ��#��U �Ӽ��+�2��i���`�U�~gJ֑e�X�������z��D�$H��hU�t�|�X�ʂD/_��@v��F�kMp�$�G0�C��Ӆ�Y*4o�8\�wj�Y�M�	Ye�9��rآN� �^��@�X���ap�����g�% �R���:��蒚S�'�.�5��b��Jm��������mB6������團g���cji�!#�����ͨ�А���5ʥ#�C?4t���H����ɘo���f��r����;$�E����HW�}_ݼ�5�"1�>��&Ta%v�3�L�\��fY6�|÷n�����نF�N��[�ѧLO9�"��ӻ�Ɵ�n88!��4S��4�4��UR|�mEA�'��O��&��j[�8��
��'v+ȍց��h��j"q<֎'}J�����\�)����E����MuHb�'_�c6��%��L��]��G���Ό�H��3P<���؝r���}��L�_� ��B0t�y�Vߋ1�$���u-+xԼW}9�X���E`��(����A���7���|N�.��7l}�R��p����'d��Į���[춼T!$���M#+�%�M泦���r9Vl���({����XG���G��$�u?�(Ί!KO�I ~v2Xp�)�bb�8�>�<�y�(r�ּ�s^{��_��n�i�m�TS���e�P��qH�	nʅx����L���k��H<�Bw_��jLWN~����C�%�$��I��!ڧJ�%���@U�.�&Į�o&�������De)rY]cG���9������j�QL�!gݠ��ą=R@�xh�)�]�3���o����Q!�� v���tKl6����Ê��L��W����<f�i%�}�T���ȒZ%�卛�i��+gr�DH���7��DE.�#�m$���P9I�˘)�,�V�v���.�C5&��������"�{թ���`$���_�P�HXd����ެ���HH�٨� ��*��u\��'���g�=��G��~̙�-Z�B�!�%�-zh�
���I�l�#��Vd>&V9��:y��g�y�q�s�ǘ���0�n�ƍ���p&
��!-3��@U���}I��9�TdWS�b�[��3b\3�;z.���{�>����P�j,ƥ���-I���$"t���`�0dD������Z�]�G�WR��F�M̔��������t)�C�'�p�@ 9���ʰ|���D|Ϊ�'���9�G���7���r�֯/%ʎ=�P(O"�����ϱt���(�S�@�����dlY����h��uA�w��z����+\B�Za�e�.7}u"��Q�O����P�L<e���Q����K~��߫�w@����kS�]�)�����wS��菠c��QH��F����}c��$p�����g��̩|%ee�dL<.��qU�Υ�C��qqt\|�w��3�j�Y[�}O|T�ף���H�����ʣ'Q]>�Hf��v ���.��;�dL��l�*hM� �4�Pү��u��yp:���3�\�֩�UI�>�_>
u��J��X�R��V�Q Z�\����;d��o[߭��H��'P�� ��@
�?�DCo�|���P	��$���JTB�s�et,�s���_��4[�
_M� �QQ]3����wFhLԠ��� �g��x��isx�g��4��
���A��9�߂�u�Y����;������'8G�����Q�ƞ�9��cs֦�������
����m:�C��}I����/�M"���u�d|ӓHq�7R)<k9���V�$��4Z_B�Knh>���b��A���4W�n1l�P�Fd�N��Vgl�f���ա�~ɉ95Z����Ӛb:���8���j��Գ�M��Q��2�:��]
#�s`ߞ�j~(2����6��׽�]��6�׽+����N*me\^�����#�
��"8�	_�?Dm���-@zG���7C�y�>w@v�R}!��16B����S��gn̰����zC��e4hW��*�Q��G��/�u��.�Ξ҂�_A�3�B��MÄ�*�5w0�/�o�:5���+@�MeFX�$