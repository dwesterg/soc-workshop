��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+tu�[tog9��ް�Y�ۇ��I@���eUF�Pw���&�KBBq�R�	Y&<kVsh��c���Rk
7�I�1m;ʨ'��ܮ`����c�TYl��D�a�#�+�D-�,��X�b�CV����3��}CA�h���r�}Kp�W%��v�O 0�}OE�!���Q�CjE�K[��|�%ÏUH�㛇
	����}+��.G��=5ȸ�������fmU��Ԭ�"W*:<��_`DVb�e��_���}�S�pX�jS⁙>�rU]5o�y#8W�A��b�{l�
�
vu�Ezǩ8�d8��(����'lX@}����ܜ�ʍ�&�m����OB�����֠��C��fS�:�C)0�&�f��|k�����LY�J�h-?�⤰�?�T�\_���7�g[�}�f��6T�إ�k�����<�.t_0������r��>��0��ἶq���sڷ�'C빃|m��j};�X��|�X�K�J�Bum�Zh���p��_��dܻr�5��[>�ߨ�������˓�6����p>�pשS�����c��l�H��`Řׂ"ϗ*`@���RȚ����_�yY30N`��2-0�(V���F�|����]\(����g&�ku�f�Ԏ�қ-�Ԕ��B}=�ʂ��8D*�N��w\��R<t�ʘͬ*�g�`�9����J@�V���������"���2R��n��D��m��$D㝄P�W�U�G{�;��̒lҎk���8ݫ�0��x�W�BDz�f\V��B�1>��/(�����͉�' Q�ha� �X�OQ��8��de��8��d�y�hj�U�hl�����JB�ߡ������ǘ"KdhM7mZ;J�g�*�ǟ�7Τ�� ���`xa�m�o/O\p�h�LB����50�4�3Dz#����Ѩ�TJaQz��P�����Ma���m� b�����D����\,�=�p�J)��L�Fq��$�:�~+�<t�!�Џ%ĸrCOV�y#�z�h����Y"� �
��rvK���Ϊ���Gz��f�u�r�=����F��nC!f;a!��a�x����6ٰ3e���c�f�zd�b�
ń��uU��U:�|*F�j��X�)��hO)O$u�&c��7�lS�E4�(�-�i�����ymO���H�
�C� V �䂏�Cur��K&����e�������!z�]т��VC�$�{ќ�L�Bq����i=/�ۺ?]�cҌ>���L�{?l�!��_�����3�#����-�}.��i��(��H�N����9����D�����ů�0�d�M2�� u��`�������OBw�� �JS��ƍY�j�|:�Xqp'�-���%�g�M�-ɯy7�6�;���{N��E�T���I�+�s�å��8�(B74#r�e6q*�w���@�qY�|�ݹ��5���]�`�g�LsÍ B��O�|l8����P�E�N�ŋ�v�Q��"j���U5��ң�}ޅ�qÓ�p�d9��v.ͷ��v���1�&.Ѥ^��{b��΄�m�d�EܩN��\)�M>"m͵�.t��6n����V6�|e�t
}α�"�i���I�y� ��A�"��=��ty�)��%���Žy������կ��A}�Z�6�������Au������+��O�!W���	��~y���%	���X��{:��2�'S�k���ѶO��F;���S�a�*�����-�' �4�AJ��h2ͯh�hɌ\�a`؁
[����p�H�Ȋ��r�r�����z?�� �B|���g[Yb;Z�q����n�<M��Ttr����zlK�J�ȣ���ޟ)���U�,��%pVRО�	R��#ڎ�Q�vt0�^��\;�N�r��\e��3���AZ����W������##+��/١�f#�oC��y�3�ۆ���k�LYk��$�;�-Q���ظ���T���[���	c�F����a�/�\��z���V����g(���ሮe��oڤmwB,h
4���~��[3�n0ҝǆ����t���t��%�#���c�Zwg��芯^KN�R��:J՝��c��=	IL�I&��9q��+�G�Py;umh�l��f��a��j���1��v_0*�� ~��qGeUx���\��I�䓩=���C#ǅ����<-�����S��F��#��	����
*���<�,���]�+��� fg��rq�bf%)`ٚ�݉���~�.�7U�},�0x�(/�E�*U�F�g��X��%M��28� ���A�h,��J?%3�gU\�|I9�0~�\�؞����޸�ڄ+z����X΄v\dBm�L��h�yv#�nAd�u��f�n�.��-��k�n�uO�$ZB�4"D�%�X#�)u#F?d���h@e�v���E�14�x+;qG�G�GR��B�)@7�?.o���Nv�������Î�w�yG����]�G(�����`�p�|�3E����J���xv����#c��w��N����)�Cf�釦��%�Ժl�o��A��bB��g����VԈݥ��VB&8:7��)�\x�+&�	�aI�adE���$R� �h$�ϵ@��v�Q�$��[�Ҷ3sC5S˄�h$���b��%���n�X�~Pz�}(����{;7�t�>��O�8t�4�G��D��w�~D?k��JN���Y=�O�XS�luh�D�HJp�#C	!�&t8�	���Ji�y�m����<k�<�O�
��`Φ�\��$������	,�NP )��w���>$+3n�{��d�P#�im�O4�5�p�����r.i��\I,����3��v����j8�ȲVD]����η�L=t�鹓%����+EU�뜘�r�~L��~)y���bn����ܖ��L��C� S���P[���n��ʶT@tg:��R�4��rQ&�}��o��g�	��b�Rx�F`��Y�q�- ��@���8Pz�xSFg�]i2�dJ��������)�����_R|�����(e;C���?�o�����Ġͩ_�d��d�n�R �r݁p2S]V��Y�nS�?|qh���oF57CE\w��Hm��+
E�D}���3f���t��y��4�<�r��Sd��3�-Bz�O3��𕎖=id���j��X��GCG|�;Zu�Us�c�"������o������yʮ��!]����9�}�ˣH�D��	9��ޖ��v����ּCND ���rW⟪�xA,l�P����-HQx�sL��a���/d�3�OF��r|n�)6sPa�E�jA���%��P
eȞd���B@���nO�S�pz���"B�l�?�� �����=
�[sf�@W���k�t�x{��0�X[@$�M��r7�XiB�괨�q=G�w�R���j��.����_Z�C�Aڭ���C(�'=�ٹ����L�a;��eO�����f���!x#c�Ү��~P�I�6�Ͷ�w k@^��4P�1K@�F;�1]���3��baW�����/|��\vp)`T������|)������4!3���E�x��F���9a�ic	p�F�A��(�y��:ፈUO�O�./]|)�R#�u�������QO�uQ�UJw_XooUh���V�.����h��PG&��G������j3���t�-�)�	y�ĸ�=n��!�12��
���_M兖�.g/Z�yW��Qxs��g�'Ȯ���iL�-�@Az��(Z޾)k@0�Qp�oW��q������[����3e�Q��W&Gƨg�g��C�:�p!"8vQdGqj�*�)��
��!��"�gߦ��j�^�KD�E��