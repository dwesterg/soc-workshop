��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���ORagowG�C����o�[�����r��`�.:�+��R^H��b��uꏌ�A�+n�D���S(�ӟxDM=����:6z�&�r���A�l�Ұ,;�p��2
����@���ٞp�E㝀D0����L��A	�vT`'�ws�r[h4���
�c�;�r�b�L�V>�=��睛bA��!���W?�G��	�o�W֋5�Iz����e?�뤡'�Kyv���ZLF�z]��7�n�[';��OV�n_P���xřׂ��A��~rV�O�Z�{�]�i�?���Z�Y��=��£^r��J�F:X�I��_G�ɡ�.f�
���"M>ѡ͚�	�b�h�=&Р<i�]x)�����>�w��=	�IC�@��Q��&.��{�f$T��rg#�߰�xpN��s&��Ǟ
���0�X��ͱ ,K�<���Z�0c�iaB�A ����Oz|���ˑ
�5���|�n��f��� bp�V��[E4������;��!��ۛ�07�|��@��d��cإ|��%�^�Yc= /�]�,AƢ�Ж�w���l;hL�M֖�K��� �K=���pd#� �6W`

:_֯�Y�]���e�sW%�V�e�����h�����j�� 0���	Slcd8h��Z�#ϕ�D=�6Vm{��B�g�!�7��%u6�:
�I�~���QF-�y:����ǫ$5pE6w�g=C��X*p�bY.���ci�ม��;�ifӄ���^��;�s=�u��cڿ���d���*��J��v/^���ގب8n&�t�S�S�P�Pڭ�2����� ���O2K���o:i��@5�0ĵ��8���q��}�N#��sU ���_�=��(G�/�1?_&nRl|�L��-L���^�p���#r�$�!�$+q��	$�P��߲�v�*HTȱ�������T��G��������pL�_
1�aȽ/ ���ʕŶ�/�]
B^~�d�2� �f�!l�5�~�J8��|w,=d#��NN�p��Xd��>3��C����d��d����w�j�[���� ]���	���"�G�2/��@��^ȑ�rp�,nc_�����}��4)��/���P����n[r�T����	@�S�vÊ��sM���	�e�P98�/am�'B))P����ҙ����7��)�4v�>���a�t���f���:IE���+0��GlK �bu��ʘ�GB��>���J�_��i�%���:&�4'RW�}��>W�����.�����g��"���Ѿ���乪����j��4:���o\�H�#�t�����/�|������N����i��ms��9�s�N�cW'��4?�r�o˅�;�.?Q��{'�)}�*�Ӕ��X��6�!��a��:��^�H%咔�e�0^Ϩ���3��:ѹ������%����pi�a�eN�MT�H��o�L�߲� w	L�F�<����ׅ��6J�,��-��2����]3��6V�s�e}7>ޛ���~��d�/3}�Y(�[�<�� "S3KICqmD��`Y�zNό�D=��ixH����5�E�
1D��� 9D^��U^,ǋ ş�i��H� ~O�һ�N��ڝ��QC���P;Eѯ��I�$�>��:Or�Κ
�P��4|��k��⪨��ѭj3����SI�VQ?��;��7]�v������U�}B�ϱSǄ
dGQ���T.�E*a�����k�;�W�Y���}�Qn��d�����d��������Zƚ�0DA���*�NB�d�J��@ �v�Ho��$�c��������<����V�"�h4X�~��Z�
�����wN/��)���HxkИ�h �d���G*F@[+D�ޜq����f�	j��$���0�
`�[wOc�4�mc� 6���*;��񝋎;E*�m�M�V�y�+:�����8@M:�#<�*q�v��ot*$�L����g@ɷRBlM�9�ޖz��p�md�Ǡ��Ep�=�H�ή����&�Kf��:z{!%�xՀd��XG2�v%@��n�?�l[o���q�Jнz҃�`��z�X
+Ġ��*�͠zĜ�y���7�P'��G�gR�ք�ѐ���[(�h�������ŷ���o�Z�?~2	�&�͏��\h���}R���N�!_<���7�W�߬j���{�����p���'W�^Z��><�ZC�x���tiQ	v�xԅ�f�����
/E$�س���WA[��ew������,Hb^�l&�X/�2�AjI��ņ�vIQ�s|�۩xZ�ˆQ�����]8����:_m[Ikd�׏oȊ��^�u.�q��nJ�i��NW&.A�7.�ǽ��ș�Ц��FqR��l!O��V1����Ҵ�8S(:	�6�O�횉��H��QI%��L���8�#��G#O.�c����$��-�	�7��&��m��X+���@�=�Z��w[KM�C�0���_w�lB��~�]��{$S.���ͯ���-=�?�֧&�Z�cm�[@X4��J���C����/愞�R؝]'����(+�ͳgR�r)������3��L P5�� �$�c����! 0j>�?aXS�0�ك��|��z2�b퐨�)cٗ���ΰϪ��JAU���_�� ���7	8��{Ag�U�a�y�o���C����=TجX���I�Y7Rd{�'��?_u���mLW�\>[|����b�#�^��iX�(��4|nk�i�Ήԝ��M�J?�i�1�h��.Xv�ѯ�|s�}1�Ԣ�Zj��ś6�ݠ��cY�}T�s�$����+H��;c����kq�8���avP��܏�d?b�����1������A;q�wO�<z42dܭ��#e�Ӻ����+[C��zT��c�U�����E���S�N�0���6�w����Ǽ�zEK�yF=���u��C>�7p���y��6�N���R�E{Y3V���eP�ύ�h����~Æ\S���Le�7����� PX.K���q5�ލTᕐ`O�I����~�->���d�3�͏a�bZ�زI��h�]5ܠ��5m�!f�JjZ(x/^݀�dxfNF����׏
8�C��R��(Y���/_1����N;r�{WF�^}�e�׶x����Y�<1���M��@�n]����C��9���
��BP;~vX�`0˄Z2�����L��Zq��_5QW���HE�]������?�n���Q���!;�<�*�k�� ��{P��4x�5gbAe��6�$�&,l�j$A�V5�ҋs�2�߈2{-t�"1�xE�,V�w���
4��r �-����
�D6�ս�Ɵb#|���Ԗ��~���S͑�[��0o�򞱳_^���>�n�<M��fH �ϊ�;�����8� <��-� �K�i�s������Vp��s�|99�� yv{]6y��ەB�{t���ԋ���*F,U.<�r��RޕZ�h�l�T�Y ���	���]���ͥ �	?]����2�=Q샙���\n{׶�x��Q��f���Ş^�נ'�R-ͩ� ��c�$�$�*�"�K���Qʢ�6d�v0	���D�K�ۼ�g�C����Nb�YcM �g�sx�jЄ�톧Q&�$�o��p}	�d�,Y�:����/��@�j�Z~�W;�-<�D6��+�%4�/-)�ߣV�u�k�M��^#�S��fmo��=6�"��ԣ���N������ ��V ��V���q�^����xA�Y�k�$^:���s�v��M��I;L��Z��L�sϐ���	�b�|њ�,���"K}<�]�%[���S�b��R�n�$�o��1Ϩ|_aJ�9����-���.�Il�}��±��;^B�tӷ&ԉ��?���a�tɷ�����m��xV#��!����໇��g�!��`F���8��H���O��ܣ��g�=�ɋ���pI�Ӈ�����Sx/��d�W�#s�?��e��9��9�TҪ�L���~a�6	����`z�L.٫�,6'ZN1@�r'@7K���$��H	�P5��+� %�b��A!i�H�[���6ɯ�d��dm_����
���k��7�e�G$��V�7��+�n̘�Ӆբv�H�w��b�4��]��B_BT�\H��ujR��=Ss����Q�|�tGIoW���b�C����V�p�Dm��+���u���#��e�֍4P�g+,��3I�K�� ��S+!�j�IYK���O��z�)6��X�i�P��թ���תkK�-���~dh� ����p��b�cjã��?�f�W
}`/��Dd���@����03�d�AF����>�����^�HEU!��9����:�Y4����ȃ��o�uh�8�!��tVtry�����hT D[�ME�+����v�ӗ}+zNAlz�O��`�O^�VI��wD���jh����З�NVɣ����N-J�=R�˘����?�����hF�;䇤�s��A���Es��|
�p�.��X����(s<-ߟ$`��re*��=��D~���C�z���t��}E\H+)�4��W
��s��#:=Vng�;�K�Ê{����vf�P���N�n<&��AMYZ���2ÀY,���?�:�;�x�/#Qaa�9����Ə*�?��P�<�'К$"aq����5�"O��ç�%A��[��p6�~�?r����j��&�q�f�+�����&�]��2��q�aU_Y0�E�U�� ����]�u&|%NM6��-�A�X \ :���t���3�tR�~�l�\���]NlF��`�W迫JFP� �Tf��}����C�%ݟh�=�R=��Y�Iג�*�H�������b�( C�;`�i[�4���E;l�[S2j��
TٯD[����R���Ƶ�4���,�N3o������C�!UM^p$V,h��F:`��F�!>���O����z2?Z��q|b��$��'���2v3`����v{���q�*ilJƊ������-ڷ��Mƫ�\��_"�� [�q�f�6�=P��@�y>W��X}��<���18���R�ٗ-�RK��$a�L4r*W�vs6מ��N` w�T�[ZW
����� A�F�����׶�q�A^
ڽ�j�w�9��[Q4�75��a�	i��"#�=�?�w�8j'��>h��4�B���z��d�"n0���>E�}�ۖ�nv���.�t9��@��>2ꟷ�-1x_��Z�+���[�dYӗј�Y���,�u%o�s����fVjԘq�;	����k~#�H��I	����@'G��\�o�-%�~�e*2�;�Tr��H��H[�w	��TW��R�Xr�"�^�i�l��0u��ǭG9�&�z�i��/�0����_�+-�*"<�k7ȔA���K�r�{�|�W��636'�n�<��*�P���4f��<� ���[l� g��#H�%i� �K���q��I�k�T��_���z��J��e��R�@�?)�vv�)c�a ���2e�'����ƻ�U`�Z��E����K]�&H�VS�S"8qׯC��~�6�ǂ{~��Vwvquư}1yA�5��N��Dfet�ho_��(a#ګ���(o8���[�1���u�A�5�=��t3���B�jU|�.��C��͓x����q �9:����U��oT��-5En]T�y����0��N	���"��u9�������ʠ����1����)a#��0��)��"���J	��b{܍>L���PU�x?P�<����i�}��?��M�,�ױn��_���n��IЇ�L�AU\y�I�3�klH �C*+�<�q�X!ph�{s;w}��B���ߏ+�"�@jc���=�����h~@�
�����A�:�Cb�_})t�bo=��[Jf�����Ա'k�Zq+T��m]@"=���9�����.��i��O.A-�"&#۞�i��}�8��@�
��(�=���JS���n�v5c��[�)�e�'��vu�a����#�
�ZĹP�����5���L�A�/	�שׂ�J�z�j�ʗ����9���S�&<�*� ����Rs�:��<��FJ��p1� &�NP�M�3�u����8|���AJ�Y�<^Nh=�RͶx���e6?ϫ������Ml���@jlUK�Wǽ���U)qe�*D�]P�X[L��d����+�ѭ�޲�0yF����V�`-W���M�!U֙����'"���oh�{�{Ę F�.��(��[�{h���Suk����}u�Zē$��U���Z�H4��� �T���D���h�E���+��$N�p#i�@�����,|��m�[8C�M�ٜh]ƽ˛gr������ I}��$Oo8�R�pE��� &���.�i=k"���W�L%�<�Ww��\#�b�cl��Έe�x��$�\���Iy�忏4VNVy�Q|!�Z���#å�EP5ǻ5]m���V�'G�(�zYo�2>�t�c���,�4�7��r�����a'��
�*F����7���)���>"��e&N"x,Lԧ���#k��l%�S�Q��*ˡgk;�P�h�Lw3�X��ΌS����ￄJ+�tǬ<Rm׍�Wu�Y�3� �.b�d<&x�E��@�Sl8��z�6��l��5Cm��SL(<z�aJ�uF�Z�1�-7$���n(ރ���h�w�/�R
=29Q�=Ы$%k��l���G��r3�)�'�����J��p@�S�B�{�j[�ȉL�!�h�M%�^�@Du'�	�T�i$"9�z+/|��Y�����>����=0�ZH�#5M�.ހ:�P/�olB���l/�k\BY �	MΠ���� �&��f�|�t���G�,r�p:�-ƴ��Mc���+>H��)��a�[]��2� ln$�D��6[��@�ϡ�:`�D��B
Y@�lN�I�a-Y�jD�"t܄!|���i`�+�S���:3�������3°tA�nǓ�����m���<m6Ô'���aV'�>��N��`�i��ÌL�8�eh0��<�l�i8��#�G�!i�A~�Hv���n��F}�\l�������ѳ�κ�Łd��m���/#)}w����"Y�ė;&!@�õ�Eϋ��u�F1�2���LY�~�G�#���pq@;-!bH��m]V��M8����*��>J��0�~�K�
�-[j-��q�S_ˠ�N�E�B��o�R����6T>x`�/�y�#��U��7{���+_��8L�$�ԡ�#���d@������e�¹�m$3:���P��z��5K�.�;ZT�i#��)�:��F��[�?>��i�kG|@��v�]�������8����X�ª{1�9ѯ�Z5<�rM�<J; �~�l��|��qP�vi��@�w���R�yt�W(��u�{�{+/��B�/{i\f��Uj�)�)uCW��<�w�q�{P�[���|(c���r���`E+n���X�!Bh����"���Y�2T�Q������#�g��r͓�t�[� g�[��7�M\���s���][B?jW�/+�֖~;\k��/}��>c�^.��â�Z� O�G�x����5j�p�Ԓ�ct�`�z�3��a�R�ok@�4�{V^�:1ؼ�~M���F��f�m�{f	�%r�B��%�MDX�5��E��2�{<-�.�]z��})�#V����K���ҡib���(𱉰G���t��G]$����'���3�.�%�m!Kd�(�� �4��Ym[:��l,j��'���u�mbˉ#�`��	F�@6�9š}�����"
�.J������\�	��뗊}K��r21���t]srl��������N��\P��E�����u�x��G���,���eϫ�nP�2�����=b	 �c୍x��A�������t�E�P��0���)'WK��:���iѰ����M�0����a���!�l4�r{���]^ݣ��0?�*r�.�ݢ�s�	hv��L��bE�%w%5�`v�$�*���jޥ����;�J�zj&�/�B�=�b�z�qoba���U�؊�R5ݬY��ٜ���ى��_���퍜Җ�����|_��&I�X��J��Mf�������J���s�:��/�{w3q2�&�v��l������M�������̊x+l@D1������\a}EݝMZMH}�<�
�����㟷%�ٿ�V�h��}��H�.��B���6�~z6�v�c"�n� �$��`ij�fUu�����σ�A@�M�ʕ$�G�2�S>P�{���(�n_gD�J_��j�EK	T6��>��c����F��i��s����⹈��ū������v����9����ʜ�MM�K��.��l���Z;s�q��2��-H�<�L�d�Z�\��vV�����l��F�Zr����J|�����!PG�6�{�sݩ�n�Q�f�g��b��	�5�u� \����<���o�l�A�X��߯�"ǽ��UoK_\8�]�!�k�3� *���D��5&��J��"_�Zzt��GF��r�մ�R�U���.F ?o֢~T��g91��um�{�Qf���&�=�Y.����Td�Քnk/�<Cn�B�u����P�`����Ot#���ր؍�PG����%V�j��$��H��0���p���^q�&z����ă��擑��kC�r���B�q�F49��]����!�?��x<X&�D����8_����E���0����������AVN2h�*��ђ�� �i�<��6���<�Ͱ��u5���˽'is_r��HR�C����i��E {X_�_��l�WC�0{\�������Vk���u�Sý�zǯ���[ ט��Y����@c�$5T���)yږ-���U5zvW?��S�pu-N�v�_L���qh������ԟQq��6�{�
]P{h�����8���3���2���2�L����#��sw0���N	)���X]a�
VS��2���5_pX	�
r��p��z-l.h��4�I	�|�zN�Hn�Cr?;Xb�[�{O������2��fr9/��\����ͪɜ�/T������ş̠(��H��z�T���р\<�H��a�s�����]�01w�$nxC���?:��/�%��j܀nG��Y0�G���⫛[��h�ٿ� jG��5#� ��!ĩ���#�!]�v,&yjtT���^��&$
3�Z۝�_�ېŐY����"�Ɔ�F���B���~8��T�(2�e��N�ĊVJ���K5	R�O��i{yx�iL���	;�L/�9�Oi9I����(\�8c��e��n��̷���#��S^ܡ㷾W��EL#Qo��5/xM}W��ڋC�2��<�*�ډ�"u� 2G��_���R�P^�F��1���I��W0���r>X71��>�h[O�:����N���������0�r��-D�^rw��e��p\�?*@�$~�h��)?��L>����^�󊕥Um#���d�vX7#�Hs6󔦽�NE�W��u+��N�����k��s'q����y^��Fk,g�l7����0��_�=M��g�%GÓO�%D��  �	��o<�Dm]��<4��@0ժ�lTŇ��iŞ��_'eUXD�y&UHv>�ɼr��N�	U�(s�b5<���́�q��,5�{p�\� ���GO��YPޕ�El�����T�V� |u�Q'��d���q�ZOV��[[��>�6������&��u`�#u�v�S:l{A�9 D8==4��`|HԵ�BY����v���_f��E��넼��;W�FD�ƶ�P�^�"�2"��2�94b��p���`����S���f�B�}�����(E���Z� e��2`�|Y$������'ܜVo���f���{ڤ���_��,fv �Σ���UF�C����!@v��f����׼Q���VOӃ:��+�^��qc@҉�*�����H'���/ 쓞X���*��b�~�zvA�w�Wl�.;��X8������� �9 �>�Ϥ�/���DpI��7�z��L�������i�IYS����ڿ���־w�P@�)�H�*Ζ�v�ҥ��-qI��×/��F���/���s��"(mV!��7����ȯC���M��e�e�G�+�Xf����=�[g��O�r�z7v��\.5�~�)�Q��h愋i�G9�c=>0��_�uX�8���$�$%B�A��v�H��p���X+��2�q�4��r/�b�p�3f`K0U�8,6C�#v�p��9�EX�1����Y�pPV��Y>�g\��j�k�-}{��7��o�ň�k,�mv�#��i�B����X#����ɬ�.��]fv�1[���tXV��h��[�ϗ�����.�����g�!���nU���җ�ο(�Q�B䧺]X_$�_G���W�%]�01�/��\0����L����WJg�"U��
X#�	�TZis+.+u+yc��<�R5�����!5���hM�C�V;U����3��JP��� �|�<��w�̿�jsp������c%�G�J�5-���.]��V# }؍�K�¥�*s�#��ޮ��);�����؈�0�,��>`�\�2�>�Ʈ��X�"bV$k�������j�t����d�Dk�����3ho���5`Gw�� �_��Փ�T�M���թ���S"��Pd�X����FZnR���{M���Dz$�����oV��9Vs�]��_�0��D��Ň~�h�\H2D)E��Z��x�$��i��ht��#C�Lc�x|.NF��5P�N(�3˙̀R��|��cܱ���3^a�����Fa���=
�_!�xy��hkz�����8\}g����.<�иN������nd�A��Uџ�14��˴�[��2�o<�;Nf������g�yi�U��l�#��0���~��1֖~q��FHL��;g)3A��Y_k�J���O�_Н��pf��pQ�����|t�'���o�g��$y�+����cw���d��Ɂ�v�*�L��T�/�E����|�SYW����D�B~gZ��p@yilK&ΡS���{�"�����Z�����PY��Z�_t��<��xp�Qt�@ӟo9�~Z�ۨ3���/rDJgcT�����;c�����E�x�
�bs�-8d&H��_-��u�΢��--C���~v��H[�P9��WkhT���Uڜ�I�J-�z𿧏�|���7y���k��@7�z�~	�T�EՄv���^Mg��L�}� K��j��ӈ��x=NE�#���Si�\�{��'j}��|ڿ�Dꂣx��}a�g�`�k8c硂Ck/+����m��<������p>�CX���A����������I^�ѽ�N�a���ބ�7iON�ŉ�ݨ��>̾�7},S��N�άgS��I���V���{/ 9 ���J�g��F�QTwL�e(���$���p�H�j���鱠UH�s�%2�� Ӭ��)��1 �~����=��[sE����^/���V�4A�.!Nd��@H2����1��2���UBe��D�A:��WꙘ,z�� #k���rQªW��p�B0���+�Ac�յ�A#eQ6���E���Є8kk�'�6_�㇂!g��.T��ؾs�+�y�� m���=��`"�����B��(���!0E>$�0$l��|��-�^��FGb=�唗���;A�P�ךi��%��ǘ�e�&$��n�F�/w	�Au��FP)�ch&�4Ta=}2�I�bc���"\G�ҡ,^t���þ��f҄���N�#�!��i)	94B2�d�,�x[����/��~Mm�P���i�fl̥�����'Q��&d�㵽���~+��t����q�/Ѯ���Wj�%-LL��TKj�z^:�;w��];Fbw�9�j��ں�*�%�Gn���l/� D1����ˤ�ϲ2̗��������0�P�!"��)�̴y�K���똦L��`Z�>�������Kn4o�w�c��[�������6��V���՜ ��a����ٞ�顣���H�L��T��\a0�$��\6l�N�?��z,L�f�e�7`ev��6����`���;86�?1��s#��]������8\>�g9���f�&'�eyl�a���C''a���?�O��i�����MR		�MK�\!F��I�zC�+�|<��E"�存{hYK��h��'�G2�7t�s�qɉ)"7P�ܳY����v���Ǖs��%�e�-wj �H��bq����Q�� 
�=����i�5�x�ڌ+�.��ǎB@Ǩsv�Mޏ�X�_盲�L6%}�0�
��xeK�p�� m:f�V���֠@�Z�Q�ZB�D`.]�;?������s|ў�2��M�g��3g��N���qno�l��Ёmev��3yß��y�K��gv|�������1�m�c"u�&�4�����>3��&c��`����T��u�j����tFv ���,��,���y؏�Ն~_��#a�N����w��ӊy��_����Ly�D�ћ��u�⌤~�a-	P�Ǉn�	�}����9��CWQ��#�H+UC'�a�>�_���?�i|z��2����⩔�i��L���� ��Yy0	#W�7#K�\�L$:Y�옠�7A� lkT���V���CК��#.����;o�x��FJg[h��8��-j�k���_�����Ѵ�"�A����i�p�@�����Rﳘ趶{}��1׬L�e��n��M~/�l���g�=o���4�3.w>#�L�Q (6�,�JyR͡�\��֎,:hL��ђ׮�Y彠f�HрtiD�]G���
/�Г�g0���,��,���=�k�":W�T*�s)̙�+OUuX�T~B��6�vB���j��}[�;��֫����q��4:��Q��p��"|��9~^���>��<�W�3WϠ1��>!~l�!�E'3	Y��	k��w�7�3�	n �[�o��T��'ZU����o�/w) �]$��o�B�����s���5/���}�Qx�HpH��ޑ�5qq������K�6�D�R���u߹#���i�S#��=�?9�2SG,���+�׍(�o��/c1���ibIno�<����AJ͞0���)��V���.ڷ}�dCSsF¸<~?�Nq��������#���`�Ρ&��ay4����`��Zr���X������R���o�)?e����O��#�3��,W��wT��	I�_,����q�M(Vt�;P�!�_��&(���?&�L�:�	lA���T�?��t���:N5Lԟ�%0pg�o5Q@ZB�_�YW�M�ʊi� ����.]UDU(�:��6�B=ac�Ng�z׃�e_�[��O�$&��uΚޞe�%U+�M���J
�G������h�m�c���+�9F��WƈЖy8t��Ň ��su"1�!f8k$z�Li��{6�~)���z.�C�IV��)3�$�bX*�g�&�������>��)��}�ئ���F�zuU"��C�l�3��"�2����{�I/���/U�X�*v``����F$+�>�=�;��	&�>��MC�2�̃�[꾳��Lp�Z��/}�H��eb9r`,�w�����L�튫��G���IŽ�Ks�޹��TCy��9�w.��ۖ�F}P�}~Sr�/J��r� �u�5I���F�,y��3���|O���DW���7�
ʃOUg��ʥA�e�r�bt޼�EY�)�͹;�|�V�0�H���A��x9`�T�W��T>3`f����_U�@�Gj�r��@�):�Fۇ�q�V�v�C&E���b�
��K�1�e�g�p%�t!�{*�^}J:�P�J���@�L��.��"Y�/1�!�8U+<��`u��S⁡��ژx�;J���G3�gjgT�O��\xw��$���G��V��8����6V|�ښ�@$h�����5��Y}�E�en*T�d�-��4�^�O�[���1�5iV~qdʆ�p��1e_��N	Î��_I0!樓�F`��6|���M������*�+ɶc9�q��cL@�3����OY,�����cCE�
�͙�aX`������R��A�Q~�����Ҕ�������Iw�<�A��T9�$� �9�7N��n�9���~� ����������v�����^��Y���ֽ��,Udr�ue�F����1P�u�+fDϧ#Xܛ�B,��$�t�H��7����7��&��H+3Y"��~��;��Ǔ��*��Iy��п�*Y�Qլ��9.)�&�F��ɽ&�L�E��ݮa��9�,��M�-;��=VR�?�����u����#��{����+V[W�OA��E����0n��ͰQ���F.L���	1��壑�3�MS2�'�}i�~~�
�HW	'6�s �y���s�� ����B��E2=��6�ޝ�n�S{���C �.���PK`�s؂�s�p�c��t>�������Ƙ�6A�Q9��d=�ڍ�_D~�(U��r�o�2�5�X�ȍ�#G��̴�6~��{,��`tk[�0a�S��{���t����y��6��:o��o�Ǹ��ϐz�
�M5G��B9q.	�����98�������$Y�/T"s����Q�O����u^�<��gN���8�k�.�0b;,1,�7QV���(�I���}���V�-�>�)Jڻ]"`�'�1�"�}`�w&QD�D4;��?$C���u\��������P��?�7w�	���C�W��pĐ�;�>�Ez�M��������4�'��FG(-�S���ϦH�̙w��. ��h��(��:I}����%�p�����LWͣwc�k �%^��"t?�	hE��S��NlQ�N#��?���	�ⳒIha)k��{y����l�ߚ���Iq���uT�bꬋ��[`��*�v��n{��2X9*�d`����Z��1X�Q�Q�������L���L�NPJ���G�P_���H)E{��@i�j�d,V^j��	���{���R�¹?��:��L�4�h?(p��K<�3���C�����^�E��O���m���o4f���������$��Tp��R�I%jg�����4c��Z���s�ş�>��!��k9�����ў�,5J⾜��M)@6�����(.|m4���	�����L��������_���e`r`�Qk_�ŀ���[M��DzdեdrQ�U8b��׳�ԧ� \W�#�co�Cu_
-�-���
|�����:�i��Z!�������lMg�砗���0�ٿ%_�9QʁpA�ծ8>��%�Ɲ�a�b�˅5|�E��-�b9���3���x�γ:��.�F4f9�Kُ=�L_�Zw
�\����@�ٖ�%��ܹN1��V=��ȷ��j$pP!խrMh���VF�}�?aA2���j��9��a��R�#DV94�6�&�bI��K&�����믟Ƈd���l(IN���=14
��#_�+�ďe|�aդ�eյՋ��((�F�u �W�!��D(�Dfé�N}�%è�jU�U�?�����w� u9F�ہ�D��.��aa�*\�B��㊡F���}���<j�F�_�ǟ�:�O�K�ke�Y>�T7��$�M�A���1�.��R3�:7�i��)Xb{�I���\.��s��A<�b���;��_���}�e(RĐ���=�jKk�0�u�Jz�Q�-����� l,�o���Ɓ�4�ux��1�9�B68�ΰ�c��2��%��O�P������o[����l�p���kCn�A+F.��Bda3,V_��N�ʥ�u7�����?��<wr:��b{:����-�խ��g��s��^���6�=d@�6f'LԅQ
����X�����QI����.[l��B7 ����h"��ϫ���m�e��Y!M��G�O�� W�ui�eK���wz{c�π��~�l,�b�*�A���yNj�x#�)��l��s [4T��߅]Z�.�Й�o�=w���߁��S }�K��c.�g�D��^zW�����Q*�5����+�T������1���1LG�/j���<���Ù0o��r���I^���>�t������_��4�	�]HA���'��o��O�m/X$��� _0uoN���<��"����(+|� S��oI�x�v�I�����'��Jk���x�-ZQcp���)U�3�Jã����J.��Z���f�B�w�.k�o�4׾����ѵ1${�m���إ {��̡��r���*�\���*Xd�$��qk:ܳ�����o��d���3�;Q�!ɲl�"�Ӗ���ƕ}}���X���K�u(H(�½�Tn����,���?����THRYC�c�����؋�v�ژָ ��E��U�[b�@§Vm�B��U���1�dt�DI����m�D^�g���U�tdv�M�@'5/Mk��A���+�7�jx�g>����w�=8�G�:��g"��dhيof��Ld�#����Ց�!��)W�d���H�̹B��C��ry�b\|�©-�������A�k[A"!������%�uV����l"�ľJ�3�.���t`1oyr�̴����y[�'�Y��w�A��K%����zw®�����f�KN��;�Z��u�-�%�n���kOL~����g)��"�&��qBv�b蔧��;�ūo��x�{ƚ#���~���Z�ʆٟ6�[�M$�����y�3;��M��SPH4aKI�oC���Y��ř���U�
�õ LIK�e5���Vg���:�n��;����a�I���-��4W��Ih��޲=h�m*�b|�[J<X�;1G�z��)����E�r`�[�=�v����N\uiU��-"�FP|����5O>;{O�\��[
xB˷풊sB���}e�.S=�����EүY�Ag#x��B.��@|�I�9�*2�n�J?���l��"[W
��z����m��L�<�?����槃�l�ȸ ͜%P6��J�Z1�w��SK�����1:?uP��\������w�y������ܥI�;<C���q\����H���*�J��ul�%�������b�g�yD�Iڻ�����J�.���	��N���	�V ������������T�||&>E7�X!�`$h\�[9:�B36�/��ri+�.�&���1��7��#�j��T�񔱊��,??�uzIo�Z�\�Q3.���)��>Rr�4ܙ��PR'N�)�N�E��*u�	��C쏢�yw w3�|U�x���� @�F�̸*d����$��B%ԗ�cr�9k��iA&Eht[Ɨg�	^8�, ��^�V�_쭴)�6ƲB����e>5��dݴ�j�
/�^�����\��H����m���_�;�c�ZR�I�O��?3��u�t�vMS^�� ��j�h�٫^Q2,���ݼ[�w�O4mɍY��U�c��(�l�>5n�����{�G��F�|H{�/����x|p�Q��w�T�,̣�\�z����g��l�`^N������wǣ��-%K�\q�{.�XK�!٥y���j��89��j�x�F������_���]񐄐��˙C�~����}��4^F�]h�&��Qogi��t�_�%w �KEN/s�%���qG�_x(x>����A�< C=��]��7����-�YK��18�D���V�w�)�RNc0W��0��&v�yY�ܿ�I�8�&'ʘ�� ���16i(C��jnT�
����N��Gv���J>����↔u�ԗB���{�QS����6; �(t�����&+O�l��գ�i$��s�='A�(
�S���)�y����<6X�@�gg�W�[��!�{s�ɽk~�u�\1a
����j�KX':�A�A定�C�'��h��#��Bl�R�J3����l����e���"�)��,�k=8(�@#�����@}#ԷN���)���t%��v�e9���,c�:zS��ʨ���Ԕ5���IhɆPP�cN%/�(�"�®BH��K�����x��w}ؑ��]|�BO�b�-�Qqw��q��*�5ͼ?�D��AKk��W��M1��F0���Ov�7s0N�k\0q�HRl�`�A��A���8��d<3��}��	��7��*ں�%O�\wp�����q�ߢ{��[�[j�M�r��@4s�Z��%����D�>��+��	%
�pR��p;��	�G��1jNtCF��1�*k��le���k�{�YL�0S�(��Mu�pP�'�)?\-|?RQ��j�N^zM���v��9I 7���t��Z�d���M�<�+�����-�C�#T�d��g�6՚ P]���ZJ	O.K�DhoU�ҩ�.�&��^UF�u44\��IEL�LBB=�KP��M,�<��:���BTX�U�?�~Fam�y8�ѹ��;Y��@����$��n�E!~�D������A����o��^|�+"U�4��a��O��)ɢm�aH�����cT0JP?�457)�L��|���)P�m�Y�b�w���O�')Mů*i��Qv� �
cO�;�<+�G#�
m������ښ7�~�j���M���~	�p�l��H�����	��k�B�1�.�\�|��Xj_=�M=1��5��f�.,����9�͓Ҧ�!�"����ٯ�?Lm*8����u,<�T�g�����9�������<N\��h�rȍ����J$s�u �ևg��m҈/�2FU=	v�lXY'W�U �x��y���j�^����/�ū�z�8�~MQ����m�[�������i��o�nъu!�#8�*%d�Ӽs�j�a_�5;d3�<U�V ���:���Nk �rS��5t[�m�O���w����t��p��p;��f-��/�����/e4s�-�+f� :������4EFgѨ������ *�Hß2c�
2���C��f��Q�\��q��T��Y�i����i#�TB���畫>��!��d��Ĥ��h೹ WU�^~�j��fWapo��^�����.U�X���U�6Ȭ�WX�0*�RRɉL�\�����0d5,��ϑ/F\-z�V�%˂g�n:�T����O)��>�boT�dzV0kR�E���T��(F�&*�s�e��2N��a��V2"�oKj!��Ҍ��uV�J�m�MN]_[�3�n�7�G�~H-;od���E�ZuN%�OL��w��L�#C_.���F�S�JKu�y��8"�)�1�Ch��>�(v��7
��ޮD)+�XP��>�kJ���)N�r�,"����̦���:��d��<�A)��MEc�UF��w�i��J��)`&�	7��Su]�Z�/-:����äXa�Xk>&��bƅ�� �v鬶{����8ا�U�x�5���x<'�M���X���y�.�@����YM��v5;�5MЃ�z�W���XR�c���0��s<�ԏ��H�t���d_�N�
й����I��s/;E�}_L`d�N�d��w�v��eR��WVH'S�lO�-\yR3�!]��n��p��YiJI�6^�+�D{�960�g㥷$WG͖)���ꈘ�x�vV�e���i�`�����Bx�QD����i"
x����ր&�DXi�y�G�V �SnF-�ȟ\�R��7˧2�Ы��x�1��wi!�׮�Mu���E% ��:��sj�l����ꆦtSV=cA3��Z�3D_�]gRT=1�� �>N1���>�w���錼ro�8���([l�/[��q��u��J�#�ш�,�#$��H�΄Z��^����<���j�zq���I�<��Z�~,��<���ә�� ��E5&����D��iƨT^ĻؚQ�W_=_�Jo��Y��0o'#��:��5N_�T�b��*�xyyR�{����hS�P�ˉ�T�Iճ��+ʣ��o*�Z$�}�v�6�c�t�zot��n�p��\��W��x�L��H�{��$������6�k�*M��]�51�?���(���S������%����_!)y����Eaio�$���#��]Y������ho�>�sq�4��"����sr)f�G
�Y�Ϗ�����q���};m$%A������
a���0�a��^V���R%�~��_�%ծ�]��a	M�=qb?�U�*�`�E�£���'T�Dez7�����q��%��J�<��Ԯ7z��K�����i$�F$�#)d1�o�;���7N�.uN��+��wq���P�Gv�=���1�T�<�wm_����f:���������
�R�x�4��ב�Z$�_�S}�E��PO	��
+�U������͎n�R	��da�-���� ��p�g���v��x*P�S�T�p�J�_��w���'�
��0�S�!R�"t�7V#�_��	��>�B��++�	?�E���4�Aa#��~��d��S`�2_vd5��o���3G�0C`�9�0-�k��k~0�l6�%ΔQ���^�%����]�K�(��g��i�-�ִq��Vu��Z���C�Yaəq�� 4dq�j�W� ������!�����I �9}l`>.���H������4UX�Oz�bQ�2J��$r��N�E����b+_��9 �i���2���u^u��$�m���V�����/od/@{Ju��k��=�+��'Q������fP�6���v$��荔|���g����eΩŶ4��Qp��'O��U��O]�(�	��s��.H%y� �"�+�NB���u��c��	_��]�h��D�Ū�M��]�~���6�>[bl}m9�3S|֨�{�ڳF�h�$\Õ4�E�7+��6� 	6��y��`�SomXG�x� K�R�C�!t��.em��G���e�6=%E>�}E���e�x��Ԩ3k��}�ȳ���J<�13D7���f�Ԝ��$Q�l�eXV�J��-��Ǫ�h��?�����.�._�� P�F�o|�	�U��w�C�	�7�w�}ꖹ��P#�{���e��c���� $����%�����uV-F��H���:WB�*敤v;Y/6��0��ÞFC�F����K�C����36������a	�2�dibV���ӆ�w���.Hqk�y�ݖ�SjxP�(��{�&r���	��͸�mtd�������@]���wfz��L�Tj����s���.�Εij}{t��R�����d���#r���H��]D �8C���)wF.�TĪ��	H/'+ ���1)��7ͽO)�F�e��C�~�P�t.�D��0�)-�y��W�ڱ��`�g1)��I4��B��C���%i��n�{K������B��F�#	��h��8:�(R�v�6'T^4�w���Ke��h#��Vv� �|�F��B��U:��H�����{;1{�5�$�#�m��0�S|,�>�H��p}��PH�qn"����8���?E��7�-�9;_Wg^ݴ ��x��]S�,��UҚ��i�&wٜ��[NED�bz�@�֪v����	�N~p�	z�n�j�d�7�cp~�F�'W`��+��s�6�Cr���n�N��Ū�d���dSb���n�A%����&����\7�&������Wt�Qt��t�E���	HD#�oK%ܣ�&�յT\:�xȲ���	A.���fjR���_T��w0�U����A�Bڒ95��`��Ğ�����	U�J[B��fiWe؉��w��(P,���F�a��,.]=�<A$�o�/�弞$�=aF"�T���$�?i_�)�9#������pX�8��_w6�z9���O���"���(ɚ��hZ*4XtW�;�I98:��=ƺ��o573u{R��#u��H}P�Tsm�x� ��de}߄��&�U?W�ؾCa�u�Q�K� Mh�q���yl�b�^�G�!�L2}�!�����G����SA� '+v]���5�S
A<��XDV��EA�ω
�*π�z���$�f6U]O%�k~�y�u铆 P���Z���O�#�6"�az���xF�jg���%�b�3���ߞ3��Q�G`#�o��F��i��\$�/@)���=}]=Ӈ���G9p��8r?,r���}�0o]*}��~DG� ���Q�W���U� ��ߕ���'����e�-���	Ld�p�e��!�=�虪�_2��NB�����_�/FM�l��Ӗ�59�2�BpbO�����*��[�f��O-��)�_�g��D�3�2SpYՖ��c%uR�V�������Z�gn����L��s�%�$�s�.�����=����EOsFꥤ{��§��dpV>�����X�G�CK�&�^w�܎e�S�(���O�y�+��xB�OF�~�փ���M�a��/K$�V��5�g�%����i��cܜ�,/���Ϗ
�҈�������F՗��=h�TW�q^��q?�;���������`�j�ܽ �DO���X�(B`�7�"�s8��y3႐��Z��8�N�����Mǉ,�QG�(����.�� `�*�O2'�b*w��,f���L��8�$�Z���q0WO�ni��%�r���	#.MK���b�d����s���є�V���G�9�ذ_N��/X�����Ԥt���Ǡ曔�<W�t~��f0�KX(G�v����/c�X��(�*�kT��6WH���Tj"��˒�T�rS�	[$Ec�Qp#i:a"�9~�{�h��@�P�/���C��X��$~rn�������H} �z '�T3Ɗ�z�;�L����q�uo��$����7��n���wQ
�GI8!�ƩX���H�4���'΢`�-(����H}��p��B�X��|:���<F-
���!�)|;�L���B�H@��3�iS.k�y�XÏ�ᑴ$u'�T�,ӎ��/�����ށ4�����?�VF�"�	jx�������Yy���V���pn5��n����A���lka1�v��7)x�œ�2k�½���]^ .�ׅ��Ik���륦���L�1*����ϫ*��4�o�2SK�G~�w��1?S�����@�}1U�c@"�;��y7R�|�`Ӓ�0l~����pL�i���b,�ˠ�����C(g׌#6�O��p�)����$=ْ|5�4����'�������FK+<t��I�����I�-�|"��y1b�u
���9u_Q��8� �UĠ���S����>6B�Q���N�'�)5X�d�j�
�D ����S�A�ik���>�oEp<E�:d�q��/oQ��YȂ�xG���3%����/ҎB� �����UɃ��֖�ˢ�cj�����.~11p�[Fe�'r=8�*rY���k(2;c�1��ֳ�I��M8�u�c�\\����`�HdT>��Pb0N�X8��vQ,�����*�X�"j�Y���FlE����̐Llӯ�Dy�1�`#>b�l	;�7�Zo�,ՠ�\!�����&v5��ex����k�Ӷ��;l����T૶��N���$o
)�i���f��KL�}w�<���1�Id�Q��@��M~����`]��W
?FF�0bMW|�c���S��0p�w�l��ñ�h'�kq�W7{���,e�폁��$ע��۹T�2s�vN�������r�3����ZM�ɴ$��zᏢ�� ��-���
��2�mO_U� 5��Uc���x�1�l7�����(�o|�b`'a~M�i�ܻ�c^�'��ޓY�/��z`�p���;{v햌M�K�E�܎�\�d鶘s�!9��Y %�ۢB'Ɖ<��ӝ�\z�a2����^Z;�YLS���e�h�ƣ�,���o� P�k�����]r��!�(�{��@��,�V�.����4� ����f���FL(O��t��_��)`9����G�:�ٌ͚kxU*^�x��s�1��
F�N"����t"���ȹ?����ᄮ��&�7��g����lF3��6�K,�}�����lH���)xi�P�T��S�f'krh�'�O�{90"
R���pK�ZT��͚��Ц[��M��p�6�Zl��}�\�����5���;Β^9�Yժ �5W4�#�%1J`��e�U m��y�x*�� �(?���f*2<%�A����QjF���Vq���m���E׵h�W����I��!`�>�9Z7N[ R�+ ���	V�X�<,�rOJX�V��f��&�������W�d��p�}¯JQ�g�t�\��'�J��j�	(��j9�kOw��H���=�`��.m\�8��C��y��^��s���������v��y�F�$�9y?
�k��y��#��EY��U%�ac�<ʍ�o�f��j����;�۳
{p i^�\�ې���0	@���e��"�v�#���[rih�v��J����+h��S�̈́�>Xi�=���72Q�(���9��3!��[������f)��bc�*^S������}�IO�˳X2	�ֵ���?��\�!�G�LfѲ:��8!%���ڍ�F)��/�{��ҬF�T���2��Z��)����K����]��"l�p%�}���eQ;� ���/�����
�o��"�Ы�d�����6��f��tc����b�s&S������pb�~;m4ĩcJ��k�޷~V�Ki��g,���5oz*K�7�5zTҥ�O]�Q�<�i��E�$��=�-n�FÊr��ތ��(�hJ}������1k(
�:�r���?'5��&�#ں��6�e��0MlG�ѱ���zc7U�Bu�"n�GXL6_���iٵ���ٴbF�C��p������[nΧ��r�:���7=7hO�O6۽��Ov1��3�u@,'-[`q��/��*6djb�� |��1�#��@���s���ܼ��m�� ���6F,:���sn������_�+M����I�{Ʒ
���7L��砂錄�Z#���6��Dq��%TIe�GWc@�$�X�+r2�B2�kA(q)�23b�l�a��X)�[��a�!1KX����/*��KD+�>`��ô��T	_,G�ky�ַ��IN�|qUXq�I���f�geF ͐�]�l�6�W�nNgA��6Z�w��z�S��%'>Z,y-�`?N�ZR��#�&k	S]��F2>�D�V뼩�pN/�a]Ʉ���<~%S���V�h��7���*���!r�~���;v�>�k�A�mmpշ��v���6\�� Or��
�A-/�$���Ӊ�Ӛ�"����p�8ƿ�kv�gq*�8����6�,p�.v�n��}���D�R@Մvx����t�rk%\��p�{U;�m��݉,(�fH�-|��	 �� `Qճ�`!6yxg&�і�BF���� qƲ�7��ߵX��h���e1�����[�3��S��:'3�&��9�>z� h�_�2A|r�
<�2I�j���GX��4�`�נ�}(�}!�B�Av>�Y�(��_v�wlMY}����O�J������lD��	D.�Hl�#�)��5����p��W?Yi����d��|'O��w֜5]��XŴ5��Ð[��?�}�2:�F���|О�����g�v��Ώ�v�X�W8���.I����=�}O�.��ү�_t���{@ne�9�Ȟ�B��ϊ�:^ڕ���Q�ſfܦ����ň�k鐸1%�ȯ�ti�\7?3�C��S~���P(S�,Z�B���w1P�7�����c���[��r��M>ˋ9� w�'��><w�9��Aӕ�8-q�G��m!��*.l�����������2�f2�-�r|�Q�~�eq�� ���Xey�e��돮C�za7��sm_�� X+,�ȔjJ��%�x�o�1����a��6����#���$6*P�¹kdFS軫�aŴ(��_��}\L���;�����^��L�>V֮üK�$��_��+g85�J���a����_ � ��v&Ե)Z��:�)��OI�+��,�p����u6�=B�a���s��ߘ����B=ٵ`��M��jQU��W���V��'�C��C��e�$iQa�ĭ�O��luw\\� �@`K�fE1�	�I�LCۀ���<�Bt��Lac~�_f�'���O��� ���fi�H�H��!��BJÀ�!�Y�Aӑ�Jj�� 
u+*ݚ	��`}�R��ܴ�uDl;��9�ｾy���f��6���eS�e�����:���
������Z��I<��6�l&�l!��k�VE"����#�S(�́�H-S�{�!���~h�x<t���͓�\G��6b�l hA�Q�!i�5�U���������.�])��P��Hl����	@k.���u�&�+-�FKGr��mj������^�q2��_�è��k]��0�9�ɑ��=��ˤ	1m:���h%B��U�f���wk�}������S�l���!8-�O�<L����.q�~���'}����J(�5]��Q.%���@Ñ�@Ɛ
]���@U2n�d����ǝ�y���h�?]�U��70[P�炙kj3�=|�/4Ե{;^���'�͆?F�\O��˃.��*7sn��vZe����3��r_��3p��j殗L3H����5����� �k���\�2��Un�6p}��=o]��1��� ��T�1��{�O�������$A7�P����O��5�i���-�ٷ㟕�U�7A������oO��
�r ��
�o"�W�Ϋ9-�,N1r,�@����5�7
�q)a�ʖ�m>U�صu?@�G��CD�w�������iUL[a�a�1�;;����*0��6������[c��
���t=�T"axy���K��ДǢH՛`P,uN�ʃ�'�]�J�fѨ*{L�F*�.��Ĥ���9��;�)�S?!\�0�oP��j�{��Ë��^�RI=ä����� ����)��W��7u�P�t֕��
>�4ϭ[��S�ia��V�3���㊌�_�;������!�Dۊ=<����"�Q�l��~�����]�������3��Y����9���d��r��<a�}�7�
|��@%�[���Vz/ݎ ���F}WǚC�fm|�ש��a89�ߵ���0��8�q4�P6�e�uK�V����Nq�/�E�QQ�La��?��~��EkR�K95��0�?��%�7墽��=�X��O�|���E��ea2B�y����3�	�	�	�$�V�Ą.҇2c�wܖG�Y���=���R�?"�sg�\Xq�-�-�#����_`l�����j�=X	:8��x
3��ȳ��$J2�x9���x����w���J�D����P��o}�-2m�֠�S��	��ö�P_����6�t�&5.�Mm�pS�sιb�17�b�r��^j�ȼ�Ø<�q55�g�)(��#z��;n7{~������a��޶��n�O�K	�&	����x��;�Z4�����"E��V|�Q��)Qj�/g��F� � ���7�B���[�=i��A������f�,χݯ"U��㻂�<�hAC�m�v��CE��D�>��j�!����R�r��S��~(G���⸸��V��ƤH� ��Ɠ�C0a6��ү}x�x�eܻ͏�ͧ;�KO˗F�.*��� �^\.�9P�0�K�H�iG��?����X��I����F>����{G@IZ7�0\/�"�1��?��ʦ�����9ɔ��R<�p%	�gI`m���nY<$8e�Lǥq���_�𪙠mp�g]�_Ik���S�ߢ���zWʫ7��M�L�"ч����jԏA�s�a&��-��T���"N�N�c|��M��f���E"T�eN�$���Z�{A� �����I�Xbp�5$�B7��)��$Ŏ^2N���.�� �;I$�9\<S�����.�5�#�i�����