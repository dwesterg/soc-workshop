��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,�9���/���]N��E�]שF����1Z�#ߢ �d��o2����TS���(� ���3N����$�F5l�@
r9|~U����Q�d�ݮ��+�4%��C�Nx"n��<�.�����U��0T��'���w�Q�z�[��q0(w&���|6BP�4=�����ٴ3���t��W	�Aت�� ��a�͌�09�\�<\����� �f�v���%�z�M�7�:A�����k�;W�qNI&�Ǽ���Oj��PuS�ق�ӆ�k�>�N�ɔpe��$�t�1ĺǎkޫ�ΔZ��I�5�u9��D汁w�#h���,e��`���/k���ſï�&Ǎ����tX�.UI)�a���t�Jq��n���tO�Ψa�70����nE@͔[�;��xq)Vot���Cg�q
A|�w���;���_;�	���ި5X�� ����/�/����`�9u�K�n��Ɩb_P�b_�`PTo)�"q��P�?$�ir�u��F�1���m0:���P�e6�J�����T������HU�s̩�^E�җ��(�6ݯ(gh<�U��&eI)��l0�����π�.����y�r����خR	>���K�I�ߊ��� ��<� �)�Txw)�Ds�EF~�l'"u\:A�IC�tX�@@�Y�ܩm�_)/-��|���~75M�.�-v��?����~��a���G�ű���!�=8�h��8mI�'(�T7�B�6^&Р�s�i1�6*�29b�ha(��lL�d�����fŜ����Ф� �d� AJf�zI�Ǥ*����M|���M�Fu��L;���2Q� �����u!�"��V�a�ؠCN�IW�����=���N-� U��!}��j�����~���d�k�ƪ�(i&�V�����ͽ�æ�K�ӻ�p��\*��5 �wʀb:�$)���<e��#�rC�B-q5���[&�Z�?� ��
ye�r��������v�3� ��Wl����ѫ�du����#h��j��͎1��<�U�.���K�4{є_�-�i7��d�����-O&1��D�޵{E6����yw'>h���#�OFx�d#�;7s�(WU�~?�������0�� &GBX����'C�~�TK��1�����T�"�~��[��;�D��#�$#���=R�&^����n��<-<==��J���X�v�l��Ic�2���`wH��&�	�)��,�B׋��=H��4TX'핸��s�E-_!�sT�n�`q������@���hۂ;"w�l+��sr;�3{}^V�8.��6��jG����GPb��qڵ}D��y0z ������ce&�Y�Rk���,S�Fc$��y��T���� �M���Q�KgD�-_�y�J\�AC%[�H�0.cǢ@��|Tf�\Q�oT�1�{ �=��pz��T��`.��)x�'�}c�`�a�o�7�N�έ�s�J���_�س���P?���BJ�ۦ�.+�b'��M��HZ�l�S3�v���pt@��sv�d?S��H�����k�Z�zA�:��K���?;��H�in�ݧA���F�>���G-����0���[dn���l�Kᔮ�9!���s�9�پ ���b�`� [�8��:��.��<�21ϐ"B����q�B8��Ҵ�h[wG�P��4?.������e&A ���)�1�`���x]�7��:$<{��V�mk�M�)���q]��N�;u%�`A;_��C��˯����lp+Q��N�8~���lKq����p��+��Mp�3q���ș��'��~�3��
n�f�l�jb�
���ޭfӂ�[6yQ��G�� w�u���p���6�࣢5�/BH��%��4���{���v�G� ��`2�]ٰ�|4}��$�qiO��Ʀ2gQ�(*X�fla�1��\+��m)�c7�~"K
	R����w(t b=�;=g2V�?q��r�胵������U`��+�%�t8T�K�`��,ŨB�>��x�Z	�5�ꀕ;�?S��aq���)}��Bw�����F*Ge+J�#�mAN�q�q���5�9�]�F�6�V���:��K[�5<+���7/���.;���mͩA���!��Fq��V�q�]F�M�N�JT�ST���,�i�#l�q ~�YO���9��Kg� d�N�-�p�@a����'�=ӯ��L���֌���T�xJ(~[��H�E���G�(�+�,n_'�-D2l�t��%m^����O�� ��%=V�A��Q���@�K���@��όV3e���i�bڗt� ��� ���A�`�nr��6T���98�`�b)mUM�$����$�ys8�J�+_�2j�6��;<�$;�KPѩ&>���d%�1�> ��ң�MS�K�۩��2/�AL���߈� ����ਰJ@�A�UW(f����6u����RU��"�N$�0\���]�$��!S�`���˰��0!4/#�d��v�ϦI9������7s6�E���1Ml���7�ƒew�ǜ$���y�r�3��I�$�|��d߈����/���� ����jf9R���[���4��]lV����=!�Ҟ#��c�x���;�h�KP���l�v�3�C�䡰|�ςLJ3U�Fr����̫���^���yB	�S�����־bV��Oz�UVד ���K�Q eM����&`�������M��-����/r�̐��i�jr"&^��С�̩��	: �@�Ch2c�A�|ð��@_�]!C�<���fi�K|�$��-������������a|f��T��:.�B���T��-���< ��!FT#D�H�:������WQ�Y�[(mt���Q�u!�жv 	=�1�M��7�N��`��:%��4T��b+���2��ݫXׅ2KP>�m���D���W?�wώn�s)�p����H*���^1��=;�����c�v߫��Á�i��g��`�dKi�p��h�V*r6���%�����m��&�K"h$��s};����Gi$�{��	��kyjv)8�r4�=�Y?X(b�QL�1�D�CȠЅ+ȳ��/��Fx�A^�-�J�l�ϫ}6$�48���O5N0L�%A��3�rOF�<��mO�N�.&�KW9B���RX�(�K����}=A������s<���(6L��=T��o������>���G!��1�ċ��<��;R�U?��.qBA/OS��$�����a�ᡄN���qLD"3P��Ha���>{Hl��PS���)�Ʌ���,���|x����/$���}�jx;� ʼ��	��/9��%Y�^��愩e��n�r�\V�M�"�1W�C�:`);��v�d�(U��L�����*��&E���0md��8' �1���DO�?��k�I$�mh�q#)�R��Љ����Gl�Q%z1���02D^^��Sp�V��,p!�es���(�"oѥ���7�m�LD>F&�(���
ge���^m�/|DS�W���	��hg�����<�3�Pa�Ej�]��u�_H�nWq�(�m��28tg�#��U����9>��HA\k�Η�븘2.�t��\���^�,�����
��]�O�)��|ʑI�Ԏ�$�F�J�?�n���hYg�������ah:�Ϭ�F!�P����(��c���7�������(�Fyg#�
�����0z�T���d�+���,9v��t��9}�b�V�_�E��Au��^�!��rN*�=ͱ���;�\�$=�|Ў���WN�I.�
8��Ҳ�`�1	W^��.Oo�-���?©{^i�2�p��g���/��deS�ֵ1}1� ��Va��t_"t��w~���d�e�ZU}��B�k��p~����G4k�V��u'�0yb�cZ�V��d�(��&�	�F���H�@����2�y��k��h�x�n�q� /o��~��ԭI��u��U�D��\�i*��ј���E��e�k��8�DӓN���b��ұH�ib�i`1�x�Q\8H7W	:*r�n���V�g_!���5���`�j3j$��=��fYK|�v.g��`��A��*E�ԃ �F�E��?f.6@�sdt�?���Nd1�8���J�m׆e�����Si�J���Z�Ы0�*G���Od�"���% }����+�-Jq�V�,!F��������y�c�	d*���`�,-�ʒv�Q����'	�bO@�ӆbJ�b�N��<hҬ�fZ>�*=`�	
?6߷��;��g5C��8r�~U�,we��"�V;g���GQ�g�S,E�,���ˬ�^��	fQ��� ���go*��[0ڐ��Aco�g�w�6�)?ƺ֊~e�M��t0�60ؖP�fxj�y��/�3X�5 u�3��p+*�6����d�e�oz� ���4��6�7J���4�-ɷ3�6�A�xj����x�@�s]9z�L0m  72$	�����+\����o�s8Z�]KP�$W�F2��\�� ��q�h�  �\�z����-:�&�̵���ޚ���tV}�w.�������y�L�Yx��]C!�Z��ꌀ�3�����w��ߎ��qz��wk�`oI2�g麉��B���nϑ"ma�I��6��l�&��7��s�{��`&�B�X����ň #-	�;��`L���}��^H4���Cw���u6�`1�2��i�XTto�[�K����~.�ԵȑMǾ�_o
�D+��Gua�O����A$S�{rƲ(B;q��I
����3G�v'eݙ�]l���)�$;QM���yf��cb�Ѯ&@�D���5�!`g"��	5�]Q0u41�.���X�4�|��%)��*��� ��8h�������6쮁�_�!\;.�%���B�[5���rV����)�Gf4EMURj��DM -GW�j�ֵe�~k������?U��G`^��z�Z]�k���gi�r�-{&<��Q$Nu��<8�e�;f�5� XzE��eF�]@7�����l�r�I?�A��O�ۨg-W�op�zee�6;�k�;jX'��ǒ�gS����%�j�BX�oBzJ; zoǁ�(GX�O����f_�on09�@�R���y�@��~ᾩ�����1�t^��+�����33blļ���P>s�$"r�1�Ȏ0�+ש��v7!���jЉ��-y���S�g����9@ή�>uHϏ#��>������(M�\�@P����|�~����;Ԇ�ʳ�; �<��|�Z��FaK��х��j�HkLWx@��; 4�F�>F�O6�(K�^2/�%�OÈM0�i������ؑ��i�$x���E85Ϡ쳫̯$|aAdiA�T�$ⷜ�o?%�=�6Y�s*�s_��	3��k2B2"|.{i�iË��}z����ˉ��qM'�R鉹)(��:.yV���=�eࢢF�v�[�lwH��fx�ȦC�pÉE|	)�1�^-�eA�C���g���W]�C����u|�k���-�ӯ������r�vm�l+�ʝ�3���R�RE��N���z�"��Wd�:���ԴSYN���
�h�a���zC>۰�7�W��[M�[x���a[��(Xg���p����߇R!f �����!=|�=��T�g�N�>Q��0���E<�0�e+��)���		R�gT����J?�T_��޲��[��90f ��S ���gF���j�ܦ4�tm�_�.u�G�./
��
3)nw(��e�%cm�%�����$\�h^h9��`J���*v�~��57���]cW�}��e�=��#�������Sf oY���а���}p��ZI Oa����To��R9��B4R!�]h	.<)��qJ�o��s�G�,f@e��~��enJ�b@ �����|
=:㈰��-����z]�hD�?�9e���r�I���nL�p�]�G@���6Y��*!+�@�e�ȼD��U� n��{]�9����$�S[n|%�aV2��d
@��+q������Zo�z@���4�/\�ʳ���B;ڭ���]��@v8�K))Nl�k����ZZbf��4��V��_���qW��0m�Oj[�����Y2\QW$��	VP-�M�W�����lM���9�DuY�u���c��g�ѪǼ��?�����q	�L��V���V�á����u'|�t%�ÁYrP�t$}��U��X'b���Ɩ�d %���Z��3��D<���t�Y����\Z�ʋ�Z�=p2�\��1��m�6j�SXh��}h���)�CF�Tp���C1(9~"a���|P�#�TlFď#��)�}�up#�X��=	�C��Q��*ĸ����v(�{Bf�Ě�A�Rp1�":H`I�����Z8��_<�#Y�����3�L� `婢��W9b��}�����h�o��ƐÐ1�X��������| g�[q����;�o�14�X)YyL4�N��|�NՃ�s�:��f��S�]�=^T�ՋKםJLd�ǣ�^T�D "����|z��O���@a4�v��� <����~�a�hްO�d(n�Dʒ����P�����L8Sb�F�J�Ҷ�[������FzE[�Ш��*x�Ex&�s���j�IE"�H�\V����Һvod!ȸ3p�c��R�;G ��6p�7�Jn>K�p?�"��r�K�[9I��I8�u�a�1��N~`_I�z �z����P^�����v=��#��{.X�吜6x��r$��A��wND�{�dnS��� ӱ�!����į�����n��z�c���P[����S�ئ�Pe+Gy�~�}5I&���2$�=����Y����%r�h?��I�vphS�M�d$�&�:Ƶ�����cBщ����֒��j�J<�>�:��'ȃK� �H��<��S�ؾ��]��Mn���<���C���:Q�W��	����W��9�������I�g�[d]��R�ϻj��DK�)�]��誵N��;_��.�,x�p�Y��xT��ܐ� �C�*�\j����`b�O$�0�#���Z�J��~-V?�0��w}��i�����%q&_9�vZx�]�+�^f�'>-_��}�0,�j3�A�0���7Ki[A%��`�m�rL�0��TL�[/h�K=J�7~�f�4FJ�!��Ũ�UB��=�1EYDc�RXE��D�к��}�p�ȯ���N�̵q� :Q��큣5���Z�",���$����*�����6�x*��}NQ�����0�h��,��ޕ (��p���,�
�5�3��N:�����nE ;Y� �|�������4��`���!�-*��J��߂S��T?̼`�~gi� ��x�/��"�����
��ǳ�fK�ی�K)��#O$�b�F�V��ƈ'��ث���X�E`;�S6Av2葺� �~X��YR��,������Z��o=Q$�V%"�J�I��}��nb��\��Q��g�mm��Չ������B���-[�i�I	խ�7n=������y̥�[��>NC)`=5��ߍMU�4=��8�"\���=�����@���Tp��J�s�:g�e���v6�;�P{��ӷ��4&�aH�/Ԅ�PLq	�a*��s�l���S,Ζ��_�+z4N�,��٨xPB94�[${N�\B�U� �V��(�Ѵ��~3X�L� .�X5�4;�CK ��lه�]9Y~���$�3���hfn1]�gmw[��uµ���&����h���D�.[��1oe�K�������]�]�x��1rp��%���["nJ O"[�6�j��(��3HV����eG�|��� �F[�(����yM�������������͕��Mf�@���~�G�Չ�`5R����M����{�э�w�I:&W�[��.�؇�5�% �U���+��b�����6t����4<�,ܘm�M(�b��{p�Y w�Z�O ?�c�=B���&�<`Ӌ�4e��w�dc�l�4I�_l*=�M�F���Xs*��oZp�x�q�N���̈́t��V��B���v��6�m�_��篯E��B���r���ύ��FF�r��w�w��'(lTq�v�2�F�O*��a�ȡv"yhy�g!v�X�Z�nY�8���F��d�ĩq�/�8
�}��5�a )e{�;��,�'��������>6n�D�{�xs�W!M�4��bf�Z#�����z�"�2̒&�H����+_�J������ U����%��g�:̒]�$�-(iJ�*q�7|T��0l�(RA�@�vl�.��==��ۻe5��0�Z��H_ 
Fq�t�V� ��%'��{����^��Ң*���0mx����O3�jg�UTv��V�a��-jO�S����;@̻7
2!��5J.ͨ"��	N�O����Uh����O1�]��H��]��]q�o�$K�
��ن�X�̿����&�o�}����2�jg�#�6��L{�_Wtc�r1�Qz���Y�5p�\� �;E|)�Se��h��ҽT�RS��@����ki���%n��ٵ=m��� �̓��&e����i�?0��V��yPY�� ��v҃rѨe�ہ�:4t�?_��
J��@�q�Yx��pτk<iç�6�j
�Rgrt:��>�߬y
ѭ��nz���(�l�l,�6rN=�Nf�	ZAQ��-�´�X�R��99[���\P˖-gf��'ѕ�5`�A�k^[�>r�N�gH��); ߚ�H0��`W�3�{&�3H�-s	�p�pB��H��Y�;X������������LR�/�,U�h	�1��Vl��"��,�q�(���la��=ed;��������XG2���J����=��ʎ��	��h>u�颬�Y��>��/�|�[�!��@ͳޝ>�A;� ��$� �C�q��k������a�"(�ע�m�K=ᖸa=�|��ῖp���h�3�+��9��I��=�%?p=D?�
�3^�}^��b��8<��IY�Y�,Y��pM@�� ��J,���1k��Wq��eET��+�><�A�X��]چ��A�l�P7_���	�v2�s�-����	b>a��+�6g���EИh���f����:�nU�Ѯ�z4��GD}1]�:����~	��θw����tA8rB�(�G�>�K(�7L�/��u����ȿ��~�X��e�21&�����f��B�?x���,�ׅ4b� ��^�\^zc}�nQF�5Fi^�z��iY����D�����ޔ�ڹ��<C�ƣ��iwL!� Kg;�}��bܐfVo�ߚ�9eDw��T폻�2�� �_�K��H������E4��_l��q\x��e�W�t?yd6�>��[^An�̅q�﫨>Sδ�O�fO����*X�f�3h����?}unMUj��xUp��'p� +Q�2�@	�+IK^ZW��t.Q��HÉ4cQ�3��x��2�=m��ʬ�����s����i2>������n��!~��).`Y<�wKy��1�͐�O��_�z���l�A�Dq8Ek�694�b���)�� ��b1M&a�M�NJd�Y�B4<�s:}�X_6

���8ٱl���ܡ�GH�7f�°�T1G��:�dcu����K��b4J�95�J`��64�'.����@���� !�ɐJC��!����g���`cj�H���&Kf�7�_kZ�@�<��� �f�`1�Z>==� Xm�PST��e�?v��>'НƐL��x_���RǵU��͇��y�D���*Z!Xw�
) �Uj��͟���Bz��sSu�1�J�e�:�8�`f=v.w�G��m ��&���2���Э,A�G��v:1ݠ��`�s��k�Aj��Oy�W�@����ʅ`8	�vO��������k�M^����5j䙟8�$�����l^C��LN�hk���bV�gD�Zڙ�U�{Y��H�|��A{y��;,�!�߲a�u=�^k�1?��!r\���	o�1U��퉭�Mr�-y�.AKM_�r�/�2�r�d°n1����䱤�ɵi�E�]pF���h�S��+�T@�jI�y�-[��`�\=$���5w��l����e�W�������t�Vdq|��M��s��r�s�����ZC�}W*s��$�AS�T'@�B��Q-pf��R��ېT��l�z��]��3�^�_iz�f�y[8�Z+-b���x�?ne�_��D�4\�̍!*]*i�18�g�N�7n�n���Ք�D
U���nf,��<��M���z/&,τ�&���Z���Vn�_(�;O3P���dIb�zQ�c�_F��R��/4a^�9��xI�����#�~XD����yT+]M��/l�,���٘�vc�$k�v�T�|g��FQ�I��b��fs��\r�� 0��@��
	�>o`}�prL�������#�8�?Y��.�O�O�Qi'݀y�|0�p���*���bC���h���ߟ�@��@�̕�y�J��n�c?��q��O�U~�,f4w�Ur�"�b�V�z/��pW�cy�2f8I�V�Н���|[����XoC�Φ��)�HfH��o pd�ɟޒRNuyB�%`[��q/KnG��-c��W7I~tPTWa�"�l�.�,��RR�^V�7�k5^N��u�S������(AE���TټސH��gLM@�[�;?�s;T9ս6'Fp~�6�(*e�.|!���:�����Ɵ��w0��~fm�a]�/mŞ�^����څ��Ų���A>g�c<0~^���\����:���r�6�G~�js���F;���,������?^�L��v,�5Un�d�Y�c�sIߒ�>dyS�)9++:��P�Q�Bq0�PE��Zl�DU;)�L�x��=3a�(������5�߉��.�"��&���n�$v��Pen��+ɯ�S�eop9Z���-��m��QؑA��q��8$�[fa�e�bӶ#u&��t�? ��5���z��y���pa]�rqL88���<UIB����
�zxCt���7�����X͜E��^��[Q��:�&Psd1�%<�BVb�嗱~�:58z���r�>����µ�[f�5�Hp ��w���������B��e�Z�ݵ��ӆ�C����N�GSֆ�����L2��p6�dM�O�N>'tq��,|��m>����x����&;��1c|`O�Am��(7�<*����II�t�vbwib�1^a�:��fC���Tq@L����D�T�|��K�̝E��v�!�K<G�!@�T�����m`�p|�t�d�[���Ko[��*���mU��`(a\�kOx#!8Ok�����!k֡�j�ڷ����ME��}ss*T#���M�6hć?��ǿ۾|.Q�"K�E��yQ;�qb$�����	���v
�z�����Y�T��+#ں�(*�p��)z��F�(w-�N��\����g�Ք��0�ë'[S!��Z��[��p/���6��v��zzL��-+|�� ʑYm���E�oJvhjY�%.4�VHqý�[GЕ�
q1)�Oh���7����%O@��҄.����+�W->
t9Օ���T�}��|	� ӧ]��QN��۪rKH���N��O����*�H��s��m��Ǫ�!�DΫU�
��n7�)O�(W��g &j�m5S�q*�)t&���E�_�1:XZp�F4j?�w+�/�
M��͒�[f=p�.K�P��Kv�)%@12��L㊀�+7:�,W%�Z�:����Q}M�B���{"��dLSo���*ӄz�O�R�f.����J�*�d�>����o�i��yh\�~-�1�nd��O���K�K���� Ɨ��j���>\5�(=ȏ>���zP\B�������U3�,p6��n�b��qa��~��S����+Rkd���9�g]0͓�pI*�xGF6���ud<Y����C�NC�/U�[ُ.=D��E�4@�"u�1|���y���Ng䐸� �h!�G�u�Z��H��St�q���"V��p�x[��~�G��i|(��ӪS�־|�Y�?<�5 )�m.�����	����f͟���>`�A.e"�Ay!8v��;�c��E�Mx	oَ(grƇhl�?�b�f�ł����C��
>���CP���U,:y�ET����3p��qޭ�J"_
��#��6m��X�l��q�>_Qō����W,����k }�N3�h_������a�;�%��i�c�cH���Gb�M�w�����Z�kq�9YO�\�u;>�D��=�W���/�/��m����ˌ�®1�c�Lj��b�r˘�U���W{x�S��
n|�2��t�(���ɢ�9BL=�=�m)����t��;#�[��7T�p�z�Ę�/���Ҋ�{���;�8;8-ԙz,���Z�lKg���V�o#����U�ևD:\�Qzm��j(�:Ī�����j�)�����)�	�z��7˭�_E��p����|`��f{��,����R��[?����@��C]G-m��>�cBo�OJʏ�X�;�Њ�D�������_�~��-�~�ܠJq��D�d���Ŵ����;�"�I���QG%M� � =E���SA��[���-�����te"�L��9�$i��^+��Xvr��5��h�DpE����;�<�*�k�́�~a%�3����r��^q.������TʟƇ�kˇ��;�ebQ n�G~t°�@�,&���}��g[*�:��e-�tF��^��x����L��)�@�� �-AeՎ�Vr@G��= t�Z3��5���
�B�����׳���O^���«@�LӋ�R
A�C�^r�|�Ki�(QpP_xgw'1�`�
�z���6q�c�������T���V���*�7��i�H'c�;C��d����f���nhE�)&.Ϝ2j�����X�{8���T *�#�T�6�����Ջ�l�řs'Wd��9�@���!]� R��"m�g������#y���.G���r6��)�S���;�< ����N�H0;�d�:4w:�����o}�5U[Ծ�x�q��^�0��V�R^����[���NY �+�-�>i����(��i>Q9�Qv#�@͌h��rwC�&�� ,�Ę�f�fN���`��������N�@1�ߑi>��l��8ʣ�qFr��kR�p��0.�VR��⯳�jɘe�W��㼽	�ݍ��h���p߇����ND9,��d"�x��+��J�%��u*I+�����]����ۊ
�a��ɋT��� �a5�`���bJ%f)ώ�űMa�f��B��EZ�7�(�.0�gۯ���X9�����R��wF�ASA�EtQ�Y>b>p�f�_ګ|c3@� �3�h����vM�(߾p�E �����05a�P2��=4�Awg�^���4��K=K�D�,�uPKWZ(DY�8
�{Ђ����Ne��ڌ|��P؇I	�<O�_3?�J�S(֊{l���W�>��#,q}�2���-���,�G�^?�F�空�µ,-�� �� l�X3���ϵ��Q\��sw��`kT]����솗[']aH:�^�4"���
 �?kb굲��[����4y�i=F��A9�ýA�0q61ͬ�p���N?����t�U���i���O�|O ��j�*�>�7���+̃zb��^�\ �5h��G��*$q$��To�Θ�G8�����R)%�{�8_�y\^����jI��&@�����Gyh����
1*���vi[��Ԫ��Y��dj�����=`16d�H,�ǆ�Ǥd��n�j�'�*9�P��{�3�u�:@��(����J1�����u�����޶��i�/�p���iev%�U�ņKh���:Mk��`|_����5��3�]��@@	�i��?W*Z??NK�3gdޘ�pf#���#��������{��Ƈ��䀖7$S�U����0��
E7=ȕ��6z�]ϟ�3�=y�B��C�	K"@_w�>V�%�*AX���c_�Zыnj�Z-�IqNC�	[������W����+�ѷ!__2�&��f�� Z�/�Ưuk/@Nk�4n��bB�s�ʔc%�.xL��ʏe~���Jqo�fV�1reǞ�?�!��0����Nun�*�ɐ9���L`h����)�#�����wߞ�����@��k(6��`���Q%�svP���|i�5��%~N|fZ_g���\J�A5.$�T� ��f+���׫�x6D,n?6��D�X"h��=u��ܮZK�$kN3K|��� �z�o��~yUX��;���%+k���6m��+v�ё�I�azϋOs��t(-6@8�q����i�s^0�_m	:�W��u���{70���BM<��0$�8XW�p��B苰����]�ˊ�fx�b ˑ'���Ӫ6i>�z+��0	��{g��Ʃ�}�o[�h�ڜ�O��2h�٧�H9��"�s���T�n�'܁��Tn����$�-��xo�CZ����l��� j\�E����3�
��ڞC�_�Q
��XJ;�$�e�T0``^�<�ɍ�m�]�̮��Tm���H%�����X�G�T�0b�%��pC�Q��TD��9�n��l�����i9�$l��!z_�q�'c�V�#V�~���{	�(!�%��F��N_	i��4�.8��̀�	�I�������O�<�>����͇�~R��aA���R�>��`RxC��"kH Bɻ��I�XC<o���	�?���N�g���,�[�K�����>��@?�D[\6ėy,�D������!rVN�����5��8��vn�L�ਾB�b�=���{�5�՚��j���K�����rjQY>�J;T��T�~'�F�Fe,��]h����F/8��ҌӬz���;+eI�q�a��kL#w�����cw@k���uxi�oDG�.�-��#啀���?���ػ�sjQ�����u��B"�¦Q�k���4��-�x�CI`���؄Cr�U�����v��^a�mP�u�`��|<D!��i 7�>�6�����dUH����uJ�����.�Tɾ f������k�P,󸑕�P�����cI𐺁C?c��-/�5�I��]�����qKSI{�j�/�=�1���ĉ�y"��tz-?Ho���HV�s����;lt�k�N�9��CD�{�?f��z)e'ʆ� �&���w�{�m$ �H@'�牷/��C�8BE*�J��-)����o/����S������@Y����"� �k�t?�Jǚ�ɩ�eu1��c.�J{�<�3�� >���>*"5�J� �BKͽT�e˘����Z����Ys������vw�����"v��b��W��GD�L^Z�����0�3A4ϋ?\��g�C���eX }��zӓ�,P�Y��w�H+�RY�ٓ���������U vp�����N��@r�R���fmv��~�v���CA�׏ZET[O�l�8������ɦm7zՊ|x��=���xz#J�����h�t_����/^S�NS�XEqto�v�ؕb�v���-�u�̝�Y,�Oo�F+�Y
")V4�%��ז��=��}�@�w�2"�G��	S
�gL��n��@���O��I��^�!���@��}���������GT~ur���wG����c��[Qǅ��m/��͆��+�m#�E	�Z�H�}G��i+�;�� I����`o/i=�9��쐴�|�W^��������N�|�q�[i2af^۬+_�2m^۲᫶hzr|�`�~'ZWYn�֪('2#5`KKbL�V2oI�|�X��u�Ђ ��V���Ҽ���"�����3o��:-�wq�+(���\�"m��ٹ!�l|aOR$v}�G�52��Y1�䶠��{�����%}8��{Z:�ؑ�ܧMQ�4�D��ȑ�(��i�)��K#�B�
���[�V���vPD³��jRt����LX�/�E���T��@�T��ͻ�^����[7��kx�\�4���L�rXe��g� ��	���r�(��5?G��B5W�w�J��Z��>��{���܆4�͙�(�N=�;}C��C;�8Ƣ�'�o�'GIj�hTŮ��j���p��~2rX�/��h9Q�$9�~U�N!���?�¬|�P]!�̶��0�ʥ�`%˴���=
���cp�"��s����ؿ�L��|���31}Q�
��Fp~�6h�;�܇C��2�;
8Ph��nnOc�<�:y�͗�����{�&�4Z��/��ǃX%�"��IP4;�)i�RK��3��,��!���n<}��O��AI��N�Y���k wϱ[��P��l��{��T]�k����nw��<@b~��F<qcT^۩;��7�^��	CW#�Ȯ��ߥLC���7&���)c2��}m�k�Gb�Ϥ�[Sf̴�h�g�I�XhABR�i��ݳ�O�/�����ž��[n�~ֿ���-�I@����?Υe^�HߴB1}���z�$�gȲ���)������zff�����>���%�����}a�?�������XI�
���MMf�z�'�}�H[�_�v2��˥��{��2q��>ɶ���V�Ly���i�����`�����l����@k���� �Dt�mO����"��"�x!��uo���A,������jc��7?>����:fq��W�p@�(Z�H�;�,2i������ �\I�=O�F�J�xh��'Mhw�W��=���>`��"Yʨ�ub�]�	}�-w�_.H�Y������b���)�Ѷ���Y�*KG:9B����r�e3���%�m*��S�+�����`9Ř94l3Tpl�(�#B� ����p��D[0�IX+` �^�;1�'n۪Sv��&v�-i|��b%h�v�c/�0�wf�߱�U�ƿ�W�4��9�[e�x��fkѰ�B�<޹
<α�8�k��H�D&{�KWdx�0�2����OWXP�8>1~@єf�F́��ir�[�ǹ[q���=0�R�|���:�x���;CE��!7:^�M��q�!�"ՅLz�~v)|�vȤ��ED��������r���ĂV����.�H��'^�'�K��!�A���	8��~>�	av���J���PT�\f��*$.��!	0���1'������$���'��9���Xެ�DLm�9^�^�)"bC�X�G�!x%]��8w*��J���x�Y����L�z,J�[>r�s���S��[��9�� ������rS	�������}8�zQ�i��Q<��]�ê��*���#_p����e�ѫ¢�7ӕt�	ƍ@��]H6Qă|g�\��5���{�����M�<���`��L�7C0ӌ��D!ҐN�v���2��(������b4y�ْǬ�Ҵ �R��P�9�?���h�m2z>gL�������t�_lE)��=�o�[�}K֓(L@3<4S�8Q���DϞ�o�� ��r�l��(t��V�a�3dS���vxlFuP�.lЧd�v� �JF,�p�O��eL��&�:`��Z�*��&sU<Ye��=~p���l���M+K @�r����S�L)\X(��pS�0u�諥e�<%���l�N�BK�]ǆ�㵡�����h��!^�-�G4�����a�%� 7�!������H帱�T⯔̈́�^P�@c��ɯ{�܁�%�Xח8��7$�Ԍ���w��JVyr��Y�)v�yl~�M�%c�P���;�w�9��EV�b$��SSLVI��Ic�s<�(��E������"Ǻϴ	M`��G������,�a���W�᳄���}7%�q���D��{�ꅓ��ō�����Ud-����i�o
�(/*Ҿ0#���&�
T�I�#�A�ᑵ}��l,����m{Ü)�,�����^4͝�b�E�0'Fe���.�Fk��	���&�H���q�Q0��w%�A<�E��'�,��x?�����N�A��P��*̱%�v0��z��@:��e�[���/AP����&cf�����"�b,�o���%�*�im�%����-�L���B=�.;�y1Q�q=xÆh�]vd�6�"���T"��I��ꁠ��{ ���.����0�Uf�)+�W� 2���G��,7X�2���`��繳�F��5�����;�x  �ן�`�t�R�����aE�=�����%5�mg��m�Ĳ&h�^�{6�~�~�!Q��=�D��}�\-P����,0���do��*ÉAe<Q��̶��o<�jEF�e�-*.���NxC� ���	'v��O��D������S�Q��/���Ø���Z��K�=�/D��\�����oEw���D��5�<�c��ڬcz��s���A!6g`P�k���NW���n9���@;b)O@^�����r
��^`�J�2�2*7���hs�"�:��3q�d�(
^J>h�H�|����Ǐk�/����s�RC�bKw�,rԤ� �!V��y�G7��Ww���MΟ��B��M�x�'��+}U P<����S���9��/9�)F�P�?��g�ǒ�&E.	��k8j=OE�9�N��A1�ǟM���Q	���UP���E�Ce��P��FmQk��W�C�͛¬��|Re�A�/�Mj�cLd{Icp�Ar�>>�Q�D\�0��j)">���}�f�cր�>0Z�W��H�*�����	),��^(�8yZME��>�pe��V�t��;���nM�Mk�K^^�C��fɑ�vk�<@%-s��,�1U�Q��%jBpi���g?�l��1<]�92�蜊d�*'��M�!X���G"�EC�N�����CA�I�5,�V�@͔T�J����$΅?`UT"	���R_�Y��O��S�xp#�/�-�����O��U4c�����,A[W�:���z�t�Q�AO�
��{I
�-:�jM��ǃ՘H���%=�W@����B�Đ�"W��-���pD͐P�t;������o��U�VV���9� AP&a�5z�����in�].Jc�]��(g�I�x�46�~2��]v_z>%�z�P����r7�i���j��%A��$�pe�3����	q�����4���B���Wa��t4�|һ�u�$lm�?�Q�x�e�i*�G~f����w⥙8�����sD]wЩ��C�Bb͚V�=�T���]�+��H�uԨ������c�̼�_�4*��\������Ё
�]�D�4�rR��������~&}g�3G��������;����R��gq},�钺��dq���$O R}���ݱ�>�����I+F�~!x�0*�����G����G�GLN�/�'��/��/]�V�^�S/fv8����d0]~� CRS&�q���S�dgT�u�݀�e3BR�z�p��g�p���M����EsFc�#}B�_�,�x�:��A�P����ؖ R�-ѻN�P<�3�,Ћ��-�P�Y¿�dؐWʛ�G*RM���C�c^J߄��JY��E%�bA��g^"`�F���-/{@q4�n���{����&�-Si6u+�:<��nV���F͋�>�E_�T��_��	�5ߦėrY|�B*ziedӵw�ʙ�ש'I���j�?�휬ׁS����V$F9����Q�2�}Oq'Tf��z�~[�$l� G���H�3{"�!�O/�5.yEJ�p��� ���Ri��-��yD��w�4���^�a�X����Y�����Tz�$H��4�;�I�a|d�";�Z�,�Y[a�Bm�o]�Iu�-WQ�igZ��R��H��a���rA�gb(V8���H?Q	��-�d:އ�r�ٙq�f{�~2�*#��&��Oa��V&<�wWxqP�[��G�B�� &��������_	��!M{��1i+d�&Jd�/�Z��K��M�;V��X�N	y�`��IYõGj��B�
�4�4��n�A���8�}��*n�x0Z*�I�
	��_�U�dU�`���B�V/C�m��L�sS���(�]��Wv�X���&�R<��i!��p @	5���%y'%��C������ڍn*�rr�^~�\�g� �����GRjf ���{@���&8=B;]ꝓS�\�k����G�t���Ne��V�i�s�"��r��!Cy.�</����E艷}B�(�B孛[���p��_L[@m��5�C,f��,�����;m��êiT�R������kE����Б#t�A��J7{��)wͼ�]���wܠ�� ��1�2F��p[����&�N��X���T-�&�2΃3�5/?��d ���}ɀ��]��Q��1�Bd���A�׃�Fx徭��,���E���q>Dצ"z|b���J�6�����@��!�Ogr�9.�ڬ�'L�=�Q���I�	G��Ъ޲���������&{~�MTWWAe�ݍqA	n��a�a UV��	��n�CSqmP&��T7 b����"����U��{f���M�Aa?��F֝����?{M��\�9qA�)�c���H'��\֬��K�[��S���0�*��z1��b<��n��)��<)��l����5
����<�;�V=}��(;����W//��02���|����b�h��<�6z!Ǹ�<�`���������7�����Ġ��A�"�qm17�1u��_mq"qk,8���!�6���̊��(;o����Z)��YT{�Q0�x�V�8�4�*��V���ku��ݑ�cN�v��[�n�b��2Z��GZK�4�\�i��r
�����(���G|*��ӟ����<MO�\'�1�V����,����! <N�_����LS��at"�փ�~R+}�pf�	�95�b�.�]�?�9�Y�hl��	R[��u�2Dء]���e�+���Ƶ���oa�]:܍��b��zݸf��h�o�g���B��c������F��]i2���*s�2K�EBO�x%��d~-J�؅��M�NJ���+Ɗ����<�`�w:m�s���M>�h�\�|3��S�f�nFݻ�X���)�k	�&p�^�3�� x�QK�1&E 3� �LB|�x�v� ��Y���z{8S*�԰,� ��<�	U�'�ZN�@���*����O$��J��{����A=i{��ALt�����7;!?<����>��
`)��Ѹ�{��[}xs�4�,O�G}�6�g�R3�֤)��0��B��q�У����NQ)ez���^ ��oՅ���}1��U2+���%v0��������e!��Ț��e�2�ҥs�w��JG�������_�-2�!��MP+^�3�[#ξh�)t
�<���.�؎�(y-�E+�}�#���kV���q���?�H� �L�*��u�)�$��J:����j�t-��sM#h����S�/�M�/�yNid%�6�x��;�q��JGܿD4U���)��u)��V�wou�� ���Kzӭ�Č�ؾSJ��<a��j�>�
�H����!2�g�$��fq���^�ˤ��߮��m[�WP��|�kQ���ͫ6�c�ɥ5qt�u�f�i�?3�ߊy1���r��%9bH�� ����&R�Þ�q}iZx���59�ǅ��s	�f���I���M����K�zE�
�A�^tת�h@G�HA�<�Ix� �;���H�U�G��$�
�\��
cz��`G���9p�P�
�5���v�6�G��AJs���'F⊳�'vV)%����~Z�����^� �.L�j?"��{%�M�����	n��T1��TVF7�Ν�
�+ �Z�Fr�p4W��ܑ�L�	ʿf�����+�E�������W_��sZ��ܝ����v}n�귄"��
z�R������!�������yA���$D���z�cw���3>�g�'p�mo�������e�n�S"��{e���D}�6)V&��18�cS�9��W�4���C�"���'���-��/�Ņ����&y��g����z��j���r;J�v{-�v'�2v����C���=ȗk}�TOEk!�.~z���6�ez�9w�k�W�a���x�E����v��B���a��&ޟ�!�eF���e��L��"�a?	���tb&��,��q��3�������j`~��O���M�	���:�N������o ֧+$֛o5��I�u-93^B��4a�R�ͼ�`j�Kp@� ��zeIRCc����wu*y.l��>�A�c��ΆM�����%&k1�� 7�wL�8�>��3Dǲ=j��!�k=�pȏ���[X�9��,y|`y�	Y}.[wAO��Rxd.�>a����"�m��Ӆ���;�%��+�� MF;���;�w�@��Sv2As�و�Y��墇�����Փ�H�Q��n���7������-)��p���Tb���K�����^�do�No�CQE&�+ҭ��Uub��k�V��a!�=�G�,j�3-�Z	��m����wM�Dm��n宧�@Z������?r�kc"�����_��s�����t�΢��C*T+8��*��)!�1+��O�(���ю��ė;���t^S�X��d���mt�Й�{�����s�/�����z�3��0�),G��l�y��!Ti�r�U@�_�k� �F�Kf����Teӳ=\;܌Z-w�"�U���}�X���wU��2.mD���@x&�p���zh��NV�n��Eh|�S!a��I�!>��t���mj �Q�^W��\`f�lm�=��ث͘�����uW�{�Cw����t@,�+ �H꠭V����x�i:(Z�O^֕����;�����ׯa�� *J�?����	��q���~�>'
��,y߁ͳ�l� �\R�h�q�3��3_�\]������+������6��L9\*H�������p������Ի�ƙp7����~���3����.�J|��DT4s�}	HM,YrN��%n�E�N��?
l�Kg��/�d��.�8��&lL�/l�+h�E�5�x����N��4U�[?�o�9�w�7h�U�Is�U�w�F�{�a1IS�U6!.4fۊ����v�Ygj����-�~Z��1r,~0��l]`Eh0nD�C����!�Gq�??�=ƾ^��J�XT�u�������u_�gB�$�I�C�%R�g�8���l2UG�Xk��h��u~��f�W��H��Dj�ý�J���^�3<zD���m���X��>�[��N8
z��$�A�� ��$�3��g�k��{pM��U�*�b����@�K.��e!��r�߅�t1�|/��$	g��
Y^�{R��f;=v�����Lm�|/�)q�uߑ�8?��멑��b�>s�^:��շ9I�-�1��>���R����Qd��@e3�_� r��e"V�wrQ�G�+�&�tn��k97��&�����E��h�8���N�N�gB��%t�43�;y�sJ�4�J=n�%&�����h��E	�����_�LR>Քw���ڂ��4`�s��A9h��"m?��?f�}�3�jnr7@1��v����j;�J���Z^�r]}\`���RLқ-�e�L&Ykt_��a[P��j�c;�"g�J��.Y��������!��w?�d#n��%�K��a{�
`�(Ǧ����\4��/�G�����xH�P��V��ot@>�
��"-�`�\R��ux^�ө�]��X��Z$��J�:��t�o�-�ߞ ��,)�a�xa7ާN �jb�r6+�+Q8	�Y�ێ^�Ը��bm�ٵ>Ƨ	�{�\��;��M�����F�U�s����_��e�-�O�ki���ԫ���8Q���A&S���>#W���� ;4N��#Y��	�H��7�-=1B�/��S�(��LT����%�z��Yn(�/��2(xM0�Yʘ�z����	�Z>*��vY)����_�+[;����A�6�{��q �:N�_X�m{/��k���/�I�M{C�T�
蒨
�^�,⃤�ʰ�V�9��?�+���yn����0�Fr�TH�
��#Ƿ���ܹZ�k�+*���9L!��v��s�D��u����o�4EU���5%���#�� ,dN:%�WV/��e��z��@���Q9${�9���(���x�'^����n-w̫�mG=���5������\�=��x�~����Lh㷘b�c֙���ݘ�U��䑅���>ۛ�z!��&�<]Lo���F�q>�"�ʯ^�����2�Ez����"�Ĕ(.�����o-q(T���W#���0�P=$�3K\z� �v)�Ҟe,h:-�o�j�R�/wǨ�L����T([�Uö|��{r�ɷ*���\���~�:'���(٠8��!q�36�ip�Zd˫��Ϡ�j��R�	_:�ћ�T���u�r�Զ0���<�=���MxF:W^؇R�3|��^�I�c��	�%�nG�������L��|�=�X�~����8��VA�[d�-Q���S�r/�D��E�h/�f�<2��Fc֊��-��f����[�?��;;9:�ZJՃ��)�;�g卵�������mȮ�t�Ӥ�i��M�O|��#Je�� [0��/�U�!�����n]��O��/�Gʇ���,��&��T�N�!�KPʳ�Љ#	H��@U*�*�A2��'S(0Wr��s��wZ�h8C8t����KF���A����2�'+��,���#�L�c1x�cw�t�������:��/�e�v�\��:}��mBM���2l��L*N��u0��h_aԩc<D�2 ��7�1���ڞ�=w���ɵI�U4ݫ$�05n���� i�D�sƄ���G�c Y0��"C���P��O�"����ժIC{'V+K��>�G�Vݢ(���>l�Đ��W�8\?��5R��Q�G�1�$�#(v�K=e�*gM\"j[�E�����$�>�Y
`HВ5����\Av�s�w\���Z�խ�m������A���(������[��o���z$�撃H�}�W�;=u�i��n��ȗ�W���,b���i,�������BOT��n<��*�F��J
��J�i���C��w6pi`���ѿ�ƀ���A㓩�x���ՆB�`F"��b ̚Q���%��G��	?���sv �
�Iҗ}���4�b ��B'��R&e0����\�@Z���뗛�Qا�L�x� |���ʸ:��*���[�B�??�����qȉ,&��x���|�W��1�!TOT��⩈���/
�
8��
R�6:X=����Ӧ��Z�>��&C�3���������N�GC�G�������L��c��w� ^\���D�tg��r�k���;�z� �a���A�xXdd�r�Q%�t�F6pe��>Te�?�X���|�4�[�1������d%��Z���R��uD��?ߘ�~Tw��m&Q�联�!�.�ِfkя��l��&�}	�� %&��P�rk�M����5�k��P�6o�?W����3�M4ڣ�N�:����d#LuS��=� �r�Qܕ�rKFR� iF�#�H�O�BV7_�ʕ��b��{/z�wʬV����;O|y��4IOv�w�z>�4�`Q��f��a�3n_/�]E�0�z���P<��bu�->�gZ�?z�3B�+Iv'�Ie~������}u��_T;�.��8#���:��o� ���{��7罍�#6�VQ_Bc�H�4Ĳ�N^ݚ�E둖�Qv_b��NJ�?}��6!��a��ZԑB�l6�/_ȳ�P��k��gT�~!!E��16d�;�=BR�~
j��/����xY��p+�Yp�E@Ҷʄ`��)�d	р
���Յ�;P�x`���(MUs����K4nP Gi�-�{W�]�Ҁ%��߸� ҉/��)f�$B��i)��`�*KVTt@O��uؐȾm�����&s��^�¼m議ïc�P��k<勌�NUo�����p��]���16}�����G��'�;k]h;�k�|/�Mů��S>����v��מk^��<$�{� �Y�5ݗ/_��{+�ro��ŕ�~�nCS%�4`�M�n�U�d-a!�_��R��ē�����H��緻 kD��0��>~�7��e�$�=J�p�G�
'� ����az�D�6l6gA��i�4��bHN�R��ru-@���pm�E��M�1�{ըAW��Gq����H�U��ݤ��3G��ˬ�T�N�1݇��ӑn�Hg��ɉ����UeFH�^t/�ʂ>�`I4yV}������p���4����)�#���r��u��u��F���Y����.�"�e#{�h����U�lo�]�|�yi�T�>���G� zU�:�\ ��	T��ؕ��E�%�ca���j�8����S��ޣ�N�M�7iA©���K�d�<LX�</!OB���:�f&ў���O��}��l4]Z$�re�+��S�o�ͤ����?�aY~`x�������= Li�G�Ћ�!s�K���R�s�6C�<��q9|����?�g}��?L�:�.h�c��'�?!��<�ϰ�j�z���헡��:�Ns���K���,�R����C_�ռ� �s��r��c0�r����rq�Z�Ţ��/@%��K���f�5췜����m�hE1��3b7NU�~;11T����.�煑����(1ר��7+*S��k����T"���ܛ^_92�:������R��)<������?���-I�`�Y��f�W6�G�!-6�����VJ�aVo�z�W�Ͽ?��Y�PlSñ�#� �x���|3���<�uh�eI�?̧�k�=�Y
!����ʣ�Iu�F�Ki��#t>&±�$J�'�
�����m�� pE��5���rC�|ra�| zp��O���ju���z7(�i4�=/c��{w
������%��P�n���`��o3g�j�D�Rj�rߗ@�<֏U�FN�z/��kk��@Т9�F���n�(�CK!�S��Y�?���i/�DM����� ��Y�Q�8�.>.�|�-��k\=�� �)t�0��;n�RQp�L��T��ǉ��cU���������'F��7tsD�,rF;�'�ݽE(5�X��g��;�(��euw���̍2�(�Bm�e=�[R�������>��x��)��T�B,_QJq���S��s��a�}!��U E�a���g*l~��aY�;s�Р-�޴��,�A?
���k��*�L���b��֛N��ǯ¯���M7��'d�Cܿ�+�1��v�s
��e������5�`B%�{�$8��s\�ɵŦ���Z~.�
�?����}�Z
������XZ��*q�pi�}�H����.@yU�"�����A�B񣖂y0T?�܈���� +�IZS��q��'ʚ��ɝ�Ȧ`L�NKW��. /�ま@�)�.36������<
�@�"dՁ��Y��=�V���Q=�@�̈��Pԁ�)ub���c"��^��b�q��/��=��`�7Ou,g����O��wO�7!���O*vr��>	H>C�Q'���\}��C��śn+�a��@ 2p<���;�= �kQ�b�^su��_;�jC���D&B���8�M�s6�g���3�sSU@4F\��8����ii�%B@�&w�
Y�U�Jc�_�?j:�(�c�bf�tf���6�`L�VA���[} ;��w��Mɥ��a�k6��kWI��Y/�h�������߶^d�����jH%���(٣J�a	����@�MNe{{���4��4Y��W諦�C�9��Y�$O��-��N�� ��թmVr�z��cY
�|����5�4a��T�$4e��L���L~��}�]����aļ;4+}�ir�|�qܺ~�h�/D�D�q�'��h�S�85M�۸Ac]膖w�l>�9�1n�{m���{rc�"���'�9�ZV�?	��-[**�K�*�������ʦe�SB�}h�x&}��� SZ����k����l!��;��0:�0�
u{)6���iB;���˜ba1�_ʞ5�m�
<�aW+���i�G�=N�'2y�� ������`�'��B��j��FTڬj9����(�A�N�3~����M�I
yݭ����˹1WU�TԸQ��ڌ��(�GbV�L�V��>@�5���G�a�}݌�U��D��4���8��R�����84@��<2�}Hz� ���S5��,��L @H��82�X4��A����S�}A�i�}c�!���u9w�G��*::
֍�֩t�Z�?D�n%��;<�$"h�uS�}���D�J�u驉��A�)�u�.�c���YW����EMi�'��Z��Ə@*:ѲcJ���78�iƬ*۽DL�Dl�!z�a�Y�8��ޡ@O�Lw�bE��H!P�3����i!��V���]a�4�a6�|F`�ĶN��
 ���67A_>�7�W�n2:&�[>ʱ����@D/�;�����ÇFmǩ��9����=<�k1(@0�L1�^9`��zv�	U}�o���p��"7���e�|~����'�q������p�B�C~��B����{�j=�D��k0�x��3� �:D��)_�:r^�Y� -��s$b,�T�K=߻�KS�^����f������ܖ�=(I.�4߉��a��\�L�O���*H��7]rDk=KY���v�L��IZ>���'w,l���
	LX�d���6�-�B VD$?��Ƀ�F��}��D�X�j�`�F��,Yl/��-�'11߅���xC�R�k�k�:�=pf� ��m+��E�a57{���@WW�*W�6��C����j���k(KP��m+��u>4� ��Ơ��gBh��6H�%�uD��2����C {�0�H$�</������R�2�r0؈��e�Y����KױM��
H6D�K��DJ�z@I�6���,_H!��Ŵ�eo	p�t������5�=�q�������G���c&V�D�ƲůÌ��S>�µ$I>u5�;\��l����ڔ�'�r�Y�}�|���iPl�hXqu���D(�?@*� ��9���0�P����������~y_�$ab�����a��O��Hwk1w)F��!�Xs�X|� im�s�aK��|� �+�����(���u��p�;�S�k�B\�3���Q��������'n"��� ���r���W'��KO�?��$/��6B�s���u��q��=�5���"�#�� �W�Z�}�%`ri��e���{�=��#�R³�xm�R:ubT�����V����Μ1�F�����1��{6ax�����:�Y��� ~���g*���}be\B%��y��>�.zI}���TQ�r���b�[��"���� �K�[�m���#�e�(��n�s��^�r�u�*}��-���p��ge?��0���d�4�cS�mߙ�U�˂8K��ޕꛆ�?&�=\�Y-���&z�"�
�������~A���N*7�UM4���叉�[�D�`S\4����I可q��j��L�D*rHQ{��"���������O\�����N�I�6M[�1���C�������ݾE?y0���*D ������[�Q,��~^���r�����2�!�:#>�P�β>�w#�d%ݩU�g�C��0�0�z`&@�f��ݰ5べ}��l�4�������s#;Kv�ǳS�.��@��ApP���z�g�j	��s�U/@`磀J�����w�Hn�-H	�C�����}�5zАe�,�"�J*R�^ݿ�G�HEd'���I�o�r�H��F-� �+2���£6��)C�X �)���m��㝊Z�P��wS�[s���k�=�k{������R�M�&�gN�h�&j�A���O��l��%�%��]�
���@����]�`:[�t����)�@�"צKHվ��s+�����)���jv���*fx根�\�9�	>�WՉ���ioU5̛�L	����Z�c^[�i�ܿ2�׸����<���P�9�'�,�=A$��
�N�����ڛ'ӑ1������y�m���s.�@	�.%�>�<�Թ.Y�x`Ԗ�O��h��t�4t3�^��nh��ɘ��H/�`�_���Fͭ(�'�,��u��cU���#I���g@R#�O�L=P�a�#��4�A�m4���!����׆�>-��ToZ��E�
�6v�Z���2�{`��M��T�l�K#.@5��.Qv �0��ִ���'8�*k	{���cn���.�3���^9��{~$��<ecl
�҇,�9TR�]���2eR��W��`r�n�K/���R+MS��d�}�\1�>�R���w==T���H:�������Y�L��ۯ#j\����d.������=�WҼ*#>.�]�v���)}�n_�P����/s>�T��?)sh8`�u�D������Y����j �%I�y��&�/��C&�z[���N9���?@�m1�i�X:�.��7���X��	1 ���/o1Ӧ�F�w���>�Ml��j��k�zg�GM@����6(E���V���3Ns5�15�9V�7;�P;�Y"��o�秚y"5���b�.�-"[7z���}aQN�ꢢb�\� ɺ҉�"K�^�`�ϏC'��o<44'ԯ����K��ҷɶs5�5�N�S�R��
���߇�?�2o�.nQ����|�_���7�����+Eg�x��/��`��%)��N)���ʀWݰ"��L�Ԗ��9�2�i!}�'��Tk�i�h_�|xش._���|�>���e9�%�2�"�'�z�ɹ� e��.��Y3.%���`���rC�`W6�)���	h`I�b��2�j
\P9>P��,�a���s��V޳Y���aoG8ߜ�V�]�+j%r=Բ'�gDb���xi��Q��-
��M7ݙs�7�݆���9���s̜NƊ�wlJ�����׀`4�Bpe�5,��3��9n~�Z���� �wZ�|?Ƅ�%NLS��ɖ��X�kM�=�����umU6���u��z��+����N7�)�_EϜ4酫�U!���=ͺ/��m)O�]�� �=�N+�,,�4�Y�Zv"?�ܰD�n3XaJUJ&:�a��oZ^g������¢0Mp��0u�U�%�f�6��y�6$*!>5<-(Y9L!�n�p-Z�}�`Ĝ�z���o��~�Ob�8�`�@�>�Z�����u�!���#~�@������4�S��F�����,.r
�K5]^�^���g�$�@o�<�U���Ƣ�<SSZ��P5�t��"��E.�/�E�J�Eëv�����f��B�{��f�4���!�>�Vm�3=��Nm� Q'A��D�V�ހ~h85�p�n����$��]w`�hY,����pDR�j9����2G��5O�I(�W��z3����x�^Hv�%���V��J�ɭu��+oHգ��}��*@����D�5�Ҿ�������0�m��v��~�TI�k��iÿ�0$FO��&1��V����w˿2�k��l= �y����rg���< ��.�+���{*��EĠ�H�Ɔ�Ui�qr�ѬN]^i�B�t��͑,��Ke	]���������VbiV��W3	���A&M��&j&f� jֶKy$=�G��������=*�(P��>f���ꛐ(��X� �j>�jV�4��N��29Q���8�]�����u�ۄ7h"���xL܄Q�b̯��f44������&��k�E`Ւ����-<a�>:x;7��]����ǫ�Bk��B��G�q3Q��{M���*p�xlkD2nN';Ѹ�u���1����}�ͩ%j�;��3���l]>���-�ލ�y�7�Tľ��0դ�����\��XE�T 1��m�����/Z&[k�-����[�աwL!��@w;�!��t�Lě%Q�q��\�����˖F:kX�#H*ng1��Iw��^�\�����BWq�3S�Y\����S�J�jn�Qh{m�^�T�g�����t�)�~�,�R6RD��Z��E-Y��������\W�I��ӄ��X<��P���ٍ�&���UwnK}}i��jk�/��!l�#��6� ����Tg�Ez$U��E1�\�X42v44���Ğ��~��]�h]B?���NG��s����8�H��*%����.1���}A! �_�hd���� 6޹���	�����~�C�5P8hL?�� l(<g`����P��/a�6}S	��<jb����#���f�mI�Ô��/�,YEO� b��p���������']��(�W�rD��&~T�F=�0�f�.u\��nȈ;N��#(��n�̠ql�+�����0�e�uT�@=���Nf���tWF�JS q%�9R}�}���l�D�g�������/��/me1�{*0wa�z�J�Wdp̖�=S;	sd�ֽ�����ʪ
nE��*뗙����ք����`g2t^��״�� ����Q���;� ��Q�(�5��vİNWر�TB��TZ���i�)�\o�g��6~�Z� ���$s��C���@Ԓ���7Ѥ�l����9�߆�����N���?�n�E4ɀu�T���/!&3�ߡ���B�[8��c-\����ik���x����X�Uh��d_���N�P�D��QT���g��Y=�� �;3�r��[k%>����H2�?XE��"7PCQ�s�����DK�5 ��'>�Ds%G��b��k4!�⭉��&��>ĕh�-q$傻4:_|�WI�C�=�(&R��՜,��һ��T-��2J�R��X����M|���������7ǁ��d'Ϥx����`.��O.�i�d=z���<��xU�e�t�1�ڨ�����;�%�j��Ku)T�L�xʓ�����P�� �ml������p�Ͼ;�9ysf�����Ɵ�Zx#��0-��pj89��Z@SG.S�-�@�̫�M����/@��_�"��Q�p��p��X�ܯ�:�F�w��,�g��	od&:�p�ٴ#|;�K���X H.�%���~��<r���m��^���p��+}�*���>�-as���>��X�����;lD|�l84�dȇJy�v���<�� B��٭X;��?C�4��gZ���v�»����w����Ro�,�)`����k�Q	(�q�� Վ$�%Y��J�_=�5*}t����qjtV�\���}� �_�MPu;RV DCzU7�t�oL��u�m^����j��l��N����µ��D��.J��e���j�m�u=�ᬟnE��1\GD%��S���׍eNP)lUl;[mB�/n�Y!on���a�:'�孕��b�R���
1Y��eF�9p�?��Ҡ��h��k�E�����l�v�X5^�6��Arc�!�,X�X�ˈ߹���B����Ja�h�p�ڬ��bD����J��8C���j)B�u��'�4�Q�AN�sn�)�'�޲ϵ�}�N]�
��a�����5����c_���{������*꫎Ej�l�`u�l���7A0�a���'���I�dM ŷae�as,�j?񅋚|�E�A��6�:O�V�tͬ�>���/i��/S��|�3�:ga��'��>�y ��@����O3r��2�!��{���M�R��|'�Ewڃd��V���H�\���|:��/]S�&_At�h�77�q��K�C�8*#l�7  �bh0^��Q�v^p�aַ�
�>s�^�<,��}Usչ
��7	����0�RE�(6�H�ܺ�~ӫ�AO1�[�R[�b�6�j �;����'H�@��]�{.�o�)�Y�J�#ξ���U��তd-A��UZ�=�z�	:����n� 7"��a)׃٣�bg�7;��Y�@D*,@��:N�gTGJ��L��?�H�j�j�$(��
3ێO��m�;^�J�� 6� E�;dP��6���'��=��h��(Dy}+T�f�}�����ɢ5��!Wz͛���[pS32�t�*L�l�OW��l� HQ<�V���v���v(E0�H�}��ӏ�}A�l�/����7�]5 �B�B����\+���v�;:��f- ���2*>�����J�Ooaz�=�/~�'�$L�A��'��t�w��I|%9Oa2uj.o%��K�C~j�&5���䁋�$�W���Gw��m&*�M2+	2=���G]�n��q�MFsnt(�ДN5Dj��?I�I�����2*� �h�5*ۻܱ��`�;����u >�_� h�)��� aQyIR�$�aGx��´0�1����DFc #�IU�G�!GD�f�%��)y�י����;(7�H�棠hjA��4�	����+>m��T&����L4��V;֬�P)4##φW�+l��I/?��co����0-��Tr߱ P�DQ�i���)w���r��e�{�k7�~����	!�����ޱⵈ���ʔ֍/���ud�-��uըЀ��j�w3#~���|
Rۏ�s>�+ӧ��ٖ�:@D|z�.��B����6��R����@���o����e�����!^[��ӟ&�D>�X���7��!@�`L?3v�I�zU��t
q
S�:��u�
?�ڸ�v��a���PA�#{ZJ��+����Ud<��HI��.:%V��1���WX;]l�Å�*Yw���?��_\G�q^@�v���ĺ+�'W�� ,b�Id���Ƙn>E��Y��YP/�'���jG7DE�����ê��u���������<Ƨ&49\�r�J"�\;����w,XS�P�3u�a�l�W�������;��{W�!����r�i��g��ŝx�e�3�{��J�j�dzňN6�����)(��o��*����k�|HS���+�a�Ns��<(��Iؙ�ұu��@�&B
`��?�Ig��w�����9�YX�n4.�(�iT늟0����O��������e�����C�����g���4��.�f���F]{`)�o�Mz�(4�e�1`�#rA��qN��/V�?ܕ�	
L������a���5(a~��g��Q��ߵ
l���b+��7�����P�җ<IT��9�[�~麳e?�D����F�C�|z$�r����)\������X#+���z#u��c�)~�k����)�|�bڵj de�L�7�(B�%���;2��a�+W.��(F�A�'-�U])#^��~q��p�iXd%�p΍��\m�
��æ���J�6��K�m!wux���W}�(�s�?칦�)f>�<�ȋ�#6���1����+6��@I��f�� RBC� �Чe�s�jeEt��mΓ�ZV���vFؐ̍��w@8�WR�ez���w�����B`g#�g� 1%p!1jQ5�i�m�~����x����1
��˫|����t�{G�ɺ��z<�i��d��H��J�b�4B�8q9�#^J��N�=�^�l}��R�ά���E��Cj#�� F [<�LǏ�nS�3�L�����l��KG�ۘ�*�f����y�-T+�/��Zǽj�$����T�j�
�W���s^�&��h��;3b�'���g�����?b�9jbї�%{-��3{b=9�����Yt�o�nN�=�;�3A,H���)�H�#܁q��=��j]��o��xC�O�l��<"^����iK2P���o����.B�;�E��`ǀ�	���Np|�g�͡RZ��ګ�z�h>���%�Bv���E���<����ML>�GFJQ�(���P\Kd�ӕF��������+�]i����_��XZ�wA
�O�؞yX0��ӧ�S�}�nNC˧ݡ͒��*�i]U+6K<��RǬA���ǃ����[��ńN���V����F��p�����^j�Z���PQ!�l���k�D�n^l?����Q�DT�f��狋s�
'?���'�U��.4
Ǒ?�	�(�41���LB_Ph+�my�2~�e�j{�5��ꇒÈ����J��^'Ws�t���z)���~v��m���ල�	#�fv���	R� a�lC���|��B�Ě�EW����O*M[���N�u��U�	4/�|w��u���^����'�
f��U �5d���C	RY�oF�����(�Mm�9�u�rCH�a�+R}����|co�:�a������$����x&5���7�n�\�A��u�����'�@��~x� :�mݳG�] 5���Ղ�+� ��;����.�<�]�x�I�4�p� XB�v+��q���趷���e�[�c�\E�ϸJ2܏��-ݣ�T��F������2y,��Z
�P���`�,a�ppUF��*�,���29��x� �ތR,�]%}�q�Gp�h.�B�YI ��I6C4	��@p���(޳6�d�ww)�,��$�_�%
�r��W��<�jdP��"����>�2	����T`�s��_[�9���ݭ	{��$���zG�bBQ�=�ײ>d9��	_��'�i�� 4pF���.%�8"e�E�.}Y��*�|J��<1��W�����X�&�� #T�Fat[{��8�;Q��������|*$��cZ�W�o��l�TĐ�`k	g�[D Y��)	�d#�^��=r���W3A'"��� (�(+�[�V�$k)�|XKb�އ��X�q"�,e)3JI$�L :!��K�a���@�e?����siT�����k�l�ps%�B�Vث,�;����9~=z�pX��;W3�G��n:N$��h|��ďB+%{I��p��x��A�LC�#{Yo�g��EmJCYb�L�ͼh,3`D;�.�K�T��=��:������@�l����\ˌt��dB"�}��7}�������:6����b"�h9v�����9�
#�r�T9'�0�K�t.�o۠9=_/0�~VY.��4��[��Q.O���vSվn���W[Yȟi��(*v!��믉��ߕq2��{��ȡ�㉋Ց�xR)�/v����C).s��׺�?��[���ck?����z�^�hy�+���\v˱��al&��vq(FQ������4Q�Л�<u���ƨ�h8'!Ԗ��E^"t3FJ��x0tv�U���|kw�!O3�\k�d�9����	�T���n߶}����L�#@h2Έ�Ë ��贾���5=iw'V��p��Y2�@c���b�����13;9�����{T�2�rO�J*���}���Nj��U"���$u��>Wo9B���X��l�1���;Q*��y�e�䤵[b�Y�\M�Y;��B"��+��$�pw�L�̇41�7��-�@�����f���3f�_R�H�~�ڷ���A`^@ȣ:I$-�y�Š/��2�����d�GAPP22�k��*웖q��q�}�v5�x`"V��Uw$tdĴ��Qɧ�"F�o	� �����77���D-������4��,�汍K�c��1����o���Kk!��4�ي,K�"�ߒ5\�s;��Ŷu_�3 V������~��R��j����F+2��oEO�`O��Ư��-�2��G�-�#0�N�~�ŊMҋ���q��,��`߬V PP���v_��楴���?��:�S��0y����.�s�t��l,��XC�O��,V��_U�bq����pf�V9$S���b�G[%p*2e<�u��6�Nä) ? ��~7�^a�Ĝ^д@��S �W�j���+O�N;���Y�r7��g�o垙Q�SU6wL�^:�� �۞�%�|F0U#e*?S�T���?���л� ~�������VSi�1�$t��8׿t�W�_ԥ���)�wܣ�-f<���S'�T��0B���:�t�����MOv����T�Hҋ���j̏�W�2/���4,��{F-DڠLx���݅��G�f��xʎC 9F�p���vD�G~��.�P��Q�<��!���ϹPc�|p�_����1P�M^����iڧ�Tt:���>��P��z��;.�����O(���+]���N��Rɮـ�g�g�M#�Zh1��� ��u�ZUF� �k��bH�7�Z�Zd�w.�u�e��c�K��� jg{<,�E_hg�R���U����i�Z*K��uv��%4�_���"_̩\YR���+�d�vZ�]�bmI��4He��ܛ�鉈I�ٍ)jT��k����<�n�;tS��ot�%���cd�&�w��;4���ͤT:��G�j�.;C��;��(&��y87/�r6߼-g�6%�h���NAi���@+�E��u��j`��T�yDc3�E�H�ޞ6 ��j7��oQ���٘���eT$�E�~���#&�W����������1qY�jȇ�ovo���6F�C�g�[����X�X����냽n�_w p�N\HSѹ�l	�]p1&>��=�:pA2�W��GB�H����w��7q������y��# ȭ+e���Mh�s��{G�i
H�p��-�'Ǭ�)u��&��9Pq���^J�d����W�=�GEN�p��rJ')���n�H[�4�.j���+Ы9�a�J�@�2/CU_M5��o���U��$.%B�u��R�:�¾�]Ug���{��ͮ蕀�֬�Ǐ���ݑ���\�z�<�M�:n!�ܯ/yQmw.�ך���A��%`e(td�_4�4`�O�@KU%1�}�8�(ゐ����{��Q�ms�v%ӪW�L�2�o{w9z���ej�ב�3��Yx��]�@#���ɂ�$ h>~�J�A-�%EbU����צق�"3�����4D-Ì�VHH�;;u�l���j*:��
 )��M�e�&	��l�ϧ�oZ�#P9a��������?>I���ی-�q���I�YͰ��."��V���v>"(�X�<B�Vy�ƯT��>+��f6�����7��3@���<ۢ��'�R����|�آD+��<���	�w�ޠ�.zf�����r�8E��]?'ig`H[��$�y���[��#��O,����5�5��l�|} mcܿ����O^���q3i�����`���$��;����K�&r�|v���Q� \��OgH�P��p�G.���!p���Q�z�o=1B�R3��G��:�n�t�l�[��6���`��0o�� �Y1�
��J���@;
KF�oO��%{|g�2���,�X��ʂA'-
g���ef �e�p$M?�ZJ8D_q��%��rDի����N�q��	Yw"4�\�|TJ���D�O�9�o0j�+�}����i�i:�CY0X��1�^��G��J��W$Nċ�lĀL�e�*A���)uk�J��D�?��ٲu��)*tO�oU	ѧ�n)Ǘ�1����˭ݬ.q�5���J�j�`|��P]Q+%��Ǆ��&A�/@)�s-�%B��cxݵrm��l�T�$�1�,��6��ື�O�-v��-���(�E��H�3�*T���[�φ�5�
���e���W'FȎG>r�E�NV��L�:�*��<԰����.)��x)�C�sTU��k�fW�kg�)qO��r|�|�zf��:�,�7��!?myU��J7������v������Owk���y�G���#��k��a��F�y|3=����Z�z�Ӊ���a�C~�}`̍4DF��+~b�uV�g�c��C��S�X���01�=���B��y��*�i�_H�7���U�.�dܨ���yZ͠�3N��!����±��V&B��ݛ>��^�Z��ָ�`.�m��+��BMk�g�~J	�*5�*��!yD"K������g���\��M�VJ{ޞ#z%d��>��z?�p�������:2|�.W�?�L���*�����RHph#���,���K���42�| �q� ���-��:�,!��iTP|�1_gf`��6d͑�q���u�5�sY˸���S����!s�}D10T�[����ȷ�� ��aFPę:
u�W� C��:.��p�����M��Mc�� �Wڭ�R����VrS:���,x��e_�0:-@7[�֚��-�o����НO���E�
�hZsnr�P8�jE�Ey�.7l�����+�Q]c�������e�3O�������;JL����ס%�3brP�kOD���;��#�(�E��1(3���sms��&�%'��꺝yL(�V:s��ف�/'+j�.~�	!诨�|.�Zc}Dk�5tN�b(nVSeo_��d���o.2�KB���u�&���I��@+�G���8�*3$^��6��nB� �m?_�[/��
ë�m����X��=:�>�!"��;�Ӂ:>?��ۺ)�D��ݝ�+r�`��9��]�%�>*��j��o�����4��������`S�䃼0D`6��{������(��ۆ�v�_�������
v��vaÜ}�W7S�R���a��� )�`�38 2l����Q�>:������U�����i"!�Q��U$�ߊ��r���Iw+��?�����������kxqb���j;;T� ݾZ�&��c�zh|(�����`������]q��Q�u&;��R�{���Q�{���F�\MO� ���7Z���Y�9�|��F5�s,�Ώ��8t���q���\���E� �ܷ9�z<���<j���F�1�.��}qIbk)$I�P�BE&�\��h�w�&�v��h�v=U5����D$CL�P[�C�ϦaQ�-(#����ت�?A�e�Qq)�T�t_$�l���O�NǴa���'�<�.��hO���Dq�������g�WAG�	:��TK���;�H��:���g�}=�'�C�?S�,��ɟ���1�y�A�n���LɈ�����#�^CX��]�F�O	!'�1��͛���T�����q�)~o�F~lp9����A
ґ�݅����urT�=��@_Gx_��Kh��{����8s���	��j��T~cmv�nkǳ����>��bK^��tkȚM'om�osP���K��B�H2�+X� µ8���u��e1([~_� ��B����=��P��|�o�b; O���ݨ�ŵdԋu���1�/��>!|z���{�]�dOIK�6A�0�q��<6���ܐI!�&�f���Ƙ����Πa�0��urp��(^����I�Iu(�*� ���=�ܪoA�~�ȭ��0�����#��O�L���He�徏���p3�Y�-� ��Mͷy��H6�w�s�O~0t�-esR�7��
��d�nJ)#��~}�J�+��xG�$�բ�Ub������� �c�4����� �+�C��	�����Ž�>�m�Т��!������2��4L��ן�*b'X=�ɤHj�9*���~�J�luގy�5,�&27�F
��2B5�A�p|��#��Ѩ+a_b�l�z�匡���~��=�z��r�D�k�j1�����*��",�#����g�>��\#��'�����i�Q��)�n��RD�WL˻��R<�07CI�Zב���������V�����#4aUC F�
�b7瘰j=*> }�N�~`�ˑ����~ĵPWG� ��T��eȢ��ޕ�I��K=�k~��)0%��i$`���#l]j���f\�"B�BpF�3z;!K.(����.J�'Ҫc��R~��V���R1}q�G�'e�C�҃>�7����K��Ŵ���X��$wX=a~p}ɡr 9�D�C_n�I|g=X�5��a$��s���Ԍ���[�xE�c�����~7�\��{���0�3}���R���+٥��7}�X���_������wZЃ�� �G�=�'�Ug���|)�L���b��)��D�p�ӌm��jҡ�t�"0b���[e�cRU��s�f\��C*���|-����E�NZHȈ)&E��"�֨Fp�ï��ݞ؅��q�����{j�f��� ҕyI��,�Y��? �峒�r�a���븕��KR:��᩠r�WrK�.c���Z�adhp�	�4��	�㚶P�.H�B?���102���M�6!R�f�r�&`P��@4{�3�\mLv���&���ٟ�3���3�Pp��k-��璎�f�2�0 �i�s!_��7�x�#�~��e!/4�11&�
�p�t�n�CdCj0G����Q��e��M�e�P l��v�V>��Nv<5�u?�y�5j'0�#9�:V�圭!�����"��qh��u��)����C�}(�ҵ�;b!��*�x&�(s�d��;V~�a�)[T�f7�M	�m=h�i;d~s�N(�A,�f!��bD�W���N̄`�#Ds���V~�hӪώCG�'�W���4m��o������������?���)�v�
S}�mm� R�,*/��=�����[������91K�M3�RD�Ӂ�I.vr&��_�>q�|�T���5�u`C]Y����-�#v��j�����T`ʽu��D#җ8�]�nt���Nc������,GKN /�����K.V��r�4w~d�c�Χ�Q�XH!o[da���ҋ�q��M���s.�4���.Л�<�`����遼�f$}�����<9�uZ]�~�E��j:��krDZ�WqUX�Zk��xz:���@�CDMp�h�Q�|wQ�� c�I�'G�Z�7�	Y�¼�wJX�ǆ�{�w֐�#�)��QvU��W`�`�#0�sI�0�;��腤��_�2�T|M�(�T��f*��A�43W{ԭ��9�Z���v��=�g����ɓ�w�酺����V���8�)1�O0�!�b���>�iV}ldd�Cх�Ѕ6�իߦw�}�KAmì>�	�a�"�;�g�׾�J.��^���w"T+�l���AT��g�Э�z���3v�A���A�Y�V����6����D���ѶuJ#W����ề+ܧ�ٰ���H�œ�k\d����p��걐�AiEja��6KIN�f�Ľ����A�m�H��cR���e�&�9f<9��|�P�0cXSjN�*+����,lW��=�j�8tLa p��	�5��S�n-�/,�bw�f�Gk��)ʲ=L��g̍P9GX��96ta �yN�P�8������6�Jo�O�Ŋ���C�Mġ��N��qd}5Х��JC.��R�	�8�ZDa����c+e-(��d�}B*Y�ۉ�e&q�Bx��u"����-͛���,eȠ�
���FW��9�v[�Is����Í��y	�/�mPi��͠��IN֨�[�=$�@���6��%[q���`Ry�9n���H�b%�'���W�P{C+<�z�;�y����g�����>��ٚ�$榱�~,pJ�JR�0�X�5r��E��3I�ؒ9ғ��	8�ǈ_��o!���i����s�����C0Y�� Ó8��,��ת�]�cn��ml��p��J���|T&�"V�v6r���KЋI��f�]�l6���&O�SC��#:����۾fY̯յ�GR�/��ĕ@'�f�q�ٵ ���mۗ�P6�i�d�[�t�����'/�mP���V=/�-&�v����4Er>\ ����Z%t��P���O|F�����E�D�[��Q�Uk��bڮ�I�,��J��@�}a&=�v��8�4ͨ�N!Dd���D\":��Q���"�� ����ן�8����x�m�l��Lw��ܪ�[��6>6��$�@ �Ó(ٓ^z�V��M�- �y)�IF�#h��4QM�#o�G���c�#�t\��-Ƀ,�����j��v3�wYR��uW*ؕ���dǫ^��}��q��*�	��3�	�������x��sdy�Qt�� �6$n��/�f�s}aUr�ړ,�?ӳ��z�F|6�޹"��1����a�\B��ń� N�N�b��8���dg�I|u���vG�m��hF���{��;(-�`���h�b�ӵ��-�7�t���ˣ����C�n����}6^+>��k�U�{~�7��,3q.������Ц@Ke�{�>x/~���L'�ݹ%�S��wi[B5����f^֥3�>��F\�f��A����G�@�������Ǿ�A�ĝ�L��Q�1���ӆ���-R$�R�� (zE��/F3'�)�ǆ�J�&_b�c��;�����a��+*���$�����*E �4yL�q�;�+�N�L�l �u[�P�|3p��_[v qM�nlӞU����
?0�-vN��O� b����mI��gj��3��J�9�gM�Ѳ=�q wr�BJ��p�SpRm���J5k���IH$Q��2&�,j��]9O�kЪ�ޑ�&�m�=��$!��4_8*M��a�"����CG#�-����j��R�7VdE݉��Y?A�#I�~1w���깘�x�zC��!c�.��|�����ȑ��jaU²��ӑ��&��9�>n43wKal�"���|޴Mf0Qv��[��h�ѽ���x�Dy{V����w��(Ξ\q�܅u}���I�����ai�I�n��e��,*�h2�^I��gdീ�0�?b��5p��ʷ��}R�B2��A
�,�c<߰�62�~��ԫ�S�=�g-k���O�5i��j=d�fX���a�H�Ŝ���^����h�e3g�h]�s�Y,&}mh����ڞL`a���Ǣ��㺮?�B&���>s��*�&6b8q8,,�3���@v�� ��o��wڃ#�'�
/J1������+�ZD�G44`� x�-�N����m�i,��+Դ4B��ǌ�ߑ�lYR�?��GC�X:r�TW���<�Yi�@+����ш!fo�y����x�Cރ�E!��U8�Q?c�`��o���S�ټ�'tO��=�B��vˤY���moJņ���"lz��$�J��z���l��]9���	.�1ŀ���I�+�p��፿>���p�q��ǣ4X�̑���%��b�����Z3�����9���YW-}|�a;�X>���Ҿ�_��ĸ���ށ�é�Z�o=����e�p�{[��VQ4v��+��|Ah��-J����I����J��Z�Ly��Ss��n����>�N�_�?���9��E��Cm��m�,+���5�D�x��b�����ܥ8{������,�����������`���dH�m��uh�Ǵ�\�	�j�\���F+p59��"߅��w��zZ�/����B� V�x����b���Z�J}�~Bb�~���e�t��D�_ps����f��2u�ﾦ�gdu�a��%���Yj���j}�CK������wk�з�3ϖ,*1�SgqëE|��`�f�9I]�j2��V[��(���ry��т��^p��'���#Jwѝh��qzg����P��{r�8@CO������������T�O%�ug¢h�~ ��%�KV��9�����2���A��W�]�a�n,]�~M��$�A?̾k���7�f�,y���!@��]`* �m�K^�SX��R��uN5���_��[����}�|���ged�T���n���4_ڙ�fe�񔠸�����Q91۸�4��	1���^��|A�����[��y�&�'N �o�w9���b�K������F)�������wK0����vcj�o�3u�qȁvW@�R� ��%�����������ch��<�\��Z?Jm��ԓ^A�1g�lB�Í�f���� ��:0c]�XϦ{�f?�� -�8u��$�f��XD���y��L��r+��:Vvz�?f(�<�k}��* j�"�#��<"�wa�v�&4(��H���q;X���랩Կc�G��8�Ax�O o.�T��*�=J�HL���a�O��V���U�����-m��4��|��a2-����
0��^��.�2���d����n����Gˋ�Ŏ}�9�i�D)S�'�.��+a�8��g۸�)�,�3>��س��NM��� 6���E'"�����w�_�Dx�W��T'>�$4��dWA"�LL��ok?�WJ@����!������P���.Y���0�Ps����:K!�C�-�Ϸ��\� �b�ث�*�^��	�A-��Ο�iw��H��@�#�=� �D�#+� �fII�s6�A��������ʭ�����[z��WG/g7(�K9�7#8�N���$�Үm\G�T��k`1�7n���V�)����>�nߔR�<��R�>Ce譗��-X���뿚ս�ۈV:Lf���/�;y&v5(����~�A'C��|ƐP���C�P��6%}�JE�SǤ�'����F��jff��$�H�s�+�Ӽ�c��5?)a�/Q0�/9���[�B{b�Sqt�5��B����S�}�1� ��@�:5Xщ�?"��1�bos�^
���q������Fl���e�bF1�6G�H�+?-������YI�B����
�q'���J\��n�����*
����dH���Kg���-3����A{_��"m��oU7f���7�)��
(�n��&f��p�&C{@A�W��O�d�S�k�Bz��G��|M@�A�fj�[ůQ!��%��h�a��+#.��'��E���_ �[��5�]�3�xBT@��R�2��\2|������OGJ�0"�����֫#U�oZ�/=21���p�_ݰ�v�1JQb�m���j���9�c3.�9T�+�v���5�\k� y~z�ѱY>`���*+���/�*��H�w�zY�9���ųN�� �o��������5y����df�T��5��sE���E++�[D�d��������9"7�2{���Ƭ���$��F���	�4x�?� BTW�s��)!W�;?U��s�ݯ�WM )?^���J��0��xH@��^�d�3{�O�j��d�������kcU-�0�#�+�8{Y�	�e&�n�qik\�V�P9�i��� ��h=-�=��
�D�Y�g�z��cL���ឣ���o��2�gZ�P�`�jqg瓗��ix����W��I���"8���M���=��[�E���v�3�O�KC�z1TVU����t?��{g� q�h�w��|�a��x�'�:Z��A��x�5�9L]�T�`c�C�X�����q�k&�{8<��*�2��/h,y�c�<�H6��X���@�p&-�=+���76�%Bl�$9 .b5 9�Nk����u.���+^[���{h�|�4vaXr��MFYߏ���4~2�0�,�:1��n<L�.A����
eQ�֍&�b��$�`�1�����wKW�|����$��R7�d�#c��	�͍��.ǎm@իvW3��H��;1�R�>����z�qa0���B�n����C��uw��ҰlI㒭a�#g���=/ [��OF�ʧ��Z�j,�I�"�L�Q<������Tl����u���������������<��)�<g�;���2��H���֗'û��^9̇!\	��nY�7ڗJ�ʧg�
hb£x
,���T��I�G��+F�[�'��M��;R�	HdS�X�T:�X޺��#�=-3