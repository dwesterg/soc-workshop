��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�������{����(\A�+�^���CQG��%6(�l${��	�H-1�\���.q0e���pce����5y��%�6�!�70�EX,z�t6L���q
�f�vpz�f��Z��z�,:�.[�Ck��q�lw�7TD9���@���q4���
��%mN/P�.��)@�P��Z��UB�"��0�L7d����A��,^��}�I>p�O������4���e�%7&�g ���޴�k�W� �t6{�^�n��(?�@�8_B&����h]m9�M��a������?�O����*]�r|�֛��L�y��H��?��=g�}A8���Nʅ_�\�aj����E��>m���8v8���(~���7�a��-���Ox]2����%�:K����_kLDrI�>��R�:�߶��=hYN5F���*a(�r�����?�T���i�X�3��}k����*����B$s�W#GW���[�Х��ޱk����e2g8їw��g�Qt�4�n8����Kɑ��Bn�d�q�	��˻���v2�A��S :>eդAQg�~l)�	+&P�]�;V7�ւ�F�����& 9=A rڣ��Z���!�׾�A�\]>7X~��|ܼ�MvhQ���ƒ�"���Й��g�}�
��7�Z�ȵs����(c`}�`V`���vd�O���ƛ�5]�q�7+]�Cf0�����n�;:�B6��X��Q����ԎO&��5�}c�����q�G��
�Qjm���'��<�Nx�r�xՀ���|�N��9?A-@B��КPG��9�?��dRF�v��F�	!��X���P�Pt��Y��^���5��!q��p;�c<�-��[�!�f�������J0�s��Rk;�t���#��rcJ�nv7 �٤�Հ��a�v���J�-6��݄��Sz��3U����0#3x��`xK\s�I�������Q�oU��`�@�j0<e��'&�V��O��u$h��>�c��U`�p6>c��x�^��T#�,z	���F���i/-1WJm��Z~������ᦜX�b��PEQ\�]8����+SR��1�/�q�_�
�e�f�=k��,�u|UO�u�ok�D���)����w�i�	.�������K�`�a�j���j�=?�2�a\�(*<o���j���mWDKb��!�6vۖqD�n�.w;
�Uߒ�W�w�r���ǅӜRJ'�j�F,ZO<\�f�J�Ϟ��~]FL[�L�ϩ�^���Xx��7�O3*ٻ�D\�';_NPە��,Gh+8��%2�u��C�r%8�+G��E0��PZl�z1+X���Šqej޽5�����7S�y����<���b}"�L���/MN�o(p
�e[^��}w@�b�k)����i��4���}��1��'\Mj���t涚%�ki(9$�;T����][!��ġ\Q��j���@���ӡy�E��W��kH1���	���j��A�e��+:�m����H\o�Qx[m�/�tz�����t��+&V��BX���v���^�Q�'�rG��h�6šʳ�ӎ6�[�||�I!!q��_�W��v�`D�ȫ]�g*2Ǖ����~��xg:2N��A��@JBK�Ա�Sl��Z�ɬ�,�ˏ'5q�Xk��h�Qj�^�<^�{P ��3�����-Z~�a�4[�����oS@D��M��m�0�����YzI'y	���˼�w�hg� ��6l�	;:hH�zIn-����� �'+���V�y��<T~�|� ���9�~���MƲj�Q4*��p���v1�A�nY�}䫌��f�H��[Ұ*��5�6��
�]\?�+�d��W��a#~C��J��X|���菧H(�V��+h'�mߕs��i�o�	P�]6HL�G���/wb��(F2B%D����j�U~�"�b�ږ����}^(τ��-�B]-�i�i�(����%���q �d m6�9�-A�?Nn�om��;���˜$�p�f��8���\��	Q�;��5�_�����!^������Ԉ���������@� W�W�Ϝrfa*�Ec���=���Svohr���h��z@�'�v�Q����È��1���ů"�/=r`E�^"�������~6i�e�/��e	P!��B)\DȄ�d�^�[��"���:��K��qY��j�U|&�NԱ��w�Pk��2B���ױb�-yU�JWbaO���D�����:���;�s]�LN�%�2'��^��6"r��3�+��5������>�ňe\��j�zj�%:���NC���w�^��Вa0�S_;8��_��
������L(�:N����ah���|&��L�C�ʕ5��h=�9���-��'D�Bͩ�Ϟ���葘^L�Ab/���,\	1s��Q_<���7'_�1ֹf���/y�њ��9�Դ���. ���?����V�� �%��*����3���aT��^X�Ƿ�=F9�2���W�<�s`ūE ,�PVn�V������ŀF>vosk����5ʕ�����W���AJ���2�K.]�hК�H#ճ H7X�z���d���������K�9B�S-�R���j�t�[��e���{�]=#��gn�
�Q�/�����-�b~X\�j,��_�GYU���?�X�rt���E�y��8&��f��E�8�l(�B��"����o"�]��A	Z�b���K�X<QuX��i7j�ƛuK��J�OŬ�����q<�e�u���m���~���Ԏ�!��FO�� P��A} ���>ߣ��^�S��zU��b�%���A�ec�dF��d�py+�M?"�_�gWB���"b�[�ά�ۻ��y���:\��.d�����H�#%��{06�A���A�L&��!��ZjH^Qq���!'��>�?��=���(��#q
�����~��HMҷ�Bc�3������`m�t��#{�=E�/�4K�y��#�:�/��'��� ���-�3/�-�Z�jB�s��	����v�R
x�צ:��P_� ��8[��m�%>Ib|�ze�C	7��`U!p�������]��ۍЀ��=�ͱ5�G)(mL��Oa����o��'�I�ih-1G�������㾆�\B��X��!��p^4n�%Qg\�a���Rp��՚���\'<�23�������;�D�8��g.��0���o�u_G�}�6،A����i���I�+= �m9���h���*�:C��g\}�u�Y��&Iޖ�cq�ju��Q#>Nx�XΕR� a�u����`/e��< �2[l�	��jļ@��rz��y՛
�wQm9��g�����W�J~�$�+や�4�}W�E��ؓ�(ֿ�@b��1롄BCgPjc�u����c��ĄSг�5޾�{�v�,^d����D��0�ؤ�g�l?]��e���P�-�\?�=�mqx�W) \������L �O����(���VQ˜ނ�2�?~O�;F�t ^�OD<fo�x�|e���9n��a|�FexI�@�K�O�W�O�������,�<�uK3�)����b�إ�_@+���i�QW�D�H%�NK����($򿡪PgEv�WI��=a�K�
@1o���:�vi�E��p�Pj�P�9�9��������Ĭ���(�%����<,�d�r�_��M��L��ҿǁqX���,	NT؋����Y��n}V�L�yR7�>𰳮mw�Ӏ�
Uh�
t���o�vp�fz����P>��XWMD��}&��w��*Mu,W+
�)���4`s�Y8l�pV�z\�IF��Lw}F�&M
[�Qa� ��fd����+���p!�+��0�2���L\�4e�VJh����v�d3ӨD��y�A�	i�`�t#�4a	���F�s׶�"R��6����Y�z�|ӑڰ���DbuX��K�GjW�������]�Q�,0PK���B��"�����+�5��.��F7�r��1<��sƵ���������!\l����p0����*�UHI�H�q�Sr���\����9�����2��7����=��>�Q�jnXʼ�ƀ0�<��`��������Gz
��~��=q��N�^�"H��u���K�%YQ)�l�u+�	d���[7a,��Jf�획�d��q�Unw9D�e���&-�����0�����ňo�}�9�l�n�G��Ti��z��cE��젘7����J&'�]M� �<B��P����a��\8	q���6�o�[h��
4=��.	�sZ�E���TU���K�Y�y�m3�����Z�H`$=�����1���B��O�qo�}őeN�<�
��D�Py�n
ʾIC��ڬg����8K0��rd��n^��_C�HfL��X��� ���x5�Ĩk%�������{���̉��ّ�U�;I��+��b�`�o�]DK�26\��U��6�|�ۮ�U�ϙ�wf��"�Df�X�% @5S��UPU������5{!�-*��j��(D�����E���K�+˼]Phm����C�<*j�"C�6>	r�	���1��sE%��f�@�3��lY��:�D�0t�(���:��B�֒/��Γ���T���N��mS�n��;��خ��a�B�yj�q�����V�P�����,?�K$��ڈ����^�/
�	�x.�r��h�|�6[�����ʯ�y�rܚf�K���R��� ���L�
�q���R�s�D �1F�' �5�ֱ��v89]+W)nZлF4�5̈́Z�5��c����:7W��%�yNV�=P�� +�Ֆ-e��k�w����N�&���.��y��1_C��������;s�	��)�Ϧ��)SWQ�6��r2���b�z���H�}S�0�QR��D�1.mQ�Ai(8�}��lc����u�#���2�ڦ�C�A�m�\��._�I��a����.P�/�N,vC$�Au
Υ}%�^p����(W��rD�*QD�~,[�]�ղAE�@�$��|6{ſ�py榗ve�&.�ոw��@p��>��UѱX�oC$�_���'��n�"
��9���r>�k�) �~Ҟ�y�EC��Cɝ��8�l��D`i�10M�v/^+r������d�Gl1��@���i@Z�����.�t��7E�h�3���_[��� ]$����l,��~RG��
y����Nzl��W���v2��Eğ1�.t��|V�����W>L=iR��7�:�!�BH IBu~Dw�$��֠���|Љ[pF���.�:�G�ض�T�⎇ڇ�QG��Ӡ`�>4�&�Ly�5�u�A~3��f�ȇ�	Kq�(1�[�0=6Q�y6r>���s����y�r�L�y))�G���M�/�F1��Ia,�62�զ�����d�JT0�tm�lH�.z��j)���)�?ݍ�Cc�_��@t����J�����̕��@�]��]��s] !��R�%��>�`����I|�J�tɋ�I����n	�ݓ�^���T���"�L��k�����L'����8"x�LG�u;�oPV�����+����D��br���3�����VT�+G�MZ�%/k������.@�gV�a�gt�'p�Ԓ}beys�yiS{
��2/1��QX3(�Ŕ}�{(�0aB}�Ԫ�ҧu���z�`r�?b��[��U  o�@�s���R��p����*���2)���9"6���*ӣ�n��iu�o��z���C<�Rn-+\Q� H���d%��Ɯ�v˿�F�k~�d2M��b(�C���"S_������fx�~���A�Ƹ���BC�H���P�5��ƌk����8��K('��S���+gĊ����t�Ry��O��+�a'*��5��	����1oZ|tA�s�q�$@�Z���γy���k`��� /S�B(V��p�Zq�09Ȓ�dIg4[~c��"T[j��84t�yf�m����� ģvx�E�몮O��Z ���ވs�C�W���h{�-ovR$o���U1��Ӄ��>i
��/��7�i_��!�OZ¿���Z��-�¿�䥇�a�k�Ĳ��w<v���<�)*-�z<[1�/�4[�o?�:�CKps�U/����=|��T���P�J�Fz�Z�!<���\��b�m��.	tT�\a7��w`�5����;�,k@/�Mg�)N����齆"w�/V�v?d#�C�'�u�Y��RMτ˂O,0���Ք�
�V������b:�Xh H�&���C(t���9�hƟ��`S�N�̖�8��`�u�?�z��w�!e)Xp�j��{�9�1&kW\ʥ-��K�� -p_�UTT�NO8Z�촶@�QLS@���꨺ZM���Зܣ�x�]�6�go� s���U+�D�܎��V�Xl��z�u�J�'X������'�����$ÇtT�(��|Y���[Fָ7*��o��&*:�Y[Z
=*�� ]秀�J��
h�ݽ��Q���!/]�vM(A5��Tp��,l�c��ˬv��e�(e^����8�i~S��C�b,��X6qn��{©����Q����K�	k���I�
�v�\9PW�fgz[�q��}�ߺ�JAMO�t�8��M~@������lg�PGN�����13��կOG48:�㊘Pt���-a.h�ѹ]����v).�/�2���w|��\2#<Y������t.�O��5-�]{f�'j��BC ��Aݐ�עA�&͂��k`���睰�����i�WM��F��d��=�s�w��	��t�zA!��6�b �������UzZ�!x:ي~�?���/�ڌN� k�)OO00�5$|�l\�C� ^��q|�*����LB�l<��8�H�F!�\��J��]�sy�|m�[|^�Q����JDf!������Q��ҷ?������S��,
OW�5j�y�W#��؜��K)�i����4Nl�Ύ����Ob�33٩�[�} ��k�o98R����rpC�5'el�" cD�����Gg�7H��9+���*�����̓��r�^�`�RTD|m(&J�g��0V��j��eMX��a,5֞@/�ϑ��A��&F^�p!h�j`�*$�xAO�^��8�͐I��պ� 00��Ü��.`e.ǲ�}�����1GlN�e��_���V?�HTYa'�S�A���pe��O���գ�
�Y��3��^���)�"�^89e��z�
z!��������5�@"?�)]��J�wB�D�d��)�匁�xͶ|i�t�ƍ��]����L�t	����o��-�.]*�2�k�MMn� [HX�o��ɺ���@ۣ�l��'I}�����
��c�����"�u�~�5\�]���N���%R�y���||��9L4R�RMb���/㈳��ޅ��;���fҍuǷ������D��=7 D[9�)D�NA.��[�Y��	I���X4�P���ߤ���;1��z���)��F��5E13�\j�7;�k�SVV��G�/w�� %?�G���-^?�n!(\?���'}y�*���B��H�	Ӏ�{��2x�Y���q�p���U��������/��6��sQ�ݫ+��c��0��n��MaC�7��~�h���	y��Ŋ�<�D���ףM7�K����i�B�����0�?�_v�ef`�+�hLZ��e'��vOeϊl�]���ڑr�U��l&CY��c'U����z�d�GmZ`��g�2�$3��	��Fյ��m�赋�S�C*����GNG�,;{9g�PW�?�����b�a$���`��or;�U���dW�q�!���!����GsA�T���~�h7Ya�O%��2v�;�!τ�4G:���o���o�`k+芃�� �NXC�W:��a���ԏ�6\߫�#��/7�@6�o�c;-*�K�%�͉W�&ʮ�6�K��PtS��k�n�����w5�w�-�&�
8���j,�,�ﺻ鵨�8�G�J��2T;!��_c� S�@���6��(+�;�&��}F]�TL�}��M�UXN\���`��!J�%��� \	Y2�LͧEb-]���vȃȸ��f{�k2k)ܙ�\q�YLc�vJ�>y/m⊶K���������'j�h l�
��V�~��z}�_��kB1��(��q�
PG���3l���Q�Aa����UD+�qJ.G�0���RHN��+9^�|=�%w�P��v��_�$n�zc�I�ܕ <Q�8_�"3i�-�1��!�?�
v���Z���@)W�$/km)�����2w̸YY��~[P�_�&�&;���b��v>a�+0t�ה/gb1f����Qg�n����,��{��u��Ұ�LEË<X ����e]�Ž���E�$�r{܎ֻ����7��a��Ҧ*"��r���&�E�J�5��q�3���,*jh	=߇VxC�,\��Mcu@�,.� � yx#FU���*���I� ���zk��R�.��s��ʨ2q�0��y���l�6�In��G7aQ�P/�}��g9�G4d �����'�r�.A[�	ˮJ�g޵s���H�%b�4���3����x'��|�˶L�
e��m#�|l��=��f"�����!mEAf� 5��vsw��"W�F<4�O���$��|6�ٱRn�b1c�/^3d�*�e������QQ���ƛ"�s��hZTs8��;@�ɿ=\�.b����q��4G�/�ww �'�*�("�*��dR�wT.���.�\�x��է�ݏ�d�w7��1�@�k��&緾x(�:������'��Зfk��ml������e_)8Ϝ��� >H1>[.��d&� '��n9a_2g�g�.fO�c�m��È���g���1�z�0��FI`�-;��zQ��O�c�#Z$��P���5F|���{WR�7P�w�H��=@���;�δ���5%�d#�gm
���2Kq�6�.�p���3L�ʄi�0A���^6��B�\�ծ��]��dtP�Z�T����}E6��	U	>o��0A������o?�$���,Ub�46��͝8;� ���{�V���9x��A`��ڜ�.����9���g8�B�w
.�.�,o �u�u8"6��>��~0ƾX�3y�Y@`�.Ҧ\u&.�������yw8O��:̗>��`�(B�A� ��N[$ձ0�c�|�0'w��>�v7�-[��99qܨ�E�mҒ�fdDIͣ�"�5T���1C$U�ֽ ��;t4�r�����wOW��{2�,`b.m�dER\���F��N���i�#�Ԑ͑���bOX?�J�\�:0���m�	@�����Ѐ��_4��7�:�>*�M�:D��UƏl�H��I����S��|��}�'��ʃ�ٰ=���6�,��Z��ڱ�gp{k[�n�-��8I�S��(:��[W6�i�<xR/e��Y��=gK�9�T�U��?�������F�ht E!`��nE�����iaW�.jZTd��ۙs�gVy9:s�O(��e�W#@�V�I�A{�S�f����7W����w�Y=�o�o=L9,�ĞPLa$�*)֚�ַ��SQpy��ɂ���>:{��
��+\̰u����9�3�΂����d�ع�t�e��tנ��h=Δ�����S�ƺ��m�Sʚ+̽0�|�I	J�-m}�O;Z�z�,�g҂6��6;[t�z��)�T�h%�!��ʪ�;��t1��`2obe�{�C����#�6+�Q}߸u=ܲ��3���t}3�%��㙷�%!��V��h1��	r���o���o��}���<�j��7���35�G־�%Hy��y�'q�:g�e������3��'{�i|M.O�2(�o�$�d����侰,_0��G��_��pJE��r���6M�bW�p�t��9�%�*����~��e}��S�I�}?������o�@|k�]���B1_�K��A��h1���A���O�j/d� C#�BJu�{I��xRǾc #_:>�|١��8p�Ֆ2 hU)�t����I	ۥ�%��x��<$1 �� �f�.M(��U�|�K��b�0I3]�&�oD>u'�����'l[�R��U�s7cbwH/.<�@��(�ZD��Ļ�h|^�rG���a�SW�w<O92�7��M�]����ݷ�qB�7�V�S���I�;���~�d�����y I����� �Ȓ��:��Z�N?�Bt�<�%].���1�\�-5\ׄ�o�!o�n�W!�֐��^�٫�R�t%kF��뉾��$���O��̟f^�K��b��\�����?jZ�����S���n�"��C�b��X�xw�St�I��H>M�t��zk,�����iC1�As"�i����-�zɬG�^���V��Too�(�V�k�,%Ȉ���g��k�xZ}�H�麥a�����ي��@��P���+�����d��]����������gx�B�.U�t'N��f�Z�x�z@Z\�e�ܰUU�*)+{'�"m�W��-��<�l=(�}]Ժ��h�!� T���4�?���{��ށ�g�k�TP�Y�zt��G�땝�����!��p�n�/���i�M�>�.����#	�.K���Nxhe�T�.2~-��V�'A��wx`fK� Tao�	ح:}�"3�D�� m6���&h[������
�e���"n_��8^1x��PJZ�h� �3j�e쳍���yu�-�Qa��)�+SfD+{�i�X,�0Qw`��݈G0VM�����_f�tA��$6'^��I�� )�~.M58%
(�5#X�?�t���G\��n�ԝ(�O嫡��#Lm[-� =���c^�  �|��n˞�zk/s㒒�[�M9(�ֹ l�˰cs�Z���ߘ��8��C������Xg��KRb�Q�ZKB�6g�A��n8lXB����h�#f�}e13o���@�-�����OQ�V�����7Y��H).�lMY5eT��9�n����W��� ��Z�_�(��S��6uX���-<��V9��ՅɎ��9����vY�Yz6�s%Y=��s��]eZX�߾��"�9Ѧ��QU��8�(�6Zv�<c����aE4tkfU0��C��'�
E&��8�-��"�01�px��yw"����NemZ!j���ɛg�_����|�1ࣱ���l6Fig�_�8�������n���i"�� �}��;n
z����ۥ�4��L���
�J��TP���i�E�C����R��Of�䓞��jJ��V�ڇ�/��2C L��,�(h�*y�|^/e��1� �1��tmR�-�)�Z�D
�~�Cλ���Uܨ��G�_F����O�I�Y�f
REf�U���������dE�����A�,Ы�H���,��c�	�^gm�ۢ��E&����C*z����ޡ%[����[���y�NA`�鱽��#��ܑ�zLh�F�}R<⏿�	�G�y�=��ѭ��[�8��|&���=@��ڒ���r���z�g.y�B�}bdθ5[��G���b��ȟ��%��#����ʀ��8\�	��f�#��r8���0�ϿN8�*}�y����(%x�&�a�>L�e@��RS�2c�%:\C�Ǌ�V#�m���z����\�h(:�6����j
9��J���a�S�05���"�%�a�q��iܵ�-��I�4J;�!���}��؈�럢�}3����,��>�3nbB������}�t��b(l�>+�O$\��#��ōh/�n��	ɩJɞ}��Tv@i��?�s8-M3�!���8��i3Z��S_�^�����x��i����ިR�������$~����ᝧ�ݯ���Ǎ}(��c-��.\p������K��Ov����-�}�ֈ���O�jy)�XxϬ�\���7֠-�&�*gLh��d	ܵU��v�Df�����g�jˉ��<6t�@^�Z5�{�������A�$ġ��������ٚ�El���d�?�&�GV|�/�fG0ڑwt<w�9�	з��s����cͭ��iX��A�[ovl({B����1t��;
M�SL5ia��*ir�
8��#v!�_8�	�	P�l���[~���������y�C��i0�p��#��i2uc�Q���'�
$�(���ox���1Rꉴ�Ȉf��̙�*pC�!�$��
���q�5I���ᅡ�i2����ۊ� Qf���*�c�����A��2�::wFz@c�߇g?��l��OFp���;_?�0:�����o�������#��>e�Բ9=�P7���¹��5=p���}2ډq�{fZD���$��\#�r������0*%�a�b=�Eʑ����\����N�SR���]�1Z����lR�"�r�M��v��v=U,w���|��M�#pQKM.F��iql�43oP�� ���?�����W1!4�$"P�Ȩ���>˳2;nN��n��y^Y/G�T[<��O�G����[�;����n�t������;�����8�����(��Ohk��۶^p�g~BI&�^3����_��q� ��������b�u�a�պ&y�y�@@[��Է��-
�=p��PO��"�~��|�T "���>h�5�i��o����6aȩ�2_3���Qi�ZB��H�Nܲ�L�~~����|�u�_{+&����u ~.exzz��& �}���X?w3l�|���}0����<���r~��rG�
4��l��2��/qk���j��s�\l	���w�frru~G;]���pit��,ܘ�:H�6�Jj�0bYS�6�^G0U����%^�M��2*��~DĤ���[۟xs�Cʕߢ-pq���k�{��Z�#�v�"�y�~�t� 1\�� ���Q��'��JRV��!D�x%�Rh�j�]D��9W�Y�ҎX"I�.�?����Q����z���W��Q�l_p�k/R��X�L�z�\��Q�m�;�E6(��4���$T͇��:Y�o�d�x�W���T��#���� ��E���^:j����(���}/��w�?�ҷ;p9��ھ�\�9���^�l���2�
VxY�wa��Sl���9Aa�\�3�,�[��zg�3`�Aa�jUa��yW�:��Q\����le��m�y�j��m�I=YH�>���ю�)��x�oE����aSY�ӯ��A�$v�`��2z��xe)Ղ�Z'm֮|B#Sx+�*�Z�s�ܶ��<F7-b!l��v��'��ؿ; ��E۬>��	o�b��ݏ�T.�*5��,��O��Xu��L">J~��Ɠ�#�z�R�4���^���w���veZ�{}S�qk9�N��<O�)<y	�)V�`���b�Ӵ�J�'Y�V�/n�(���	7���V�����>��a�^i���ҏ��U�����n�������|���;���[��]��^��$�Dv,���~#�YCe�h"�z�;�<�qcL:f�#u9��Q��0�PY�Ǆ�#��U#
�;�M�	]j2�	�w��h�Y�b!���[G`��������K���=	�TQ�<�p�����ق����A � v�L̻�\�+黈T׼C ���/�3ܶ✆�s��'���ρ�i&8>�GCNc|����Zp8K"i�,�3r�u��闠�࿖&3�e��<����pº�@NFA���;o�Z@�x�X׀9Ƹ����ֽ�Ҥ�-��EsB�'�AMUD(~ӻ�Q���֦y9-�Y����
�v!)����xϠ����58e�,������G�>5����$\-������";!��$Μ8�`~���4:[�z���	y��&��Bֲ"<����S�E�q�Xd�,=D�t�sA���9�?�:��0�@�=��6��³�_�U���GF: UXk���U��ad0�Y(D�c�N��k�%�a���=qt��4����t�ë�1�"�E�N <�S�'2�Ҭ����GʤAL!L>������(P���u4�P���X�����i�3� y�!�$ժDA�ȗ�I�0K�2l2�,��Ka�m/�>Ҁ.��92�$5�K!o:�ul� �U�}��\�PD�A���q����½������^���L�?��p�T�z���x� ��_f�<��ldx�dc5��<)���#�B�������w8�;�4�eyL�'N,CĲ�`�ir`�d1�S�@As�r��MW� ��c�oNq[�I}�'�`塎�eih��u_����p8��sw��3v�C�[�~�K��f&ݲ�(kDh��Hf8�wHI25Պ�S����zA��M;�����hM�)h��������vz}tf�tS�_x��d�1��	^m+h�����~�LHC~E�W��g�QΆ�l�X>�O��to��	 �� ��LK���T�������nj-ԣ��ïw,wR������W��l:ӝN)�a��zl-�X�An�� u���VM\mnXF�3��܃T�C}J[��ҟV��TJ&:�*�N9���p���
T�v�^�V��'�V��aee=E���LBv���2]��Eկ*��K�|KZr'r|�T��4;��{ k�8�R�/�a����l���/s~�}�v��L?,-�����߿�We$0�=�M�0�����v죡����u&����py.��ο���炋�gcO���+m�a���  KǕK-�k���諆�@F��=��"i��ǄV7<S~�.��ҫ��ݖ{�.���ErQ@	�6�C����s��i��N��Dq��f{t��u���(d��%H�|y�ӹ��wr��J	$����n�$v[kxnqu/~�c����*j��le{@����Os�0!�F�P��U&��1؅������ς���D�H��l�6:�!��:�޵��˱zAggβ�ԩ�])���c(��xX�/��D� ��$א�f*��T�z[��,+�$�p=[�eD��<�&i�+@�Kz����!�۝+�-/Rut�\;�eս�C����K�����.�)��^`ӏb28�3/�~�W� �T-X�������ҕ��*W��G� D����L��W?���D%a%���/AN��H3>T6q�j�&gԂ8�RoN��&io2�AzA�f�ބc�����M���ZiB?n5�߫�+��Awm:�@�����]�b�n�q��z#�|�cw�<��a]�B�Mot[d���̄��N�'�ȹ "��qv���j%�����-�� �1Mgh����j���Azj2{� �-�����6�=7�P��-�*��#E���PX��⣎�V�@o��^��'���L~���M���q�[@�2	���(�LcZBy���hx[т�
 �o��V��X�ԧ�nU���e|����
ί|T����g|�ُS���B�\���x�_�0��{q�����T�ԯF���n�U�NF����idk�8����^����g5�l��)�`C�uka��i�h	+�W�w�|��K�l
�����rh	���f�����[p3��_:c�jv��Q�U73Rӑ}���w�X�\�S��]�F~��&����f3�Y�L��4��{�"�h��)a���ղ�W\02~׊h�Ho`L��q��>Rښ���Y�$�3��#[)g�1�9x�.�g�ZB+)�a6�P�����.h���ոb��n/8<��hV�/���m�+(��u����a�ޣ6�r�K�٢�I�O�$��P�wJ����.JP�ڂ���ڟ�?5�GVO��<��%���I�,�9g-��0�V�aK��k��Ƣ��!�O£���$��P��d�����"�v��Ms4(Y��5IW�B��F�$��R�W�CȜ �s�p1�{s�݁	�M�J�v��	h7JzH�/��O��a��E�Pk̫����ñ������d�y��)N��;CP�dY�D�1��\�&��h�j�G�5�7�bksp-�4��tY"��`U��V^�����=2�M�
B0�$���q5�]�b{��Z�uBG��2�r��̠��Ȱ�_�ٰ)��@��d�p?��vQ1���� �y=���*"M�+.+���U�mNU�����v�0e���f% ��5