��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V�WV��3`M�KS۝��5VWVr�ndh������*����㿣K�{b�Wh��g\��a��7����_^1/d8�cQW�*�����p��m1�]XxE%ƛOh�8��8r�0�n�uv\"���mת��Jh���`>�i�y*3i$���눮O'Y\�����������'�Ϣw��E�1��]�I85�%�(�r�H_�p'�s$��(�BF>1�μ8���`���O �m�f��S�6c���,�^�KH�`�����+6ƃ�.8��9�������x��P��/��)S���$����Q o�8�)>�Y���E΍nߕw�>WS�!Hc�}�T�EG�npk�&H*/�dr"���J�L���\V���d��F��}�E��D QC�e-��̌�bv�$9��i:���1D��轵$�4/(�UD�W����������ZQm��X�t��[c"���;���]%#��ƀ���Ũ����R��0����t�?�ѧ�P3[�5?m�uVO�E����q��q���z��-d�|�,}$afd�ER��{C�$T8d�5�Ae� �	�#�F�N(�������j�0�-)o���Vz��I�VD�Y�j�vb���^)V�����xsG~r�4�m�i_m�*T�p��se�HsK9�"n)�٪�9Ӹ�������L,�ތ�3�k�!�4�JͰ5)�����f�2���q�ꖡ��W���%�Vm3�	�rX�4��1���'R���#g����9!�o�ui�W����v���o��)�6�e&�;�J�tV��c+�j��wI G��=F-4T(,wI�ṱ$-k{�zU�ǏX/�e�[	�]w��,r&��ͣ�1��-G����<��(ZÙ	�ِ4i^�w�N;� 4��?���r��C���������HW1�y� )��	�gт�$7���
�L�O��%NN���Q<^/��#d��
Y%�F�-��(��(���d����4�n��Xᔨ�Qd�E����E��Y1�n��!g�u��F�B�N�WZ�o�F�VZ������⋭L�i�rw��Q���=I��"�6��V'!�`�a]�ӳ1%���R��[��)�^�o".u�(�~N'SU��]Y!�g!��Bb�0�S�&ϯ��0-�u�������J�A�[l��.H1���?�Ro�	O���:f��̝�ͺy��O�R�����G޹(��|�;A�"�1ܶyK+�@��z�s�g�;��S1�-U[N����*���О?�nVi�p��<� U�3�\��=r`+�2=����7���^��q���{[J�7�l��6N��_�2�~�`���uU[���+�������;�H��A%�ޗ�Z�������+��&��	��E�)�Bu�`�������&cR��
?j�%��IYt)P�O��?JPQէ�<�gE�r?�nv1K��mk^ی]��Y'X`ۈ׼PmM���"x�v�u��0e���|o�^|(���Y���{�?�&�����露��_���y�KBZ-)�<�w�X��q#R�]��$��W5�!J<�Q�P@��[�MJK�I�6n5�n���+V���5�9���W�6��=~x/e";6���m�vl���Tv�%��kt�'x���-�p��.�Ǻ{9��eE	N��n`��
Wj%��&a'��p.֥Y�k&��I�%oTFjM4.����߉s$�C���W�#�bG��+W�r�_Kf�Q��c`ܭY{���u�8�%�+����iX^��xC�z�{��H����������E�l@z����V=i� ���L�
���w�_�k�
�p�Lr�7�^X�G�U/m��֡�����-\>z�k��iԅ��Z�)�[$����Y�jj�F��wΒ���F�L�|4jZ�to�E(_���[�-�C��L8$A����߾6�usJ�/s�Ex�Ed���	�{�4S�dP�y`�/M(�%��Ǝ'�i� #�����rߤ.A��`�g�t�?E
��j
���t�P�n_�!@m*6�-�,칏��� z�Ф������/\���q��1����1UQпo�K��K�3�?{s��ϫ3�>A
�K���m�d�waz���.�Xt�g`�� ���H]�=��~��f�4zGk���R�^��?6e�#��쯳:����z�l����A.�]����M��� ��p�+��,���bԇ���څ]p���7�yʓCJ{����>ѭ|~�� {��/4���]t�(?�in��#GkFd}�Fd��tbjk�������$�Ś��������y�|�Pu4L<Q���������v��{ti><UZ��O��}����o�JL�ꂁ3���C~T&!\H�{
��2��7�ŌW^ΐ�̴�lg��S����h(Gg��>��nε�T��Ų��g�,}� �
AE��g�&>�7��c�gu�e�m�M&�Kw?m�onw�7aԇ����z��Z F�(X4�x��Yh�e*���*��!s<�֋���6]3�ئ��T>��yэ�j(���t�^mYG�&���䠑)��Q�Z�9�qdۗ<-9B��vV����Qq�wwׁX_��%ú�	������>��]�+��BTd��ے,���4�1�ow�s�F`1���M5RI�.���[���@ ���r,�(X�����ѭ�y����no&nk;f���p�0�7���,?�ei�;��k������%�ЮH>[�.G�(�_Rh�\I�l�H���,�Zp��/U�瞵?���}i.ӪR:�LJ�t��M*�b����]�Jn�������Է�x�O��PGzo 踧X*zc$ӮGY��՚���_F��!OS0�!	�h?9�%7����35��ƪ�J���!���X������實�%��˹c�