��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(��ἧX��P |�`=g��P��F�qW�4qoG��\�ewQ(^n&��G�u��ة,��(\� 6�S������X�'�i�غ��ƝǞJb05���� E���P7�ii�D���uҢ�P�+м몃u_�o��K�9!r}!�lk�E a^���.iO���f��F�I�����u�%ЛӃ1�=�$���V�n۬M���O��og����1�� �[q�-T%�_m���:���YN����7�d�RxD��|Qnb��P��pV���Z����b�[g<�0��?�R��f��Q?��w0Fq�V��V+�Qf��Ĳ�(��K��j��E�YuaE���^k
3���R���J�����f����90�.��l�j�9|)iV[ ����N=7%g��zź��s8�f��Oo��r7�NV��8��>�K���������|B_n��p����o,�(caϘ�uP!�Ѽ�*N�G樧D��E��7�*�Z�s��TloM��&ʋ^)���F<y����F�<_z���(J� �����=�[�J��[��<���@x	z���������f�45T���2H����7Kb6_ɉaZ
wq}%�f��<=@��+��?��ড�]��-�����2W�\�؟ytL�Z/m��HrN��籅�5���}���� MҪkt/�0�##�dwқ˰1��T@�1�)�@�P����φ���|�RKP�B�
1��p�%����"J��-��->~S�w΂Zb�T�z�_H��|��HncwN�\�6!*El�ݟ^rؽ%eZ$�}D�s��+�� ��Q�Y��&}e��i8qs��@r.��D �)�!���iʬ:��~و��:��
�s�N�k�M�2]�NſsA7�!����眚�_�	���1���k�]��)r��qу	 �"��%x�ٕ���H�"�#���d�KDN�)�\� o�Ş�?SO���hqb
���a0��3$U���Da�+��;�ߠ�d~g�u�0�"۲���9���O�6�������a�LB�(�X�����l2�����i�F`���<�/I:�K�Zzյ��K/ζ��y��
���qb����Ngō+uՉ�N��=��>&��^��Ko���Hl�ս��.; �G�_!�� ��º�e)<��}k��@�SL��SBw����k�E���l�Z��U�"n�+ї��M����@�ڲ��W���	�����^���ڇA�`"�C'ŉ1�� fZ����ߗFgW�M�T��(/�8{��q=�����)�#����.����Cm�d��G�2
Fn��X�h��,�!�tǂ|�=<��Z�m�D_�ύ�^k��i��8{N�"��D	t����b�=,'��:�����]�b�t�V@� ��Yl�q�VM�Q��i��t��%%d圛�M��>&����X��œ���,�|HC26\q�sLTf��'EV�b�MhiY��md��)j�B<'�Q��'�8ʃۤ9��l&����-P��\�����5l����Vi���R�4����\G�q�h[ah{�h���`��i���mr��1���_��6q�*����������L3 w�U:�G�?�Jj���m�!���C8_
9h�� 7��K��`� 0�.(����+%��l\L1m��Х0����r�(T���R48:��U>�{O.�Aq��4�8�ud�6@ȫ�Rԇ�q�<�3���F/���?��6�g]&n�d�������w���X�5P1��'���8.��b��̎7�J����5����8ȡ'��܄9�B�t]�o���a��s�L��-��c))�7�O��U4��&�P��;L+(���5|��46s�ѩ�)-��ڻY|�! �`��H����~J���'С��)i�\����N�"��֘�뷥U�'�ƅg`K��u�����lrPNٰ�ښ{�|l�f�����cz�:����E��l����A�/c��fC&u����b��vb�����������J,�&�����(���&��
|W�r���%��+�~�.Ꮃ��M��;��~���y�O����"z+ܫ�����`�k�m�PT��*~[U`� � b%��>�f��D�:���~���0[�����j�Z�GQi��g�$D�~o GA2�E�Ѿ���,;����Մ�i�$�r�t{��7b�(�u�x����TV����C��x�'o�X�c�KX!ΗE��X�w�/��E�0����T�1w�5��e���c�B������d4=ɩ�>6"�=!�Wwپ����ޱ�7�d����L'n�X����)�[�F+�c��/��3ٳ\baw��"]�;���D���2��16�ݤ_N����@�^*��ܞ�YqM6�M��%WT�OJ8�A����k�
D�&���6:<\.sF����cs��������(�_\���c��~�Wm�:K~[Y�kt���h��S
��-.���<l0Q�G���~i����<=�KU	ͩ:�(�ge����K٪RrX�&��������q�Q��a9��`�[/�
�d󄿃�a*�cx��!`�L�����!�$��b\�3���=S�p�m�P�� 
�o�6�a����O���).JI���┃�S]�8k0���T�
�T"��Q�ْ�jp�;��/��������ٖ2��ST�[\��Z�X�d�=1x����7�bhY��C�T��>�є<1=>naiW]v�+��F��2B���j�K`����W�h�Տ	p'�+�PE�P84'f"�u������,}�}5�`��]����8[��*ON�Q�G�+aB��Vt��j������簍B���/g�`�Yb�G\>un'J�e�,��[p|gyC�a�ݬ{�s��� �^��)��4'6�u%!mY:҃�ғU�X9�UI������0ן�>	�Zʢ�@O�"F&��і���[diQ�z����*+�A��}q-�?�/$"��N;*wHYLXj�H�e��Ӛ�*��99'��R�%�[�:�ɉ.�+��F���~g�}IG�ܵ�^��oU���N�o�o
�{�LDK �-8r�[ٻ�V��-��A�%,-@��F�q��6f��,�	I4@Ai�,��؇j�_2�͚���������G�;h�Z��գY��7Х"�*�j�i�4:�9l��U��Xe1՚`�����3�Nz����w���ً�0�@E�J��K�i	�������{���}��8��qK���G?O��Fh&�q�o��>�ۉ��_6�t�Y�C%��ʮV�8�5�	$�>T9��8�����c/kۿc$dҐ���g�y֙����W��������)�G'��O0-K*  ��>�K<V��N���1�Έ�_ĸ�,.���a����ϼ��)�4s��v��+��+d����R�5�a���K�we9i*&�;r���`�xL_��̰m�����6f��e5V�[��d��B���3���9�RAv�2&�B>��W�ʦm������c�B���F��u����d7P�=V^4q�܄^$픿�m1T_:l��X;�Rf;���]H�����I��M��Y~'/-�;�K�&��@K��_%I��ˣ`*�o�G�y;7z�rƇA�,��"T���Q�����.J�-.h�#�K$x�n̼�^*U�I��[K�ވ����:����U����l*
?���e>�T4Ca�3����?�Ҿ5�QE�"��ߺ>]A�	��g��>�v���8`������
0mrD�f���������7]�B��t����vlh����Hm_p/�k����=[�}��5o� ��x��-"�18y����c�µ%���i�2"Oހ7�Q&G��嘒۶���%��{���=U	���fo)c�#]3}�����y\�Q�fl���Pk����>�+�T��1v�IЏ�' c�� � (�Y�Dg�:�m���=��%!@�sH+E
+@�w���h�?j���㰺��@�2���ʞ�T;�q�9֣o+!ø�n��#�ҵ	���wN�A��roM�������
y���WIrkr)�.I97��J�����f���{#�SFD��L�p�S�˲1m��z�V�i�O����m�3	�mk�(�"n�CR��.?��%��aM��H�� E:kھ�u�0����a�7�ǁ&���E�6�b�7��2�Tp����xu�(E#�_�ov��c_L<�R�� �ˬ��Ξ���O�f$%U�V���h�䎗���k� �+�G�{52��ƫ<�D�c��eV&�D;O�73�]�*�@~���u!}l:A/�r���.5�С���r"��Y��7���Y]�i�'Ҭ=S</��F���|F��Eu�P儕v�qc|p�6GD�X��������g�z^���e�_@�,�Vs�HP8irɯ���n�?V3����Y�L��u���̟R��L$�KXj�֭9UF2��diD�JTl:"D���,�$IK�<`��!�*&I�IQՖh	+�XC�4j2)��g��u/�v���p���5��d|�X��+���=�|�?�5��s�p��Xg>�7��1�WW�j��
XQkr�a���r6���R����v���|*����reL-�j�`�����2'W��A�j?>z���ʋT��x騃X�݃, ����(q�d���-lm=81�x���{�ɨ&,Yٺ�oTu3����SH�ےGy�� :�%|q�
�P�P�������Np1y&5�� ވ(��bR���s9��~s9b�J^��\��7FȚ�ƹ��e
����{}�Na�:D��/�_�t�0��ng���J9�3�s(���9PI��C���F,'��������Y�D��,�.G ]��ս?�%���f8�я����'�{6�-\,���"�FGuAP�oc��(�l�/Fj>���HT��ܞv���$r2�4�P���  �<.����3�V�مd�"%5�R��l
�a��;����l4;��}���J���T/i�Da�5���zG�T����)oT���E�.�y�:r��Z�����f1y'nU��Vt|o�HF� V��"�5�F�V5�:=�2�[��S,lLy����T�	ƅ�Z�b_H{�u[��;Jx�����Z�� ���&Ǫwf�����L[)Ml���Ջ?v{Q��9��gv=�t��Q� |�>�Y����'�_f]Ś�NI�7�<Y�Y�~C���<*!��_�1Fw��HwL���K ������m�}����0R�d�3���%�6�^v��U=U��f9��m�=��C�3��x���p�b�����2.����a#�k�t�ž��\Z)�)�~��3����Hv3���?x��Ð�� ��z�|�0��b{�� ����sZ�y���w��>��$c��B�n:-��2S��rD �E��I�―�츶������%Cs�>R��%�u�=��V��<aFJ�,d፯�
���� �%����d:{ۤ�TȐm'�yPN��*S���˵��K>^�P�|�AӍ(�V��g۟�Sr��������p�<��#���w�����ȄUلm���g�h����f���p��K*
�E�9�&-�l����|D�M�a�>Y�
H��mb"�q�� ;E`�(�dyl�7�����x�4�Ӳ�rt����L%�dL�t�#�w��ϸ�����0�r||ԁ`�-n*BY�&�(�8�7#yĴP�2l��\�O.\%�t�����h�kK�]PsX1y��%/�:���.�=3�$[p�!?��1R�]�I>� Ǎ]�C��L	�{�Z���*Mu�![�z�bP.�`�NBӊ��*=Z�'����픅ل�;��z*��2��?"G[k���`S�%�|w&�H5��FUh����{SF�� V"ζn��⇪���3nN�)�!K��ԢЩ���M��O
ݭu�8z`�E9�% ����ţ*�6-Z��[Z~�2~�Tx�͘��$ryeu3B��㉹�|��d���7Xtz��j<=�Pۯ9_�n��/t"��y,�z�z�������hA��K�ђX��T����hxvx9�����)��Wrj���?z�S�'����7g�9��I�U0P��:0�%���FN�t�&�q���g���Ό� ���r�p���W�6�T����$�2�/3�\��W�뜞�ж��p�oF�Ҽ_�s�i�X(��������Ix�O�kG6�(=��m/`c��>+%,��z�0 6���=��m4���:f�Z�)Rhm�&r�F�WΣ��5Eǹ����:����߼QƐA[�r�q�Nb���y�rƨ{c��:�ݹ�cq_F�����^
I�EVR'&Cq�
�i��Ҍb��Vs���Lz���?_|�A����鸌���J�R`�\g,���m��S?�A7g�}�u�w)����p'r!t��>9܏��ܭuP~`�ß�Z���ЦKz�om�K�|�z��]��q�R.T6�
�$���M�rL�d�Ed�&|�2�|�̃��%�7��K�O�J���mG�V^�P����X��-+v�C�����=w��s�3?�~s������9	�$�of�ƪk�F]g�ȏ��)����)f�v�,x��l���CJ�Q��ݨ�p�D�1�m��վu��Xjb�p�t��h�l@hϥ)S:s��P&+v��ܹb�D-OyU�p�n���u�rWH"�{J�(��Z���	s����"�Y�cdj�X��4P3-1&���s���O�����~h��ye������狅��bG��c�����bxB�x:���U�U ��g�h]]�Lw��W9z���X�,�wjl�~4@K��m�<Z��[�!;�d��@T�O��""�!�#ESPy�	b/�\���E��E�*�O�D��Q��M2*,�b�6-��}����:���٪Jq8A,Cj��nG��v�.#�yjoyl����y�fyO�٠�b�������nR�p�Q'9CƗ����7U�q����%���Zp��j��(���Ƹ+�f�I�)>3�u�
��T���}����u�����h��"];�]ȟm�FF��(%W&�v����:��5ٹ%�NB!��q@��}�R-|K�k�p'�(��������_�����W�Kp�r�!�g`u�Y�$a׼�>����#���F
ChJ�vb��V��Kq�(�-u]�~}��fZ�s�����"�&��|嬁�*����%��q����lGR�4��ǟ���,��Q�~��/
х�W ���>���vu��H�-��N�
r��$��#�Io��eT��d�;��M�C<���������o�i�e��2PU�e�NWE��{z�ۻ�fVɥt�LG9��3��ݓ��t��ﳹ��XƲ��t�@�d�l
O������?��TT�@�,*�M ���X��B�x�)�p�@���8��b�M��Q����4�E�h3�BW\���m����Qb,FZ|�صܨ�����F1:]��>;�D����j��oe�z�vŎL���m�y�{�M��m��c9}qcz�v��ٿ�_a�(BD�O��M�fR�l�3&���=r�w�F��!���UX��)W@c��j���O���X����� <4��H#��9��� �g�_���PbB���4z�{��i�d��~��>�,d�������6���'��)�nX��"1���`M��Q� ��3�`F'K���N�H<p�bMCz�s�xgIq�a��!�P@&Zw�����O�s�K���W�s�B������$烺S3�,J2{̨�����]UR ��}G����s�A�D�������Х���bK'ć����z�TЛZ�#�F��)HR(��Zj�uUaҿ��h>L�}"D�b�A\KPj���EQTs���pg�BĪ���&��sFJ>+i��;[��ܖ'�� r�o����S��p��?d����ʵ~]�����V7ax���A��=P��?�7�,0�����U]���oY5IS��p�v�l�������u�mΪ���e�?�n4ᣙ6�l� �'�Jv\�Hf�����/@i�]��k��f�l8������{������-뼑�Ux� ;��$������I��h�����	���\b.���*�/z)I:�)*:��ܽ_4	=Ի8�֚��J8cXO9�����j�v30ێ�2%q>��x�!H���Q���Q->��.Mu_kP�T������*�^,1��v�`5!���0�K���sm���4L�Q'-F7$�29�ք���ޤ�a(��ߕ���C�'T����a��@�9�?���s!d/���|�(���H�ZI��"A�K��冖N^���;�����`��f��R%څl�����mG�/�A��ђv*�f(T�D@&����D�ۋ.�[��'z`�����=Zr�mH�	Q,�Y��'^��aL�9T�j_ ,����p�N���|7�����>��c	*����!�i��t��m����7�h�j7����L�����Zժ���y�n{�95F����{Ia�� �3J��`\=3�EAa�����k��S-�T�A��+C�1�zJЕ"4%�����Ņr�X�él{���7�R�b�]ԱIw�C_�!h3��Q lE���4���5��aM!�Ƌ��?e����P�鎺��l ��[ J�9_�b`F�kF<���9�bi��i���+ǒЎ�Q"�r:����D&}����r+0�)η��Г��ɦ�R��@�BM|"H=��y��V�=X9��g�H݃޿hf���c��$�#�F�{��nY���Ș�����l�r��,.��V����͸�^�}�˧�;�F����������A��t�QP�����Q�҃/xx�D�UveZ�6�vϖ���I.�	>�o���lNN�T��-��#�4��C63����/�{*v8�5	?1LC�k�K�ȧ���= VXO;��<wY,n��#���3	��\Zރw.�
��Kz��b�I� L=U�f��⡱<9��[��ȰVX�c2߼)r�eF�x$E!
čc$UC���݀�6`�@ ȟb��ۀ�n����Hq����2�v�y;�n`��VDE������H^��gڐ�p,��N0��F�>.�q�O��K��+�k�V�~<Qy�1��� ����@8G��=Rm�-2s�f�n���T�ܩ���g�ݛ�6����bymDH���{k����X�*���<ne�5ޒ[�v�]L^\����T��@L��!D}�j�V�Fݝ_� a���E��N��"�8w��נ*�ƭo��:�2���/�֤���d���N5T�UŴ}}^l1欄-�\ߠ��/�����m�_c۝�����*���q�RX���cŰ0R�G����R;���O��3�F���e4OB���!G��~��+4���qy��;�af�q�$� `Lb���g.T۽d*��k��i[���D�{��C������t ;b%/� ��z3��C��[8Id��Nd�|I��H�[�0bf��T �vvevq��#�_:�#G����U��a�~F2J�5�� ����K[����h�|��r���T�5Ⱦ��eg�?`�4����}/ҙnxhmO3h�=�j3FJ�rj*�v|��>�f�]U���T����iM�5�i�|q��O�]�m�;j�	Q�3���v<�{S�mZ�b+���]�{�������W�.����7��dY���M��Ή qh����ȆC�"��"����,�\ث���	�fW�h�X��� H��.�V��$�?	�⟨�:��n�k�˲ki5v�jl�"�58�݃�5�Ѷ�5%������D���0Cb%�Zf�
���AC�P�k�d���%�k{�\~^7���Zq
�ڢ}�L��:_o0����_P� �X�XQF���a��p;W��G�r��k2+���$&L�{�݃���w�|ـ��"9*�G`����t%X+)�T�7�>���-�W*�M�}q	[��;)i��k:�|��t>�T���)Q�\�
ϴ�bc���Ja�^�}�Y�a���l�-�S��<���r�G W�ٴhX��t5e'���Y��t;J=�TqN�<����jfc�Ε�V��9e�εhn�Ãrk+a�ԧB.���E�}��S�}3� 	رet�E�.�\3�;$�0���<�sc+��fr��Tm�Hk�n:+��k�ψ� 1+�����ׅ��$����b�������*}�y��L+�u6$@�N���Zl�1�m�6V��S�_�/��՛��M��ۓ�eFnm6hq;z�prd�dl��� ��+��"��c3x�rhU�2n"2�p�K��#)�M��Tv�p��)��~�K�w
�;�,wZ�e��O1)���y�+2eFR�SLX��I91�h��:���HÇ+���&�|m�w Z'nP�G/,�L6����l�tW��Ϊ�Ʒv������Zj=�bk�?cT� ������C���|j�g�����U���Rd�r7�󙷰��^�!�h7b[z���X��J�h���!�ӯ'��d�L5��{0q�졺,{�$M[u�	�F���ה��Tn��A�S���yܻ⣰�<��:����3%z�Z~V|��<4��1���!6�����	�����)��E2�=*���ٮ�� e�����[wI��E���IΤ���<<��!M�(���'��j��s�Y�2dY�i������jA�n	?���1�;��}{a��HN�r'�M��6��5�S+Jp���V��p�]��W��^���ZT9�b���L�7�������&��N�tx�$��=ү�gh��_(z?�N�dܔi���0�.��Bn�РG�}��V,,-Cn+�J�|���#�	�,*��|Z��������Hz
n�'%Iy�ͣ�o��t��W�����b-�/�t��~��ɩN����=�L?��8��a�|P���:Ba}��xi�X�J��'I�u�+�<Ѿ�Ǒ����f��ˁg�s���5HkH{~�K�=Q��F_|4)�<`�������v�t;ʌw4���rA4�a�%��	j1H˯{��C�9��������OO��\{�}4�O��6�`T����.y���j߳U�zadeٙ�y�UK աF�� J�
M0.�o5�B2�"�]���}�G��mI���X�it��� �ݓ����	J���v>�G0}��mn�X�d���t����i6��I�P���w_6�߬��^��5UՁq��%��/�]Cd�2_T�T¤n�j�9�j��(6{P(.���[p8$u��:�F�Z�|)�T`���(3'A�5Z�P\�Nt-�8�(��p�A���N>ó�Ue��j�{��8���~����#X��s4q�&xK��{�4`$"SJx���Z~>o�3�@���-Z�2=�[_ާ�5!�C�E�,YY�h��%��S�?�7�:��>0J���q�����g�oQ�:�ݗ��������U%��Ȁ�.ڻ�6���E����ס4v���|� U��>������+���6�E�;^��:.�h �'�f�|@��%[�:#��F�رTh��b��ǣ�w�7ge\��6�K�#󑣹�e�	�X*}�йP@��;��pc�AՉ`�o��9�EN�i���CcHH�`ho��T4A+_�*�������}wĝ��6c(q�Aw+��0P�F#��r̞��|Ey�g�"j���!���?44���#���IH��\���ݜ�g,_8�u�',�ɬM�$��iz��G6��/7��q���(Z�_��͞�`z���x�z���3�9wp�4� R��j;D:�E.��	V��<໏ػO��2��B|���hfFO�.�1Vؕ�;��=�հ����R��X;�ߛ���:�� �.v,�� c��ckd�[�ѹ���*�F%�ț�,��Ű��|+k�*�� vO�O�^O�,.����v��{f�j8�a�aW�������0�q+��t��n��Z8���7w�>������V�ц_Rm�0s�b�5N�U��DW�*+�_�_c�;4⬷�C1g1j�&�k�a��Uޢu��sJ��n�*	��脬Tr�'?����\��ZPD�grf��q�l��J�:X�����A�m.�P�Z֮=��^T��S(<`	�#����'��$�����R�+��ε/O����we�(b�cOgm��4DX!�|h�
7��t5��B5JnM�i�I�J���T�*cj�����b�UW:�O�uF	r�"�*��Z8��Iֈ�<�YB�^���V����DG�s����h�'��ï?�ю��