��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bdj#E�]����u�,޵;0�{Z�����xK�,���u����{��Z^UؠE�񑬉c_�pjT��l�+AL����瘺�`q��2z����������:�ی�[ɯ�l=z����w
"4�"�B�����(3�r���kf�i����Qv�Q���V�e�7c�A��(ܷ�R��eS���Ҟ�&�j�P������8�� E�L�@��B��{�B;���$kRd;���/�����a��� á@X���w0/�b4�l���j��p|0=I�7��n�'�H]+"��_e�ian9������DN��jmF(U��~���/�)b:�B���G�N»��.�ør�V<m��	j���9�se O&bU�O���(@��z>��xz4��k������h�$Ջ��sI�Q1�
 g�u�n�!W�	���h��t֒+Yǖ������JQ��ɝ�t��t@I#�ϳP���[1>(��H_�t��.�z���5[��),��Q�,/�%|���m��_� �c�����A���Qa�o��֏wo��K�- a����	��k�����c\�ň�yh� #�	ȗ�g�$��|Br��*�gj.�Ln1h�{��,��u>&$�a�ε���A��t�_-�A����_��O��їc!y`��ڰA?�ϡ���rJL�;ý8�ߛLf$���G���y*��#g���Ƞ�#�d����{���Q��+f�)��a�W���v>k�j�M,%19T�B�_�A�v��	|t'�׏���t9̘�M��Sxr�`�;\�(��s�u�Z��R��&�֧�Νȫ�)[@;���Q��������M�r}�e)Os�c��!�O�WJ�q�.S�r�?4����p+���i�<5㒤�Ta���6+~*o}��l�Y"�$ľ��bH�Ꞝ�畺ࢎ'�[y�\���Rt ЈnM�F�_.N�!.�X��?���Ul�(sҍ�����w�oy��q��^����7�N���D�v|�����X^^+�X��A"̨Z��?$W�s�ӄ��+w��Ts]L��ۀJ�"�)�`�ħ�o�ݷ�������e�H��U��G���Ȝ��lKf���*�1m�Fˀte�*L-?�3O����L��;�ޓ�����W�:��#��|���Y�/>���v�𛬧K������Z���!ۛ\�[R���u�+b�^�}|j��k��@���nge��\��ok��Kˑ��尣���R�?�n����8QT1�Î ��s8��'L7g�#����/�,$��3蔦�#>,P�{���c�1(�y���l�t���*^�o�2�wg�S�9G���;(6$�1�o?Z�'��������1v��=T��I����+Wo��qeu@����k��>�Л��^(��bnU�������{3��G����ƵE�t�,`�dԝ{�M<řyǚ�-����e��x�hycľ4<�bk�	������l�@a�%��#瑣1]��Ն\��a��}���D~��p/)rM	=��q���ӌbXP]V��g���2�?�4���^�����f�����*���E8N�Z�o'��Zo����nW������Q��ۄ�J+��663����囅�H�=�)�Re�[�M��F���
�t{�k�
z�Q A��N
���AE� #[��=�;]h��4�a��I�
����#�QT�P?[����.4���7M0ģ�b��`��c�M?��v�D�'K��XRu��ѣ�E �8%7 "2�x�s�y�G����gZ��5�$kXy����RƠD�U�6�%����f[�L���U<�?e_���'�Fr�Q��;~�̮5F��8���+FYN����b�ϱ����(~�!�J�=e�6�gr�jL����Su�+S;��`F�盌�ư��1�6|=!}ш?jn@�d�C���)�t���m:Y8x��x�E/�W	*t���;,i`�qlmf�1�Q�ue==@L�"�Q��?%~��a�3�;�u{0}�,/P�{W5`�9x���w�_���[㇖������|�h�^=2S��s퓻B+禁�uKi<	�0�����2 d������w��Q(��I=�!u�?�M��k��Ď�I�j&H��.�8Γox6Apʆ#��u}���a�[�aa�{EG������3��icn�6�ҟD�A��^�<��'�sn���3���!�{4gتp�����Y��m�fyM+}�ki��명lb~]����ˏD��:ѹ��;ݫ�+�Mg���k�t0B�*�.^тx�����a�n���.��I|\57�n1W�pb,gL��V�ގ"Z,��W{��<�S�ؽB}�[��hX��T݆�y��ц�%J\�B��,|��WiJ��b�C�[	?�s��%xE��f����/�l'��$��E��2iKVQX����v�E���G��N�W��Њ	�&ºW�X���Ka���NKQ06�v����O<fj���œ���[����T��m[gk�B��V�J��%���6ܩ�t%/�j3O�O�;���ܺ�ӥ��8Pm���-���-���ȿ�$Űd��"��$U~c+���!{\��2 �	�a ���=�J�V�;�{O��jgBo:��U�ড=�K���$�L����P="bM���xY��`L��GU	���l���E˕G�;|e�� ���iNc�F��0H�٨��-��w���#�=�ۘ�s�u�	!���=5]�o.ͤW���	=hX
nG�Jz��"����J�Yf.|�B�\Z2�mv�w �`�&���ӕ��i,�y\�1���7 ˬ��-�W|9W�ԃxYK�P���O���P��j�>�tėH��SF��&�ӻuΩ�;_�v��ƪX��0�Y��=g�u�2�����L�aX:o@mV{�d��%l
:ƿ�L��g$?�k��h$0 <(��Ά�B�Z�8"�;��B�e��E�7J�?L��}�஁�t؉�����Fn9���4�� ��5�
�!ClD�.�#y7 �Q�F��X��^�����}b�^&��0oͦz5b�>�c������*&V�ء��OjR�u֫�	�{��2|A���p���Q��H$�e�p��fV��#}]	�3G��{���^�щd8�10`7���8�E�K�z�'d���^7eN��P��o��<F<�	CN0�U�C��x���1<6��^�R+	�Q�э�� �r��c����T�+8*kH��r: �-����!����{����P�"��g��7�i�=������%�u.���wF��M(��t�����a��f>,v2:6����K%W���Q��T�{�U*�
 _�7�w�T����˶*��	��Z7W�<*�g��U�@j
h���Ӑnjל�o�b�R���R�{��~X7��ɳ>ː�S_rI3�A��l�AEp�u�@oz���l�y��n5MJ�{c����Q�$-��r_`�����X�~����;ޏ�%B�� ��N�lJ1��h�б����R��r�R8��a����>A]�If�ȩ�F�:��WI@ݙ"�k��׳��?k����}Vi����!*rZ��[C_�T����5�$��F,�7�$���h�I��?Q<����a!ۇӜ�<&Tj�h
U���Ĵ�W�b���^d@}-�"��/��ԅ��/t����]=���+w+�l��a��p�h��Tl�6#	��%�]�}ue�ɫ�e�X^��5��At@�X)PϤ���L�p��LЮ]�nȢ��K<�%p�ѵ�P�$ݝ+��$�������d��Σ{��}m��a�k��:�=U��l����NS��T�]ڳU9aX0Z[����N���t�+8 ��P.mr`}��1�cG"+}�P���W�gyF��:S��c9lmkk%*v�����i-u�lr� �`jF����G�м���J�Y��*Tn1�c�!��3f�s=֍	�)��j��O
�%�E��E���/.g�]�!#��&�I��*t�^���;�ω$>��Iঁ�$HE��{%Q/;_�t�@���sV��7f��{P'̯tŇ)-Y��e4G� �l5��\
{(I�.����dm�X��� �/!�s��y�x�Pg��i�!�<i��Y�]|g�	e�uV�d��~XG�
]R�O�x(B%�s�A�d��j�M��;��P�Z�I2��o%�S� �%�����[���̲;G���� �d��W��f��}���1i�B��L$`�&�H[ ���[E�t��d��>�����Z�3�z�b��� |S�5]���x���D�!������M9a�	,�E���sWi�u4���0�+_m�_�^s8�)�eN��/� B�Z@N�"q�ɧ�8���D�N^� ���+Y#
()�_�,֮n���nn/j�PYYKj��؜��-�;Hh��l����W*%�98}����阌r���@��U�n6bJ�َ$Tx�aNWEY�zIQn�f�tp�}o�[���/���"z�������T��U;�V�[��}��B�M��~ ��7�~�/�*h��>�H̤�U�- O�H��9�H�.�iK|+� ��@NW����#AM�,�������t�g]�M�B��]�p��. *�}f޸[�(�r���Y�"~����_@w���CN���p���/[hS'1:$�����TQ������R�Y[�=�ڃ���@����0M��TV#y�k{���c΁I���+O\�cE��������͂�'J�:��l���2>�8�����Q�+�,'8��P�*>�;^���W]��{9�+4�B_aG��o�>s�<@�9���0'��V�{��Yg���1��Gn�`[�^-�^K�)��ŋ��	ɽ	j��h�V971�
���We'�a3}�=?��x��,h,�ܿ��0��h�c���:�z��4_�P��s4+��R.��(0�-ب+T���c��i���|�:���ĭ[aA�"X2*	Y�'�����\�����z�12m�a$]tv�Y)��P<��ݝ���8��`��X�t��^�<LH����g:�Y#"Sc;N?'������g����(N��L) ���ޭR-�z�B����tŴ�A���+c�aW	����Y�S_0A�b%r���>s�Fkp�ع��@�/��2�ƿ^p���)xA��',��zi-��U��\~PaDoa�n�4ջ�jR�ZMP���e�/��H��tG��a��,��K;���_�U�J<F�I���T��$A�W8gMe�� h>>�1��n�tڐ ~5���lm:�%��e�+��렵��Sbߘ���Pyv��9�������W<9f��K������}�x�K"k���t����&e���%�S�zm�a�ջE�W`�'�����u��@]S3�ϧ�/u4r��5d�^M�f-O%�dz�u�6)��!%(J��<��3[�`o�M�E]������l��h"䆳�ךd0�l��^{Y��9�� �<��]r��q��b�0H�"�����LZ�+��J4.yhPz{Mz�� ,����Ѻ�"�:��WI1�p����4z��[DX�5@���ˍY���� %�yMożw�S�w��bu)�x��T�p�s{�дN���k��)�S&r�&�Z8�G��$^��Y�>�d*C�?�K���w�ٹ��2���[�=Y������V��t;�覍{hYx�w�\W��)u�W��R�z>��Nw�^�'<�k'��� ���f]ewY�J;ǧ�m�&��Q{ ����Ϋq����}���܄��	঳Ab�\�q�p���"�L	��4f���UUtv`'�Y����mO�'����@�AV8��g%�>0��u65����n�}1vu� ������.l��Ҩ����҅�Z�:����ĉ�}�)�V
���=��EB):+K8����]�y�=U%��Bu����Q��I�#z�S�)��¤�-�N�E.�{ň��j��j��?�v��$��Z��&l%R���p�[j�!%B�7��e��RqtL)ͳ�ƙ}d�f��J#�̏�P��rIpE���c�F����	b��{��( #'|��`�C?�b괼
�����)p;Z���bY�<�Ԙ}w���-ݤ�ZЉ��`1Yxrx`W7G��A�8h� ú�5?�B�S��Su��e�=qn�sN��������n+��(ٺ�J`3�QKivU�����[��~�C��6�~*/� CQ�kN�&E;t�4��[�<#� �=���;%�Z��|� �����q�G�F�A��̛��ٳ��^۷?˽z[�ї}=D�?��ܰ$0�)nL��Dmp
� � �.�j�L|dX�ȷ�D��!� �"� DW�$�A�3/�kc��-����c�C�}�v�,�(]}�!���1���>�w/dcep��$��]�,���Twۨ���)�J�A�s1} ���l���^�FWgݷڿ �H��K3�aA�2�8+��75���Q��v�5�@k�)���=�"�$���͒I!��L��FС�TQ�h2�4�}��Ǆ Wa�S�s������Ep힢�����^}�a-��EGIr�n�5X"�51�����[���Am,�?��n7��pKK����(ā<<{X"��g��w�?o?�o>�p�˄���T��RU�?����0W�R���B�G��uoK��ȫΖT�9_�oN�v�	[DԀ�]Wy�RV�^���_�������X���ku������k�!EV��Y�8�D}��mp��t�3j��CM�nC���E$,���e����y!u�{t�|NB+�m6�4��"}oS��5Ll��\#�'�#rG������
q)�L���F���!�{��C���J��K;��*�`\�[�y~��M���$���-!p	����"�c��v��1;��)�lhQc��VT���1r{��N�����^���y&F��h,2����Z'��{@�1�[K"V��A8N��D���S�ߥxqrI��>�?0"��zf�oXŭ}��_���"eZC]������ԭ\S��I���SDh2.b?�ܾ�!�n�����w��7 ��=����
mr�ŲՈ�s�Dd*��36��� �zb�����j�j�Q�ϣ]�I'0M�7a8�{�{^y����V��?t�쨂��A9��H�h��:���-���\��bU56x�9̹�:�~m������.dn��K�oȷ�ff$9�v���B �8^�4N��z�VN��p��ع�5d%>�3S��l�}z������u�$:��2��+d��`	��:�a���\�U3��IMp�L�Ewn_�(Z�ѵ��3���{���)�Ĉ�#+��쑭c�D�U����k<�y�d��2Z_FSu��ư[|������{���GD��XcI�f(���?��������S������0�Az �����%(x���h~g�tV�����Z�Q;Ac�q�7�8�:���G-߆ao�(J���1++"<��c仕��xu���MX�����=����M�?m?�b�oQ�%�\Z�+-ޭ\cK�E"�6�C���~{���IM'	���nF���%�ީ���<*�x����]Ӈ���}�3eQJv`�ު�E	_�ŗh�p��)����o�FɄ��fj��/�窙�&������8���S/ُ.��-θ\��B�<�Gw�4���G�4��� L"-��v�d��cJb���kn���
V��*N p�K�T&�S�6�_@���YM�t�Y���	��Q���zެt�c��x+o�9گ��k�(`;�[�(��>����o�o����BF��+v��x���l֮��#a�����˕�dm\	�v�"(���k�ll�#��ݟ$�ȧ}��'$-��!�Y_�+�a�-�K��e��Б�bɞ���zX�x�)|L����t�@��~���|+:-�k�6xw.Y�ɒ(�Y����6x�w�3�N1��7�G�xϐ�� ��jcòK��Jq����~bI���0 £�s������X0yޢI�!�e����4�F������J����0��x:Ji�G���/7JϏ�Y�l,2�'R��M/ҝ�����������2�0*|��z�HV��U�L��?�kg,�ݒ?}S�4f�.���@b���\��PQB�L��',�t�X��b���7G�"��Vrٞk�h�A7� �sJ!	(�P�q�%bl���� .�h��ݡ�j��qva`���BF:���]/��U����FWD�:&���+IY2�Ni.���A�̕$s�gǵ����}�
�m�F[[V�� x7taH{ x{��Y{�᳼�wTR�����J�?�t�)���b��o3�;����	�_w�Y���)z>M��X�"x�_)�7lI��Bf�s�1ʬ��!q��>Ʒ���\��Jfj%>p"{Q�ҟ�vY
������g�1}��zsq����B��7���O��R�f�}�Q ���Jd�6���M핣8#��UO�[|Mw�ֈ,�W#n��ǌ�K�Kfዞ�}D�B�a#��|p�U�cE��U�_��B������SM/R�vE�� �y��V�KG����m��[{����zs_5��4�q�qO"z��/�A�L����)�s�e�"j�q����V��R�L��[�
/O�d��Ϫ�|!���� m���[~-~�=ן�'
�ߧ�{(R�ى�V�o$3�5��n�����.�,�ҏQ�p$��_77з?A�ݫ7�n��.'!"0�0���nd^����7W�C��/.�P����lN�Ngb�y�	��{b+�N�Bj�t��(�x�s�� -t�1vJd�l���w��o�C��R.�S�Y��w;�Ŧ�FSTXzӷ�r�ZB+叅}[�SeR��f�C��nċ|=���	jU&
�?�!�8/��s��9��)m����3�ᳩ������a��D��i�GD��{�"`�b�V�YO��w)��ʋA�g�rjv�_���n0Y͟~渂D�	�kv�Zm�Qc�ޫ���m\�wgt.�:Gb�
�xow�R�5 �H_f`ק��иc�*Y�}�ft�G���1�у����:�C�N)�Y�6v�3�}���G�k)!�1�C��>k;�
жC�#ƀ*���,�a������X���ftr�_6�rU��pi@�A�4h�?j�q���g�W&IM�`Le�����=��r�Asj��]돛l��3=�ǅ���(��[����Ľ�
	ŶN�?�0�1]s���"d;�gn�zJBy��D��#�:��[���qb�IbҠ��В:�!��o]�EXT�)��$�(��3 +n h%�ǑL�X��=] 6��ޚ�!���W�=�����i3�e�r<��!|�;��گ�WU]������?^l�k��~q>���h����,��x�>ص�-'�D<c�^�'`ZJ9Q�{�j�Q�j>�ʫ�%�x�J�{�D	�Qo|d�(
�*�\CN��7ޮ��r���'��>W�ƴ �7�:�-�G�5��f|b���B+n�h��kJ0�SjH0���lzA�.��np<��Dk�7[}���SV��P�ˮ�=��0�������Vl�$W)ޕ͑��S�pO�P>�6�Ľ�MIs +�XW}Z7�+h6�[��_��9��wGv6�ǈ>��s �6v:O�T`������Bs5�
�.1� @��O���qT.�AX�`J�;�/���YQ���4~5�K<���4�T�^%�����ԿYZ�0�cO:��r㎓�H����a^�_U5������y����y�0��;��+�|%u/�]�2�j�����eUh͊f'!|�� Q�#��喗���U�B���a���.q���].�D/K�ۥ`�Xš�ܴ�s��9#��"�E��Nwհ;#�\;��\�Ua��c����t*��X
��C'Rt�ŭ�Mؒ�m���B^�a� �i^ϐ�<���*,���>����s��
�S9n.d�J���5��D�U5������5�~v�Wj{~�;Ѽ�.f���#w�o�����t~�?�-�0��6e�����&a��x���$���%T�������CQ�������N�Z��Ku���8��K�`�6nLY'ߋv�ojM�@�8��̹�����s<�
��_��xa;04v��}�v�S�HS�ZB�@�E�d��Z��j�"�1�'<��$�1��ғ��� ��j�5��)��zi�H����RO�2y4�&9E�,l�(L*�A��;Z��b�D����D�;�71XU5�<ˁ��gl��ER	7����~�YmV�d�����,W,=��z���:k�*��D~4��w��½`QᎷ��k���H�v��c�z,�,';�@��+FMFhr�LCs4���p�H0����/3y�WYtM^?���{���d����5v�S⯟c�.�bΛn&�W��qk�@<^�3ek�K\��c"a���c�t�=g[�#;M�'���Kynb��� �����cIuDެu/�|�,V&���8�sT* ����݄T��E�C1���Ґ"�H����gT2��౾L�Nj�
�>+��OJ���~�n5���K�R���!hD��3b�g�"n��m���U(����g�uᆀ��懒I��\	9t�`< ��0��rщB@�͢ƽ��!S���ֺE]�J�G���,�l� �N18��Ĳ�?����$?�OyT{1Gt��h5���9�_[��R��O}��H��9!K��
Ҷ��y�"�bC)[��0�H-���MR��@\�t��_�����7�-�����u$�3��`�����Ĺ	�ু�(s���K{��Jv�{�	��nO4�b����"����h��Fp�$��4��j��i���4��NQ����^���]W��D�C��p �!JJ}���J�İ/�!�f�>�Bkx<)�a�Ƨ)����԰����:Y}y�� ��Q���sdm�����s@ۃ<�����	���9���Ӻ%����|@�-��~��A�:�Y���y�7�E1�	�S3G[s�d䢔%K��??�ih��9���ǘ�#�aFnc�*�u��s�MZ����Ȩ��^����I��F&Z������'�+����؄5�{:!Zt:��TP�]�N:~�?��g���6$��c�h,\9�K��Ck��-��yT��1�^1Dwmdxų+++t����w�s��`q�y�.��pYWM` X�/�1k����Ө*��Ɗz'iM�.Y���%Q�S��{��ұ�;�LT�op�SX7�s$���N7M���	/I.E$��/X (+��*�D��o��yX��$�/N���4���b:�o:�Zz�˔>UTP/�6_^e��Fxӯ�&����� I����&�a���
&��i��⦶!}�M��T�'�d�􌽏�l$)��"4B�r�8��O$ q�,����� 	^J����y���t&�;��i�P������?[
/'n]B��T���c��ߞ0����ȵ���a���8J� 6w�k4~�5�$/JnܦݖG��[��e��"vgC��*'qCYޮ#)黹���5����	�7�b��'
@�%��u�ڎ�	�� W=!�9ؿ�ֵ8z��k����\1cPtꒅ!�\��"�#�g=�]��ri�����:��z3��kܣZ%}N[�\\���W�*֭�^���+��x�H�Z��������?�1�Uc{��s�*���r�rH�v�_ҩ=��;���*�D���S����K�6N+0LE8#�n���֢C��3�cgM�U�2M��Lx��]yp�|�76����<�ǟ$�/>��q�ۆƑ��;R=3�_�қ����>�	4���٪���l�C���8���}�/���X�x���㾶�A�$��.�槬zt��x״���P��K���^�ˇ�K�'��ȩir:vV�O"��v����y�|GY�<��&� ���m�ܪ>-3���͝=� �+U�t۳}o�9Ym�#������\� ��ѽ3�5��L9�4GEؾ�ʬZ#�Y�P!v�#��G-�+T�SY���\�����ܱ�7��aE�ZEO���ԟ�U��k��y�-�@_x!����ʔ{D ZH����v�����	Ps�s�Ŝ�A*��Vx�M���L
�Z�U�M'��V�k�uE���S�xL.ƕ�ɒWŧ!��'rlܬ�,�J���W���tR�%��C�M����NU�^�\k��q�ƹ��D��,94岽���p���;�%�����N�&Ǻ����4I_��v��<�����W��s�Q7�����$�\}�w�DZ�P��VNeJǯ67��&��S�Z�����MO/��n��~�ZkeR�����&V����r�B�Py^�_ᛰ�(�A��5B�0MF`�?2@`���R����KB�v"_:2�Y�ZM��ƿ|�%�o�:}~�����I����>v�[�zb{g��c���w��:)-B��NaTx�_s�k��ݦ��L����s��jO�/������D��*ӫc���g{,�xVO�NRM����h�c�YnH𝢨&�}I@EHϙ����ֆ�M�����jߜ�2����1��_�ho2�=�
2ji��*�ʥ��z]�9�}�R�2a�)Oг��1�1��c�L�1��z4��( ��$���&Ѐ��>�zb_�|N�m(���0�ҝ�O�^�cP~̩�E<5� ��ۄOU�d�
���\�!D���t6��l����o�L Ijjbskd���)�MY��;<{՝@fy�k�j�o`���S@���p����2ЀE�
�$%�2͞>>T��ĳ���-@W>��kf�D�ڠPHk!��3� (s�Ъ��X*���,��@<8++��	���?���9����pq2����k2\0~���r�e3���ɝ����V&U�A�
��|��Dwp>�7�>���fr�=���i½ݪ�Dk���E8%$#�����>�u͵5��wU?K�ă9v��b2/e���^_�zzi��μ%�Q��VY�2Gv#Hw�hJH,Ǫ ���`�����ytF���k��W�B����\�z��-X�V�u��ɢS�o��8
%����8�V9�EK��gE=ӫ�O�>�YAy�7~S�`�au0�
`�B��*Jp=���:���O4
��M�Bv�L-�k}��`0L�'��	&��2ե�	��l���Y��6�׾7�p~5i��k�R)U�"��e����7V}��
�8;X���	�mdo�হ�`��T�
m&Ã���k����l������܃���!��&1ج�~ K�V���XN����S©,�0��.�l�	>ٜ�JlT˄��^9�O	Z�MQ7��e"�k�Z�
��<�%p����y����4s�D7����-��mNi�9E[k���1ڸ%�0� ��H�>�ϊ�y�D��X�ﺚ-h�juD�Wm��ؼ/���Z�}ۤ#�1�g�B��OgM�����ݎŵ4��!W��g�Fi��?��:�j�����ۿG�i�7���G����D_$w�Y��
���P�Ҷ���[��F�	V)x`��ċ������s�0����}�7�3i�
��M�b��R:(�O�b��@"��/$���/�I8t-`��|C������m���b�Y�eG����S_�Np��y0>�_��w��x�����y���;֢}'`=9��;ǹ�ڞ��!�3��j�!1~h��Ќe�����Ț��/(�mu�⹫�۟����Z�#��Tnx�U�^/+1��̎�| y�)D���Y6B��%0�%�[w\��mB��8�A�Lt���T�@]H]b3s#�5]��r0{E�,���O��� �����O��� ����}��:�Fhi1~ڸ�
�<�{�ؚ /y��f��{4l�q�EJj�xtF�T�a��B�p��Kމ9N8�T&�9�2%;L��ᬃ��m2$D��5S�l��l̡����t����A7B<��HYm�G�K�֛��q�l��S\��"��yH̉�'��Ʈ�Ks�Ch�9����<���K���A��]�V=,3R��Vg�Š^��#�(�`oֽ������~|��"�+T�bt����58-�H�>��޻Cg��e�Ȍd�׺[Zף���0O�J�5��'AGjn��~v(��i�K��i���eq�'��QǟF7�J��!9olO p�"�	׊�}�i@���稒؂9�, ���<�#��c�xj��P-W�k�Ě}��Ta7/�ߟkN�ݨq��]<sC�Y�|WX�`z��?I\֖͡���q��wJ���{��*1�j"(-j-�	��#��k�����m4�ЇCY�v�
�L�W�楠˘t�J�� ����B��pB�8ѪifO��rk7����=v��A�x1�����n�@aN!���(-�I. �;�i&��W-�2�x����r2�^��4�Y� E�~ecy;~��ϑ���E�~��$��jA���$��y_����lm}禎�D�&6Rg\�@�������Wr�w��VC�a���i�� w��r8���(�0[���/���Ze� ��b�*^h��DH�5g���[���G_A�]�lbہ �TH9���a _{�n1y#KV�
����W���k�ƴ� `LG�9��y/J�+�Jt#f��syq�9EBQP�+V��C�D���/�z�۫Y�_L�����!�܈�B��&������(A8��+��`L�\§E\9�8���ޓ�h��UX��7���Y�(��&��Kـ���ZJ���MD��6r�`��mG���1� ��$�ϝ7ԧ�ᚘxE��ڢ��mY����v	�I~0{褪��L(zA���;��Z���b�L�ekL����&ǉd��i���s�&Gp�.�{u��F�= R3�������XT��Yb��$�ǉm��`�^^����H�n���A��˽�p��n���h̐1l|��.C�y��+ �
���W|��Br���o��T�+*b��訷$bu>��2;�6׌v�h�G�� �G�!�G�d0��r�K*

ޒ:��N����i����b�8�=�
�Q��a0�p�Bd�c�e:����w۸�.�@ �;��G�tmD����"��6l0ǹ�?�jr5jU��;e4��[�ܸC���h�-�,��Ƣ�}7��H/a�	�N�-��9���������)\����rܪa��Î%
$}�dl���'X9N�$�����d��3XL3wUpJ���u}��v�ȅɼBim - p´4*qY����&���.�fn����f��}�?���*u`i	�4�P�7�S�5#XHsa%�CH��	��`����*I;yq���fˎ����4���,����j���8���\S���c&WZ/�	J `6�㴀�E�{�ǜlp��BN$�6Q�	E���>#�}��U�>B��m��[~�y�+�5���|�z��.�U����_�׮>��%�b�_�vv�oe}8�%h���a��},}��C�ՓB��5LT·r�`:?��C%&�?�|ڡ�ͫ����Y�w2�	;f�%���
�� �õF���mP�qB��\��	u�i�鷏+����=�u��9��	٪�?�
evz����_��(����,f#�1fr���*_W�Ul�	�:3�qz��F�=!ؗ8,ź��D���1:��ܥ�x���6�I7��鮺�v���}�F8��$���)�a"���e`HhI<P2q��G��E=��}j��u��ď�rn�k7�������f�����+9�u:\����l�E�H���@��K�İ�6v3�a�`Z@�>��O�Z�?��ӕnw+Z=B�M_���5��`��c�=)�U#E�l�c{����4�NF_��S�褃�|,�?Z���z�,2�3���Ǡ+jo���1��Ѐ����Jb��{��-��,-җ��0��dg\4��,����3?ho�Ѿ��\.[ԫ�O������#.��$S ���#�4^�#p����l��t>r�����@M��}��3�M�i���i'ij����IQ� �ֽW�1旅F�f1���?g�% ���Ss:�@z�Nk�CގoY���"���"�л�V��u���}�cd0.�,Ma��:�e�0�������֦��͠2�<v(�V��F#�'nsV��HQ�yILO�缮����������Q�)�Q�ĸ��KF�i�����-����F�=ENH����T��e �LGm�&=���^p};d����%���l_-n¯o�Ȱ�����3!���`=��%�"��#
�!v��pcN�g��G�i� !'D0�3�f(6���|4?C7����2�Z�pO��-ᦕ[�Y3��\,�)n��jh�˪����(�`O)��ͧ�H�M����ی�R(畭���������dE;�3߈ce;(�z{���.�2�^��C5�������8�x&EeF�D=�-?[!|�ԿS6��ǭ����.ڹK|���ysU��
�X�O92U�4A,`���`1����Ռ��+pkn���Ht-�%I֖ ��Wjk;��XA� g1=Vg`nG:�\�
q�Cu���Le�OL�f���,�"������{�a� ��|4�}~��ށ��Eؙy9�.A�լ1%�S>E>ne>�5���4�#���BAz1����z�$�i��Gb,[��'������wU����[<zV�"Q���"/\;�[�xtk��f��V,B�
vm�}�Q,�4�9$29Ѿ��#�߀��"p#�}��Sty�6n5q9��Ih�Q�_+*��γ`|*�ʹ� �lނ��ԓ���Cm�V���mt���92��Z�Y�P�5>�i�\;���bM��D���!��0nkڏZ`dM�pV���`�o�!�9�Bț�������13�י��۳�<��!��:ҽy���,�l)� �eo�h�2 I��s�̸�RꙂ� " {힫j�_��g
G�gj"@K\	����y�U/�EJ�X�yWyY��L��&�*���[�	��G�����\�-�����WZ3y��`��
pi4�l�dI`�Uԧ���%�+���>I���9�#��ΐ�~:�]H0�2�>��&qӮ���d?(�u��G� �-����Źn�P��%�&��H쇍��
���ܾʅs�@�w�֥a�iGKЕ���>��d�[*3z ���=O���W~
�]엄�p��Ζ 6����;yI0S�_Ö��m`Z�2<ڒ;����赉��@/t���0���o�ض��v��]��$j)��P�����>���1�ݡ8&�4���e#�o���{W��o�Z��W�p��4�=�� �9�Eb�����܏�S	`x`����>�"���ڿ�d��I�*Lͪ|g�|Bq�[̓��ݮ�X$S]-�bW���=�
t-fV@8�����&��C�P�'�*�0��IW%¡���y@Z0�&Wy���G#x��֎��"�󼠌{U��=BQ�y��Xy�[��m�t�h!jm(�hS ����G�|�t��K�Xw��Q��_+?�w��2���R����vI��ls�h��Y�S�!�6Ɍ[�-�I���/ֳ�8}�tP�4�3��U��K���{	�wd{���,v!$4M�ui��?n}5S��m�9N���κ6M���e����=�'��os����W:�4����{U[�%�[J|���co�s�LT� ����#�v��cИ'^zT̿��+Ok�ej�Ó��yU����ʴ�Ә���J��H�{٧�h��)�/K��|��ˣ�5��0���}' K~���w�T��ٸ3����_M�ѫG�H�l�w���Leg��H��k>&Cw�0<k�5[�ϴU��#H�@�T{���a��g2�MЃ�f	�Ff+B���gCBn7�\;���d;�b�(�>�G-�<�B�:��x5�yR�~�YfM��S��$���4ҿ�5�삗_#��V���f�8/i�������F�G}V�J�������o�9�\Ǿ��Y������i5��3�L�Q��S_�++�Q蜁�tݙ �%��9�>�e���X.�6eW���n>�I�.	�1%J g�T��9Dx��|�}��$�G���ԟ�6����!"����*��J� k�-�UaF0y<-ׇ�Qcgd�1EZ����쀷�����B��v��>;�V�kـ�d���V=a�����v�a�OQ �:��R���Ľ!�ʥ�Y���p�g��~3J�[z�my�j�a��-���;�o�Mp��2�|�
���嚯�B�|]9�-�h�ޱnĞ-�F��OY�"r<��6�R�YnUYD�_�J�#G���	��dOA#�7���F��Ҷ��� Oa%����<���|cT��mQ	K��<O ����]�Mr�ԡ��^�R���9	J�m�L�v���T�$ΧP�:X���G�ߤdk���ۮ1�F���̟��|��Ew�[�]ǯ]�q���.�Q����,��������|^��RT>��h���#�^w���ش��Ϙ]���)�������l6v�^5*�;�<U\+g�F~���Z���Q)��ު��!��]"S�X{��j\ң￹��T\�rk)�讶%��(���L ,���Y#H��c�-�%"'�Xe@1	�J� %Ѧ��5�E����s�(��+�cqa��;����tŰ��wϡ�ԣ�,F}���6���ű}k��]�1���x���LF�a���7q|��]�[�T����Y���x�ݦڊ5{̏}a�}+��*��M�6	��S�"v7c�;�Q\u��J^�[�@����=����u�,dG[�-d+]h�[�����4��r4�J�{?��7���b�MRL�#oâ�M�������LN��fH�ʫ���T)#n4|������<\k-i�#���5���ad��~Q;�`���ov�3'�ͽ�#Z�i@��t9�׎V�8�%�(Uq��⥵r����\�6�`�Bv��؛
Ou�1G���.3p$O����7�?QՋ���џnd2%a*��©���m�r�G̙h�oGõP8z�F6w�u$�n( �k;�g�D/�	]Gc1_����Gs�h���2 ���2C�]�͝�@� ��Z�F��o�@t���9��Kv��K,q�!:���-�.��Q�p��R7��\-)"���,j��pW��N��r����-P��V���K�@o�#7�g�k�'ɶw�[zt�����_^D $23�贒eG���v3-��7��_�
r�a�e8�c	�m��B܊��]��RTէ�/�ׂkQI�np�	��yU��J�5�?�BAf "4�܏�AP��K8
+?���d������n�X�<�Rw�j}�;v��>H�8���X�M��>e�`��ȵc�N�]J�z�/ֺɻ�T�ۃ�b�s_���&&*�p?:��<z�.F���L��t�uϒ��:��M��Z��С�Z�rR'08��~�J�/�y2��y�����+$��bh�4.6���L����~���]&��e�Gæ+���2�k�,�B����/�����7	Uӱ�3�P����Nzw��`��y���n�0�Z߿��w��CO�	�􇧛	 �s�3�4��вГ"���J؀����&�ꃶE5��s�̥�9�' �����l�ؒ������Mb�J��곙��h�x�M1b�곍
�#\�?�3� ��v!S�$�&2�A��: {�L����x�Oj�g�W���v`x������*!ב,���M����
�i�ڔ����
� *�pخ*��m��t� @���qO|�u14�pxej~���!�c����C)b�zz2��� 8�
�i'/���ݢ!����M���Z�i!Y',��Kp�������	p��A�nX��Y���r�L��O���|�N�EH�5J��f�՛�û�¸YFR��e�ȃ��Ii6K�?�*�`:&,�Zz�K�w������%+Ed2TÌ�-�uZ�����[q��Ysw�	��]�����h���S����.gi&S�qv�F`�r^��|[pb���C|�|w%�El�դ�e�ү����{@}�
��Aָ��u������S�R�j�Ώ��_�4k���T�(}v��1#:�эQ�����p��}����=�rfM>��p�
����I��t}{�L0�e���>D��н2�_�PBm�}�=�B=�> �B���j��2r&~�'�Np�P'2��~G9�|])�ю6b����Q)QE��IH_�L�|�{�І��h�yHz��("7@0d��IFh��/
��c1(��b6����P� {u���E�8�=y���z�Y��fTclٵiveHo�����dS���OۑA�M;	�m�N�zNȮ���
������~
^'0��--�y��O�v�i�Au'�tm0jA�vU?�F��.��;��l17Y��\2%'�f��訓d���>^\������1��]�F���%��0mS���\��c�0���I�v��+�;�KSD��K�=��`��*���\�3���?&���\��{7�4�l:N�Dۑ�H�/�b��آ;Ix	\�D��q��R��$�6�Ꜥ�>����s�0%��R0SP��[ ��:��Xߺi-ԍ-���&���.=��2&@�cOQ�%��h��A�3���=�A�S����1�T���򑜺²*��赾I$jG�;���hD��Z��#�cy|p�Ű�i4��p/R���!���|��@�.����<�����MO��V�S|1�>Y�r������M��>�ʞf;}W�~��)8��(��d�to��[�u������Te�uD\o>DAa�Ȣ�|
k߮�8'�\�z�d�����!	G��i��'�ռ%9�
JEO���{�M�FW��Ӯ2A�%�ZR\�_5*q�>q\y��w����2y�A��Y��P����|�X}h2��T�䞀W�%�ŉ�1:�J$N�:ͷ�iWg��{t�s�u��|4�"/���@V�]%�i+����xsʗ�s�$w�F�����R(9�6R�$�7�@͉�֦L�� ���x7Juۊ����� �i�o˔��:Oq�2Y���\!�,S�q�,s�|��h=><����@a�
���J�Y�nIpL�Q�b�������8o
TzlUoo$^s!mǔ)��ݜ�$5c��n(@��Ucq/-ѱJP�6�us��TC�Kj��bVKs�a��ID��8X�06�`�?��sO��y����0��J��YVr�e���6�*h��ԐqY����i V2����%,.O�ޭ >�(�4� w��x��V[�t�[�/9/�@�J-y̱�e��@3F�����#]C.8���8�_��!�o���%p`a#j$oQo�p,��Q]���n�L� �Kď�6���B����xE'Z!{"6Lq��8^AQ�̙��A�DO����5�c6VM�>&�L/�򼎛B����~>���͊~j���z�u�ce����w�r4.<�[4o��k劺�2�\�O.�L�t�\�p�f��ި��f���k�I}�	E��Ќ.�d�R�2�-:�5�����'����,�\���>��c?�oE�=	�3�
�ؽt�Ց�*��^��/Sz��b(�c��*� 3������h��E�Yj>���d<��VU}���/gW�v����7�?X�RŜ$��wT�<��5l�Q8<����	ta��Ճ�K������E�$[nm��݌^JXf�/=<�vtb)�?6[���ቒV$��x�2�8��0���0~OX��J���k�w�����{���C��/l�Y2�A�ׄ��-2a���4JZ��� ¡2%ޞ���*D�pꅭp���S9� '�{?ķS��|V 4-�����/�KO�ܻT"lF��/l�����Ǹcdd���X�өse��$��-q�+#�+�Ԣ�����pgW	����$�:��R�޷B��U���_���z��W��e�]@�+��#��� �Z�Ď�g'`��]S�_��T7�w�5V4���m�px�c�hK���D�^k�b�Ta�jT?E2A���;�L��YS;@Ǟ'BG\�+��cQ�� ��w�EJN��VZQ��hK�5��T_/�����K�b�S��|��,_[	hw ��ծ��7yyP����2�_�K��zèn[B�_���w��˳�����>�f4���q�v$i�sw���A|��f�[����6 /���
4ȩ�M��`{#�HQ�q�Ȧ.OIi��#@4]�	�RFu�T`�xȂԳ��˨���{�_&h��T/��y�n$xM��؏� �Ub�2�7��-��Si��lk^�])%���T��e�F� �<7,k�ˆy��G��C(�P�����z���~L�:R�
P�i�z��E�}��{�Z��F
�$�������� F�Sj�˰O�tn���*���Hx�y�	*.�����J������ r��6��3��;����}����;������8Vv�/ X�عܧ�er*���I�i@%�b&K�8D�=�V�~H�SK�	ǌƿFPO�"(O?Kd�� T6�b)����?!�%���<N��mDO�e%�U�k��K���S6;>`���ѴsJ��_��xm��ໆEw9������F�� \��j�A<\E����S�S������3��c�U�"�Q��6�0�ISi�W����6{8���ݎ�f0Ȩ�!h�*)y��&?<��W��%;��Ϡ���J0�}�0e����T��wX�	�!,���h�`?ū��:(sv��P�o��[]B�*˵e��!�}���W�8ϩG$��k����G4T��[�N���WqmW��*�����ĝ�'2yBp(t����_,#ŦZs���('I�)�_�4׸��2|朒���#_��?k\�����F������:R��(��g���k������/��P�����\h��N��S�5]��N�3��P/�@\�#���!����)+����ɾ �Y��%�4�"�.בB"h�gXa�b�>yᖬ)e�+@y���ۢZH9�.�V�/�F\��T< �&*Ŷ��[�˷��[�����j�����S�g.��ٴF ��GH�v���Y��4ԋ��Ї����O�!	z�;Ii-��ɏ�=�,+������l+{I���v�gt8B��?�|���v\���?�K̨L�1��n�my����N&�g~&��$9:���evy
��R���ɣ�_W��G�A�b��,)\�W"(5e��P��3�B��w��]�rc/�Ug��!��3o%�����ՙc=�/6n�$�%� ����̏:�Ad;��S��ׂ��l�7o��Xm /������-0�3edxȋ�&�����)3���� 'N�l���B (/�n[���VJX��ږ]�)�}���mԳ����/�_b������T�nӜ�_�GZ�|���~� $���OR Y��T-"'���-���O9�av��ߑU�n4�{��m�N�(��+���))�'��ښh,T�4e�e�v#�("�XW�������{TC~�Nz��p�(��,a� yC�Z\�	���<��z(t�O�P��W�{5�}#��or>�j.f����h�7##�����n+�m((���D�7|�i��Sa?c�\����>���Ԧl"����pRc���Jg\g:�e�#���� �O�C��dV����d��2�Eo��c6�vXKC�"�v��]j�7o�䨍d)u=1c��� �
�ݙ>!��2;�;I�4��	�bG���]>��*R�Ee�,^��]縗{�ߎ@Kv������2}(�߫�:>_ۥ����� ���89:ԯ�d��T@dՌ�P��VPXjP�=�5՞����J��������"Ҕ�<:����������� ����p�,����PX[01�⑈ߐ9���Hx�PX�ϢÍ�!��+u���O������%ض�"{�!�ׯ���a���1�W  Y��,��ﹻ��KZ���.h0�6�ԛfE�$��	�C;yv�����uV�2$��@�E�MfrV��@� �5�����B��7��l�Q�Gj��+(��E�,�G��8��r<��ha9L�;)&���ͳ�3��6mrS�Бpp?t����3������
�&�c����C�Ti*b�'�oMb��]G*S��'���n�oP"����Y�X�p���ņ�S=���eL<�Ys����0�DK��1Xƞw�<(S�b��k���d�M�XRb��˥ H�v!����6T�-ڴOZ`��w(�Av�����	���ER���;��=#ه�Z���۴���K�Q8|�w���s�:�&�q[/ˉ��.w�	C4�2v����M���G�����x�i�66!p�CE��Ω-ۭ=�ی����s2��6!8͑!y�Vd!f�z��%,�y��@�w�/K���觛������w�5H�t�P�c�E��
Vn#q��=6��P��:v�ߘ,���fCD����p>^R2��LR��~��Q3���}K/^I�y���y~R_���"^�CL������_��N��$�}��)Ë�,������ȣa�� lY��n�c~$��10�OÚʼ�Z�$��AU
�� o�2���1W�_�+G�* �ψN��SK��2�,�P
�cnqW2��& A�o�s ��9�nҿh�$S�oSr𗨸	��`��JJ�髩3��\	�����q���"�0Kk3�Gn���X�<����H��	^��gȘKq�}.�ŗ���Wm��g�*9L)ߺ.O�Gfno§�&2��Hc����]xh����!E���]�$���G#8S�Q¶�:�1:������ R�Yv���R�������<)�v�*��������Y�]ڻ�|p���W�εKh�.��<>����hu9��F$���[�ɏ|p�y������c�sB2L����R�|(�[��� \U�r�u���+����C�P�V��F:(Xӱ(�~��ꏼ&����W̟b��pl y���q�[lJp.Y���d�Eyi�l%r��� ��`F�ɮcb���1��~�s���bC��
P��������c��_�?čˬ}6 ��R㡌>����Wq��Q��Ó�����T�$������Qx�m�9�'�:v:��q$����v'�X�Ni�}�Gy�� Iy�GxG!���R��=��۰!N�Y����`��maޅD�ˣA��x����\�o�R�Q2RJ�@_�|E�e����p{�DlS1���P���ny�����#��Ϡ���?e�z4(*�3�<�cI�h���M}�k׵u~/(<'Pgj"#�ωx+� en9m���nk��l'��š�X�4g<>}�ws4V�M��������َ@�	�vW~��>��M�%��;�yg�h/yLݰw��Jw%d�i�H��̴񿮴aQ�z�P����$4
*���R;>���{�1��PS;��m]V�|�V���voK�9�5���E��	����������/[3��t�8�C�q�<Y��>��u��w���{�J�F�n\qݖ��$�A��G0k~�o�;b;q�PJ���}��
@�.���&��?n�ɩ����3�C��yx��`C�*l8�S��#�e?\�� /l��L�YL����U���V�e��vක�W�M��śqԙ_M�9���>}?^q�9�N�|�@�2��� G)�i���?̋J�MtI_�~����a��q�>�0a�5`���L-ó���%���U��F�&ã�[Q�i�:���Rê����s�$�]�D���f���wI�΍���?�Ր�t�{e_�&�jv�'��:2����`�A������e�e�{%T�·��q�֛���O�5yc/~�������]�Ssi�����+����4Q�p�� �.1����ri�8�;���em�,��� :s;r��_�>�.7��2� ��2��E���ג\k������-��RHz!�x�̷~��<��k�-ɫ�n|�)�mI��@Bi?4a��Gp����P7�[+�֘ǚ\Z����Ƅ�� �Ɛ����7|1�q��V���.?�ii�d9RhC; t!���
��_����@0�9x��Us��������9ѓ�Mg���L���~����`������/4]+��R�!���_�FP�A:팓�/��_��:f�(�� �l�z��&��ש�B�YN:3>�,��Q~�9'l�r?4�ߦ8�!�:���̦a�%�Y3w_@��D>�;�[�]��
��p6.�l��3��=|$B[��1[y6]�+��̞����<ID�>^�>i��+DX�[Z
�)�%��YI-$��8T�r���Q�������ŃFR�?�]N������W��67P\�RT�9$��<&ߥx���/��!#ɧo�d`�d����o_�ȑ׍:F�̊�WN�h9ᷨ����4�гh��N�@�Z	U�q-I6�U�C��}Ł���O�84\�R�Z��A�ݷNb�aR6�M]g�М?`�O`�<SnD���{`Q�AbZ�Z��w��n���H�Ii�*��Z�"M�����R	*�w�<[�Z?I%����y�9ߛ��o��|�DL�M	54��?Ɵ�fb$t���!D���bSc�xծd���Puc�QN�/���<���,�r��������!

Oq B=Ty.p�_���e�]Ȉ�Um�	w���I�qt�/�r��k%�rI����H�w��BW ^����6Y��`�$3,�f^�@}$����P9�.�*M���/X���٧So�7J0��-�Z����Q�Cl�s=X�:<z �imp�I��&Ϡ�冭���F�C�0���
�L]����1p�qY�2���۽F�2�{�B	��^�Љɠ���c<xW��mD��p_6�h7��>=����݆⁑u�����H�6����,[�Q�,S��cR��=eY���m5eyP!?�ʕV�0ϱ/�#�w����)1�,mc��tJ��t�3٢T�a+.���i��@B�u�4z�p,|�G63������0��7��i��<������eʃ�Fr�k�G�[v�0]���'i˾����@%�W�Ƌ���}��M��A���y��R޾z��o�;" �WS�T�p��Of�@�~�+��,.��Y��+m�U��Lhk;tIc7C� HՕ�>f1���^�P�_���(���V���gz��a��J�~�	sE�����c�4������М���]�n��)����W�