��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�:߲Y�=��D6�n�s� �ܗ�3�*�]�Z���#�f�6�i��x$&3Wc��T-k���]��eY�
��S`��/��V�IJ��ݘW����S����f?^�da���u��Рg˽4�E/w�t��/�e�C�Q�̡�VD�tX(r���NKkR�z�WA�� �� �I#(��W���q�o�K2ֹG�P�C��@���xO�G�`�,���r-4��/���������f�&���Y�-�&^�E"h+�'+��s����7�d6���'t���۟W�3�?��B���E,Xo�D��"����4ƧՀ,SF��;o*�F+��?+�wvxXT��s>k�l�y���C�t6�HV#K�^l��,$[^���F�~��tD:��	z��s�i�ыz����b� �Mp����o[/��kv�P
4����F%)3C4q)�f�}^{9������§Vü�u+��ZA��Е�.�2ܻH�����7;�����?�l���f��ޚ=W�8��YRc$�F�r2�LP��0���G|�~�x�|a)U�?f)F��d4���K^m���nP��9t}��O�z��#ղt��}-hP�C�Nr�s�x�ӻ�J9���\Brv�³W��B0p_��*��:�+�.E\B�{�@v|qȏ QJ{F��`�Z��F�eۨ�9�&��JH���퇅D���x���=jr洽��&�Ɯ��k�*`Jsиӡ*�O.h�?Y�ￇ����m#���6?�dL�O6n9l>�3xɿ�����&̃���>�\�<�H'�0f���?~66���}�OR�X5�4/���O��o�8t��o6B���'H=v��F�	4!�69nCڱ����q���ɘ�i�q���c��Mdc9�[x�jJ.�h��������1Gf�L:���T>��\璹W�(/�a��z�F���8H;-�M�T�@-�
�U��]0�Ev��8v/��e�0Bx�@��|�L}���D{�Q/�
L}�Uɍ���^��������T~V"'�i�H�q��`;���==l���嬄\�ЁZ*�Ϙ��<9f�L��&�bأ=m%Q0�F�,hL�Dgp��\��� ��=�._f睅��!�e1�nG_M +�M����-:�L9N�Q>�e�[ݻ)�qG e�p͍sg?�U=���]���,FK�S�g�Q牠��G�ZL�"��'�Kr�d�����-N,)\�nY#���-�%9�E6"�v�ӟ�:s8���F8я��&W��o>�I���e�V
���%�jU�[�R\r�!��b�c��5���95��&	_����Yw7e���P�05���)�Ԭ��,�%�����@���n�T����i�K��y��-�H���ȋ�A3����l�&�<!ߩ�.����l��|²\�n����$|��������!� 38�}wd�2�~Ԏ^ ���L��HT�-(��@�1`�s��w�	�Q�z���Bԅ�;jh�?l���k�9�iqV���9|��.q�7M1��v��\l#�q`�?�;��\+�Ax*�����6�C�Hf�wT�iMs_��W�������^lo�~m��CtF�hQ=�=�w��D��z~}v�s���M@ҫ��,����9w������COx#�R ��a��͌L�J`�#�����%=�X4/L�w��w��Z`�5��]fM��;O]��o�-r�?��/N�2un��4R��4����VH�	��U�gY�\_6 &?���H�g�H��u2>4i��g,�I�? u&A��NQ%I�=q;����)��>���sht2�� ��m8	Ԗu���̘��1\�Hݛ)r�2�2�/?�����,���䟊�����k�4L��@�o��}!���\?��Tض����޺ʷ�@�#`r7>�ˀ㱣_nuvc�x CT�U��A�>ޝ�`:=V�SP�xo���FR���\�yoK�Ϥ�)=�>�(�-�^	H=�+�ÿ
��B��eҚ��4��N�[VQX�|��W�uO	� viz�W�g*hmNsxo�ZL�����Ĵ5&OV�H$��+GL4�v�d���?q�@X�{Då;�1�n��7�M�DJ5.,��J�<,o��X���Z�G?Hc"t���ɴ����폌K+7��,C�u��~��dv��7c-��̜������I�~r���%����INp}`�YH��Q)=��g��_ {��� �� 5��~t_{1 t��@ܬ�2^�bY�&�L�γ�/%s`N�'�����s�mp��R�8�*.�q'���\�F�D����=Xn�\1����P 鋄��p�\H�d��I�TTߩkeN�#��h^"��O�{�U��=.���.i0�&.HC�����n�AɜH����9k����8"���*��`�II�V�J� �u$CIcl��Q^c(Aew���S����JKQe2$�-Z̈��y�{�A&Ae P��G}��1=Y���[1��T_��;`��c5��x$��ʋ��K��5l�$!_��)"�"���d�]���8�V��F��E�#��AWGe�I�	��5W,�6��R�A�ч�|=���x�3<��p!�24><��v�s#lb�>4-�r B��@X2�h�[r����+�g���Ri��y�HV�9�µ&ALQ�d51������x�{;�$珩�=�89����Y7�����G ���C�X�]��Tȍ=e����Ne�1=��A�i[U�v�$e�|���k8�݄~rgC�2�K���s^H�/�"~�C��z���������g����+�O$�a��!:D˫1��H}��jqg�A�Y�E��FT���Kb?qV�	 W����%��J�&C-��܍f�n���b�а��-�S4?������{c����ޤ��u��Z,n ��F`ƍk���s���UQR�������ͣ�6���H�MDQ�Ō.g���j�ʱ�NBlv��F�t����Zd��E���^2w����wh������əB��D3�Ѳ;u?���V��+sқ��2������������4�k r�ّ~d��;�/�64׮T@,�I����[��Ί`���ju'L��"eĎ��%��@�)�	��ז�AT�����&�#�Ŭ���kU�2�l��y��D.���F4m^N�Yx���_�*�&��);@�2�='��h���K3	Q�G�-�;��p7S��;W41���%z���f����d�9�d�;8ph�Z�/W�e�YxL[2�sf���� z�p`�&��Y��'xE�.Ջ�����=3��;�d|���|ϝ��w�,i�������zbgls�Zo���O{�j��l����9�(ۍU�2�,�k�T��k�F��a'��4K厯5qb�CЪ}pZ�5a\���J#k�+c�`X+�{��½:�k�PrOMO��D���x����=�E������Q�Sg���X`��[}�lx�8�ܮ,�,T$�k���C?1�ȧD��D@�B����ߧ%�*��L��h�����t]�ǋ�Hmf��U�����s������ծO����q��୆������y�m� E�䞩��$+��7lo7
��0������˵�[��>۾��W��9����v�4#�{�-Qo G���S���h����{�=W�|����<�&�|;��(\a�2���ݱ�;`;T:���w��cҖ0(c���ϫ�FٳW����R�ׇs��)tE�漸
g�4���"�F\�������W�Yr}�;�{��D����f�=Q� h��Xj4-�Oqk/�e��5a�7i���ϸX�A�сE���	(�i���TkzT�۫�*w���t.���%��$]_��w�s%����^��[T������w+��J	�7c8�~Qv�+���0��?]��V�"q(8<���I&PE����P�Ԙ#� t��ۓ��VѴ��ۉ���c/٬6�9���:��kZ��������^�#Li�{q�����w`�~�8H����(z^z��tRvy��䲰ܲ�C�оZ�u:����r��B��*�f�O�2wMoD���R��չXV���/�Ng�ʫm���w���xP����2�D��)03PES/$.���b�!7D����kT�)|����r�'�do{�5w�KK��/e���w���;�	y�t�bD�s��K�߀��M誉L��V����iU�Qq^�c;7k�c�Y�ǽS;j�R����,��ҫ�����n��4\t��5;x'B��+}��~���}��S0۰�_�ٖ��*��;�t��9d�XP:��v�sD�)),>؂bv0���Y��p��$�3�Q:
E �
l� O#wW��I�%���|4)Y�B��%
;���e��������^T����_,�2p#�����R�u��ٮr [^o��1�tI���@2pY���xC�ؿ��|�љ�>����jj��d�o+�C��0�:t�osMLQ���̾9L�e����qm����͝z�x�A�ǐe7d�� TY+z�79Ap�&����a�E@�춬���=_�	���j0�>�΅���W�a�������� �d�F��h�$%�F�*Q@+�a�T��a����:�":�7F��-<�`;�<�_j"l�}�і�? ���5�:Dxk�/\F�Ӷ"��2�Z	L`�������4��_[�}l��l�>��k�iȯ{�M��Dں���凯�"���BU�[|"f�2�H����{�(�Y�!��hc�ZRz�N�Y
��X��9RC=�
	P�w뇹y�n��`��e������C�U'�/,S`��N�C��9:�犀EA���(���ɣZΙ�9L mntZ���N�P i����Țn��/�����������_k�7
þk5�gu���k��5P@�E�o�uIy����tzj[rq<5����
�=��pRZs�m�t�#�s���%��TP��bw�1�5Lq\,DJ[͋h��>�lE��yE���^v��������R� �f3QS��˘Lz�fxٸ|��q{�w(2�qk���F)\��u�o�Z���a��&�G�>'Ł���/�V�>_as�v�d!#����U�N	F�뵈](YJ��Uܰ�A:��È'.c�g�.��m�)Ҫ�)̖e���w��,��mf&K�)��	&��u�q�Z�ũ܄�Y��L}L�������P���*ʊ+�F�>�,ߐ�7��iL\WT
���k��O!��辖�&�]�s�6���&�Ў#�8��#��YI���j\�S�*������^{�
�Gmd`�;��^�L��/!��toe/s�A֎�>F9�����m؊N�� Uߤ_�k>,�x$"�}]�V1��]����Gݫ*t���0A���� �Ҭӝ�lע�o��~�#�w�lpS`�(5<%9S�E5�B���w�/�)�N�>��������'1I���>�k�eĄ��\���'�ݎ�������*�S`��� |[Ax3�rL9규����u���$��>�����I�.!�����h����kJ�����ٵ��5ੵ�tC&�q�X�Օ]T�-�K�,�!(��m�dh��k `s5�mB��cC,ؔR��ÜS�7DK�-��#H�xy�b(R�n=��@JD�����"��Җ!��M4��=�!F;$��. ���o�J֝f���=������p�B�cЕ�U�u��1��(�FF�<	<��r��W{W�_pPGK�ꇣy��S��e}-���#í����It���Z���9�T	UŇ>�z�𑨸�5-}i",���0<O��c�?�(��5��X�F��\,8���>4��p����5�.{�����I�啑O�Ϥ0<�{�P	X��9E2��ՙ(��u���;�Xǁކ�|��̈́���*�՘yƎ`����z%���B2�Y�aʡK���}J+�յ�_����e��ԨF`Z���<��C��_J\:���<�R*T���*�%��{�釞/>}�S>,��M�
�1�ԏ֧�$�wdYJ�>����,��:�T�|J���&l$]`����i����1-���ePӑ���_v}����.a�6[�L#��C����F̝�&_3ߌz�6D��<�[M�G�M�13���C�g����;SpԑG@=�&*���}a5�G�����o����1��d�{�u۪�0���R-b7�uq�P�7����YH	γP5�W�+}��bd>�p0|W��~n]�%nC���;N+"�>'�Z���d���w��l��|z� �6{A�Y&j���a�p_���M�s�[���D=��Y;�X�ƛI&L�bm�t��n���=�:����"��jH���;��0P��Ut�DJ_�f����If�7�L�Z�����pz�x��)#ۚ�e��q��r�3^�n�AW���S�>��M�h,����ѷ|&�ь����T�#����^��Hv��~0p�DyXK-.Ҙ-���W�J��e79'm���6������V�x�^I=�&�c?� �$<�D!���� ��r�j�vu��$o�߮��[�� ʟ��^*F\���ȗPw����
��l�k�_�۽Q�85�A*§Mգ������t��xn% ���>�`bJb�.�kh�s@���
)�n_��[~*%�uh��.K)��'��۶Md_3?�ʅ���YH�k�D�M�@e]���Ke� ��젻%RJs�풣]5��8E�Ic��Fx4C]I�7q�a�GP\��B��P�⶿咽�/<@��Ћ�?8����	 D�m��(�=��.']f3�yj�-�5D0T��=�1����f�j�+s�����{�O��KX9��n%��Z҉��{�������۝�[sf3�@�� rJ"�[��6��0��9I���B�M�ʉ�P�B�,�-�*�xZ|����o��/��u����RS/����^���&E?J{CBgl��BG��*�}"ۤ�zJ�MgA���r�����|�&�zL����X�lZdg籓:��v���MF�r�2gs�%�L�=�KT<Ȉt���]*+>Օ��G��b�oK��2��Q ds�h�/�q)ۭ^�`�nj�I�6x�����(&���\���z]17��n��%�0�JmL=��d���f�o��;[VC%/*&qzaf���m�s�����	�!X'63�#)�2W�N�z1nK���:۳d M�=Y��->�F���0
�]�D½_Y��u�T7��7���N
}����QVl���e��� uB��g��}�)���#1_��ۦ���i�������*���/8֌�UBHa��p1�]��%���6��tט(��2����Ȟ�ݫ�F��ݸ�޽�a�\�'뵋�J��2R�[�A
A�;жT�t�$&@��Y�
1#�iH��3��x��XW�%ٞ�;Qs���ҳ���\L�V�y^Ec�؃�nL���q��̴ \�+5�젣�.�\P��dH��5O��1��.�^�D���F�O� �~�n,W��Ƴ��`<np>���$��12N����w�-��;�]������A��;�4�e����a
�	�ȋ��p좷>��B�ũr̻q��E\j�|��L5o.�0�\hR�^@����O�E�~J��r��せ�l�j��:�ճ�+)��P������9rv��Ҫ�I��KzMT�Kݵ(Kl�&0a�&<?����uQ_R^�+��vJ=nlz��z�v�l��m�E*L�E���}q�Exʲ<D��7�A��ֺ; X\��m�z���-)B>C��J�]Cz�15�o�)Z�(���S/�zH�h�a2��f3N9������/��"��a�f����F*�_�M���v����� �l-��Pe�v��ѳ��1�v q�Q6�%�o��Be�t��z�����?E��oF���0^�Q>d�� �j��Ƈ0�A��C"/)�� ���(.��⍚+޵0$����(E5�����I�n���b�̥�fQ�QH�[A��^:��Ym���
�#6�ۗW�K���A�T`�e���W���R����Q�Ǌe��Q 1O�o��I@��DrU�������LSI>�|��b�=����y�h�%UgG��؛@r�r%=�qpK{��t���G�ֱc3/�lz��,���_�/�༬��KE�śE�RB�1�+=�ׂ��9z��v�r}K|�B�mA�̧}�]��<�;�r�K�%��X0N�)L����N �
��	x�j��/��3�r�����B��e��~�#� =�2p/���]y��ڴ'p�s���-=K67��.3u�τK�r�����ڹ�r���Y.��BQ�Zzx����e,R[�gf�,�|*�� ��&��-#��B\��k@mFP)��ߍ��o)�8�$MM�yl$�^S8�4�rY	��6xWm^�O�k�xEl��Q�i*4K��A��#
kc�>��!Ű�_�Ta����R%M�������Q!43Ϫ^|���9�kH����d�=��-��t6�wI��N�zǺ���#ީ����&��<k��0� 
�
��ZL��n�̴ 9o<��nG���2I�cb���z��3����e� �
	������.��'1�h^0�&�(U�/�6qq]�}�D�xl6����:���j�Y�}~�^$��H�Ƚ�9	�O�Z�����J�zE��γ3۱�q���?�c;�Vd�%tQQ�y  ���ѬJ2�F�����mR��b"SY�U������Ho׳Ex9�>�^=��m�����մD%r�V������R*�sRa���a����A��^L�π�R�#�ZP���0��M���kL�ry.C3a�`����	=���5���C�T�ӯ�$Q[Y��H���E�9�$�uf�]/2�+�g���n�?ڛ���o����?�_����8-ʸqJ��̂�o�yE&q����r	�	�����x5�VW-.k|ܹSƑ�<�� ��:�t�+�����l{?>��R�n5X%P�!�����le��5M|p09�ĄUIv�9ew��f��_a��5Ȱi�׫p�t>�~�=_�U(�˛��<��L`۝;�z�%���.6��M������g�)�qR�`���s���cw���ڜdI��|�>�������O!+�$16"'%��}�Һ\=n�	����a��QJ��Ooa:�\k�-����P�Ud3�E�l��T��i\�S�`�Xb.��b6��
�<2S�qB���V��=m��s<���}z����������'��*З�����'��Xvf�lNEТ=�O����d"
��U5J�ap�m���8��]ܴa�)�B!�5�d���R�t�.�9�ո��~���Լ-?���c�H�LAW(�6���^��;����PN�_|:C4(�{/Z�R4-�m��*���n�	*��� �a|�����R�X�'�y��^�)�iĪ�Q�'sut�l�Ɉ.L����c��dnC��x#�ꎧb���k���g���q�m���=� �`����oL���TFx�6v�+-�b��i�$1�C	���u�<+!��"��~ ��of���E)Q{F���l1�g/�ʯE�_���"�4��e��C+��ab
E[O���`�-y�љŪy��i���M&R�>,�೷M��k�!�Ѷ<oP��dȣ�\v����kv����tVy}5�kKL90���L��$�a_�Κ:�^	.G��R��q����ү������u�S��VS�����Q4-��\#8&!��\(�*O~
�".���jk�o�:�@r��0=��N��l�V��{��{����!/�n��I��2{�����,��z:�%f��������S�����6{q����t��;`��ʩ�z����������3�Al�Ӭ�J*������@XS�:O�A�F�%�0����`&�ĕ��˥)�R�e�&�R�o{��m��}6����ji�v[�~;�\��U�!�:S,�ˌ3Պ�$�fi|N 
�N��V��
�7K�ZmN��z�E�a�j�a����U���;E��z4�S�`�ÍS� 	������	Wqٶ��O��I'��1Ӽ��>����@�#��T��W"b�i��{�2jķ+?����a�uH�֢;8�)加�h6��(�wۢ�S�G���:���/5tC�'�Ӌo�3�N�Au#�{	Q:�v��u�wh-A,��jcz�{�G),\(���L��o��������;]�8���8�(s҉nE�ŀ��--�_�����{J&�E�"=��D�2-,�+���~����Gy<����(L`\��	�;1b�:�Q;�b&H��B��^�����T(���銼��Q�7ݬ�^�h�� �O�ګ�E�Q|�,,/N{�w�l&� ϙ�t�����Hļ%�+)���@�g�x���M����5/'�KqFj��W���
���S���b�8�IQ"���l���):?�'�PiA��W+~ԞD�ݹ5���mv!�!�WI�	_�ML�Ok=�*�u{.�����`�����dv��}m�,bO��~�D/��)E1j�^=���w�A�7��T6�0y���[�QtZ3�~��6�Z��-o��˨���G�n ��BHj�V�֘�;D��w��_e?�'������Į� 7a��3{�<U�z<�<Ͽ+L�_4��5W�� \*̰�2~-�jsD+��q���\;�=����7��q�p�%UT強-S�].C���*���aPC�4*����H*{���Y!�piZ)�di;w_4�q�qB��6��-����A�.�u���~��@�E�"4�	��<�-�]�*RN]��R,�������}�R��}k�+��53&��v�v�8�;Y�Y�L�f4f2�^j��6X�~c�5P�7�\=`�i?|��{���w��<�����A���^ڙ��W(u�6��J2hac��x�ǵ���%�?=u	�ˏ�8
�7��2����ch*�v$t�*�"4�s�(���8TZ�j��kD�v���#�64� ϕ���GTd��L����E�5�f�{h��nym�3}=m�*�����>�oS�}���1���A��(/����|��\@�l'�&@WO�؂����؃�Dy�!��U�ҋ}���(�jUi���\��.��+ŲUk	�3�N�z�Eé�ХCO��PT��]���<_��6������Y:IZ�0-SB&(Ç��\��>:��~�&����}1�5����pC�(f�#�d]ݳ������C�Q��1�̯2�v,�&�X�Vs�Ok5����r�O��EAkTQ�~f��+́�B����
��J��4Q�J l�VG�̄��jN����b� �T��QR�z��v]g�v�y�#�!�P�CU�͖�k��+���a�y��Y�,E|;/'=p���$��E��ǒ_t�Y�N70��_�6>6
/&��Ȼq�]�\h���=ٚ^S [�m�;]�3iR�8�' jU�`�d.T��t'rX��hč���g���_��O bn؀�~�U=��f��U�X�s���F$��u96>.�Pn�����l*4�<�a���N�ۿ���H��@V���mcH����!y�����b:p|��WWR���
�A�Y)&����l�ӓK����0�[3:����OQ*���dqδF�X�ۋw�9u6P�y2��z�l��)l�(Ҧ;4��c�湟�B�X����e��+Cl�g�VΣ�Hk�R}s�����>PQ����S7<L4*��?3��2�$��T�w��x�J��7�5�x�^��g+�#�m�pAS#)[�l�G ����o�M(/��X8��Z�LsFN�v���x��VҚ~�t��\�F���l�Hi��mT��0L���㴽d׍�k�����e@����%�@@5ffv��y?�[��<Om���B3��7��7�M^F����s�(��͞�u� ��{
��i�[}6gQ�D�f��_�+�x���~3��R2��SF��������x<�R�I1>w��?�Ɲޱu�3��'�5*�u���)�=kX�%<���b&���$�Z���_]!�,�	�>�ĸ��v�ێ�$?�m�I^���ĭ~"Ury���~���6`����:)՟���j����(Q.k[��y�O�
�U3� �����6
�@k���DF?�\�F�0��높T�<��va�=\e��h��{O��uW�ơ
^��#A�e{.��'�~���h���3�{J�c����P�uL����S�/�m(��)���Ȟ�7��xo.j���hN����c���uz3��:�/9����Ҕý �j����������������+����uvׂ(e���$�~B=$�wŢ�]�8Z+��k���v<����.�ע����~l�R�?����@����ƈ�-Q�I��O��E���k<�8L�YώTBʚ7�	�.讚�rʹ���L�H���1�����Y����Ku��q2���s��wxH��E>.����i"to�:{ .j�h6����Qv��?�6H�Z�b�x)�{���-���ccW�&�r#3-���f���mWy,��׈c�WnXiy��r�B�T�YP��6�a�.�'��.�e�w���k#��N֡�V��8�y�p҆mq;�.lJPR�a�����Ne�=�h��h%�ڹp�l�����A���<Q1 3˂34�܆'l�%�/NH��0�ǹyJ�N�_{#��]Z
������S�;Rb��2���Aר{��C�~o�f�+�A�(6�{�%Y����orH�E��;.�%S�8=�h�T�-�����q�T�*]J�ռOX:�;�]C�a�7����Suy���xa�gPx��&Ҧ�����ƅC�\����K�4�Z������x�W}5������vy��_�lȶ&��R�����b�޶9�%�e�ۚc�D�E�<#��=(ͩ(,��D�Fb�Z�<�d�\�J�5���6^Q@�b�s���;��ܘ^����99	��E�fP���RB�������䩺�UI�����W�Q�т..bv��|t�4�n�Gf(+��ЧM��.N�CN@�"ś�=h8�;��H^)E
-�Q�@مK��}yl�['�d��CO��Q�\
>�&�d��l�ҍ�)=������C&fwwy���´��!���ॽ�j�3�����	��M���4�GF��H��yTU��k�w��p�Nr�5�Y�ة�/�@c1��K�}a�S��e�6��HH%Wv��V����J@0�'VQ�&�'���6�	/N%f�${��j��2�V<����lf��+����/�U�9��e�/Y�i{�빹�T�HQ�}�f�Ƽ�v�ҎqnI����u�'c���L���&�uF͆�8d�h`Z��w*=��o��)<�7u�J�oG�9�l�V��L�ێ��D��'��c�'�����2g��qLao�UTZ�nWwB۱�d�nW����I(�{.�mϱ�g�	�^aܿF~<e��z���Zf(����"�Ӟܗc���ZUS�G�-���M��<5�����E��0���9N�w��y�e����B���5E#?xj��ӂ9=jQ24{+R3�G�bZ�@�d�4��"�F���@���3v�cC*n�f���pڻk�NJ-D��˵FS��2���^綆b��K�y�@�ɖ�S�b��g��3�  ���M�A?��?V��������B{��HH�r�+W��%�;9�l_WQ��̫��#)�g���.���a
�=вd�� ��m����t��S1�� Sv���v,��B���f�N�F6d�ݻq,ҫ��	��vI#���w�S���pɝ���S�S�����Ujzf%�n�r7<��ݻ�I��wwD�l�	�����U��(�����G:9���}���j���>�O�Տ]�3ŧ�c�c���Ҹ�4�}^A�����0,���D�-]2�
1��7�4�_֣'R�'���z� ���T�-����>� �g�1��OE��1���z\jЍ=���+g[e;u��^��b�����.t���.3W׋��2��qfH\"���B��W�rG���#jpQ}��Ut$��޴�4����Sӑ���:E�R8����e���'�b�����DT�l���<��<��L�m��J�����Iط	}��~P�����S���ER�M� ~ċ�/��������U{9��~�u�Vi��k���1-e�Y�?%
�K(��oq��򙍬�ǳ���Xۄ��2-��a�����7���O߀��eP">2@����y����!�_����[�m��!u����P��-IxoE$�����WD˶����2���p�MJ19�BR� �ۥ���6��� P�(����}�=��-#�S֯\A���k�.MXû�kQ�9[��P�dx�s�HzP/�d|�.�6w�z��Y��+(�^�� x�!��H��Gyc����q׾��^���@J̘�ĩV�j�zԬZ����w>1�I�K0�Gey�Y��Ĕ֒�2}�nD�w~�9�������ʅ���*�������?k�0޷k��&���d�hK�.��K������Ap��&/*S{fQ�z�͊�S�9 ꆌ����7��>j���A����1&S���M�ϾN;����r3I�{[-*Bb��m��C�i���v6y��i�ᕂf�1�>�QM���ն=:�I��y�T�	���Z���TN���EC�Y����q�9�Ѥ�i�PY-��j����/3�p�';���Җ}<:��#�(&�I"�Fo*�dl�H"��^ѭ7�����KP�`���S
Y�����i��~�P��V���t��Z%	e�a@�SY�{��$;&��*�ρI񛴡�E J�~�%\��þ��]�U��L�awQ#�芾Rja\�������7'�B[iZWKA�� B ��L�+��5���j��(b�xg�kP�/�2>^n�Fo�S� |��^�U@�����g���{�?ci��J҄�d���˝�^����J/BV0x�%�Í��} (G���GJ��&����:S@�L��M@��T��d�3�1-���7Z4��zD�i��p��vw��B.������im�&B�q"�xu��7?	v���x�+���:�C zR�|�
���h�z�6��g=෪���� ' l�%�0��mV�LH���7���ޗ��8��������F���9����"ck�� ������\��K���b"Յe�#?��Ry�']�}L]��xe=Y��L�#����S����/���7��r�=��:�Zɍ���i�mM�0ӄ,�g���nE!Y�*@G�ja���=nK�H���KoS/[�$,��W��n"7��2Y� �h/���q�6"�$8� 5�95����9���<%�Z����"Msv���kN����h	͂>��s�۹�f��1���I>��l.��b�-�W��]����Q��/vLD��h�=*�vS{fc����'�\c$E���h�����N��\��}��&�sJT2�m��� �{�J�'�#R%3~�Q�ɲB�L�IehE�)%-�[�����f)�������/z��cm��%���.ߕ�"(s(,�A�z�4?�^�v�����v�C����n�DL�qi�����	jR�[��g�I3���%r�z\�����5��ܺR�t�����I爑=_���7���FK�;,��&�1�t���ƒ&+;8�T?H������M�]�b�e|9���G��p��O��vr��d�r�F��w��YͧRex��@��#\Y[�m�E�+0Vf�D�ʘ��>�[�{7�*�_qT��bY�mZ��k���P������]�*�Ak-��B�I1��<Ӈ�D�gx| ����ޫ�T��J��*imsZ��k�X���j�ؙrG�}ȏ��kk�Z��v���N��*�>?> �UG�j�	l����h�~n_�g�`p���ў�m���2��a��m�N�PO�u���O��!\^�F���r���L�� ���B.��(܊L��ܳɶ��5:yfF�ϝ��	m�����:N�jt����6	:�ER�S(6�t�n·��@ʱ�����=��E�i^�`gf��]FJE���E���pl8��y��1i�[]���*� ����j[\�;O9]�fP�St��p�����!�w�J+7ӂy�/�>:Z�]� �X�+��8�o�c�~�Fg1+�.T�)vT�a��;��sJO���
�� ��+)hf
��9�/Ǡ�e��Qt�u")�[��0a�@�K�:��FӴ�x��sȃȝ1M�-��h��������X=�mP�*�3�`��&N�����+;{��H����';n;�O�k�70�ڪ B�{�"�#���u��$����/���<���
j>}�o9+W>�&��~"	<�N�w�||IR�}'��/��sl��d�Y���d�Ǵ�0�',�QQm���n��oK���4�­�br��c*̜ͨ�-�!JO�p�p$�n�=4e��7c��l��)3���=h�Uf��N��u�W�:�V�xb�X���/�!�m�#����/��L\��<x�\<�U٧xډ�����Kؿ꜃I���75$�i�8��VI�Ko�Gi��έ�-XF�q$(8/���ܷ��ĝ��2$u/ZeQ�f��}g`�Y���[�N^�QS=y��2��ݨgE����Z�*aw5�Ua�p�{7��(���},�� ��@�+T�5�G�ո�N�R���o��]D��PPUb�%����q��@��<��?�|͏�#�	2)_���i�7�ɒ<mף���-��qs�DN���f*�HݍkŦ[3���+s\�x�|��ڵ�s�����%�G���0�s��[
�3J��<��,f��iS��;4*�B�*���=習�;W����o��$��udv���W4u�1^�AY`�dh��C�35�T(M�[-j_Dv���F����떹Qd,~�=E�Y���x+�%l�=^��������>�V���A�?Ebr	I���6�<��z^���]#k����������[�,�J�T�uLK�C�6��j��Ba*(F ��aȐ���{��D�h�H(���b�u���.�w튆���^����e��26����Ǆ 3=4��ˋ�8���"\�f<� �b�������6�vʖ��uy_����v֩��8E�=�R��bƾ)������N�"�J*����p����� ��7�q�;a}B�,u�������x͠�V2*����r��z�o�uu������2����r���_p*�x�O��j]�#6������z"���:JF��������(�\V؄���v�.4���M��=�˥%����yn��d����nI�Ƣ���l㠜@��\m�ݧ���~:��n+�T������/�D,�8�^�ۡ���Y>⵱T&~O�r1G�_�^⓻�~+2Ԫ�}Uia���j)�Z��+_��{�%�]c] ,,�ȥ��Ƚ�c��G��xJD��@��;�����;�`m�6D/U	g׺��z��;`�K������\:N���)�m�	ȋ�T�SP�[߰Y! ^�vWV��m-`�����Qrx�� T]��#VD�=�v2<z��R������p p��&t� Bf�w:{YB^���Z���y9�So!�������=	�+ݶXa���G-�v"����K]����?߰^ ���f�"x"(�Xr����`�t��b��*����� {����ޢ3y�e?X��u� R\���%��D�Rt~��bP����Z_�c'&贝� �[
cn1�-b��Lʈ�js��1�$�:Lp��8I��4����2eA����)�\��4���Yj?C���<D�'":� ��Pz����R�i\stFh���VrWkz�-�n)ﶤCb�S���:�5I�Xn��jy;��J�|�o�f���cGyBP��MP�֣7�`���'���"~�~Y�H��7����eU�X����Q�A�ʆ��������P�W:����נp���h�҈���W��+J+H��滷`Gz{�"ɑ��Ȓh�*l�~.xD�ͨ��j��v�_�0*���R�@����_��&>��5X�[� ���sK�tK�բ�4;c�R9�z��#��)9�&�:������b�[�U�x5'W0o�u�6"���#v�h4�/��DL�^³5�[W�T,g��瞢A��%Myܨ�4�E��+���$L�z��+�ʍ��j�-�qptj�DT:[�����F3��n[D�i� �!��,��~���	dЏy���s�Phn:6��O����Ae������a �m��k�R�6W�^��,	���%emy\�Ӭ�T$*/d�`g�U8�����Y�@6bMr��
x�d:�����J�1�,��;~9t-U#�s�����!ڜ�v����y(~�ޢ!���%f�P�[TO�p����X%�(ktAY��0�H|lP���vc�Ik���4������Ud�g9�ҡBd]X fH�������꿂TA'�.v-�f�S���84�S{�lE2��C�6z������Z�:j�F���5ye�D�k@�j$|��j�7l�~tX�%T�u��4��M���.4�"�:��z������h��WA�v����O|E�!�|�>L`G�	�{,��;VYG��_�y홄c��yG��P�7d���'�eFIy��jZd����;�<�Lc����U�N�hx��Qaa�vw�f N����d����E�+X��z��p���:�@�_p/xֽ)oD�Oh��
[o�ĝ��z��!�\�0Q�����`o*��C���Up�3��3t�v
�.�#���.<�0v��N�lm�8�v|���ʑ�
��G=���&�����V��Ɂ63n�7 `�r����F*���	����)��a�L+<H��������f�K��gK8.X%`����[)r���ky�g���u��<����o�w��,s�C]���$���vݿ)��4�Кx���u;�O�=I~�X�1HR<I�I�[vl4p&>K�4�$m7��X������E;r	�ժn:��j�@�D�"�2�q7�1�$��t܏U�:(�p�S��ʤb+,�G4�|�ߙ�/k�g�e]!�"����E�=ۗ�et��+��l@�RZ�JKm��ȫyQ�pD�
�Ĉ_j�|� E�+�ɏ=�����^�݂�S/�/����?���UEL!��x�����̭u Y/y�X��栫��W�	�����;]4���|ɩ�@���.����ۆ�P	f�v:\;�St���_{��4H��S�y П\��8��[�k��b�Xq���d�S�g	`Q��SAF�m?��KL�5�V�_��ά����_�|��5Z�lJp�(�ji��;|��4+���"y���6tF��e�v��S<������-�����`A9��e���:��$�z�Rɛ������8�g~��@'-*�1�	��hdn���W��A�kٍ:V}�ES�C�J"�`-������'93e�_�����.�u�;9��شq1�Ja�H��&@`�Ώ�5���N|h��^�󬅁0FBb�3�U��E�D%��,k�$.+3�2���sD�?'�6x.��m#Cݨ�[k�̡Hr��О0��}�5@+��Լ_��xI�W�3�+�1G�eB\uE4��Z8��Hz����_�@ت]7G������o��ְBK�/i��5(")!?�]���6���T�~ґ���U���8h�g3� ����X�q��}i��v����G~��M�H��a� b���� {hGj-�о4�rc�3�$4�A�aR=uQZ�q��l����⪼:��Q&��-n�a�-�
�yNNy9@�}~��H`�, UP������L}��(ێ�մ�e�&�|ݻ�Y��f&8���KV�a
����+`;��H-i�+��4H�%�\�L��J�a�S{�}�LA=�2���C�1��ĥ$ыX�\y&���KF��:�:�S:
rۢB`��aF:��V��by4j���Z����ߝ3�		e��ĄƼ�ȁ,�$y�m$�N(�*�R�:S��v_�#�0�0�T�0��O�&#�8jv�q���l�})�2s'[2�@�&���kA��0�����8R��k��u�s�F���Zj�,�7J�����Y��3w�Ҏ��N�<��K�	O*�-?\Dk㪘�%0��vh����o_��X���Jq=�j����H	k�?D���I-��]�+11���Gm��`B��?6>]=�O��RLK�`0�t����@�I����.s�h�8�H���.�0����+g2F+���Im�ۈ�P�O��w��^�K\��8k��r@�s:�b�MiQf�>�^{�=���f	g���3\>�6@�K@�W��x�.�#m)G��6�XVE�7��!�p}|�FbO��aR�<\7yn�H�m�r
Iu�<������c��֊�wcV��s_=YK��!� d��3���N>>V){|?�s��t��>y�!���=�И7�]���QoH?���	��a`�¿��X��qs��m	\/�$!1��9�tC�����Hoɚ�q���0Cx�Qo��M��Ⱥ��V�i`�K��;���Z���Bբ}J�s�+ڵɮ�+?���n[M�7J=m@+�I��\��Z���[q<>t���1B�y������ȜDCaI�K�0pP��� "h5K���l��ӧz�q%S��ץW:+�=a|ٝ ޡ=�U�ߧP:�	�L�*�^&�E��m |��,SY���u+��h'�\�"�t�\���h!}�(�Kf� ����<%X �d�k���m<st��,�M!Xe��*o0s��1���8)6�NG��oX��cI���N'ئl�)�7�.�?@�ߏ��y��O�M]xb��s�ݰ�����nek�_��%��^{j�K�V>K��T�n���P�n�6g�0N7�!��Kԓ7��lj@k� j�D[�?2�&
�@M��V]?����,����\7:��y�����k�tp���^���/�':��3<�O �ҵ�@.�w�B�����s5?�d�s�ů�(�>!�8B��{=Z2�G&�r���y��!b��o�1wz����MvQ�_��������lC;����5Ei�bʞB��2���M[�.^2(5�=�����Ҹ�+ �Ǭ[!0���s�4oV��b*cKk+FK���f�V�@�6��lt�غ�QuE^չ�>L}��s��`�{���#�xGc�6�k�B��C,���lť������]�*����2�B���M�E<�Io��m-�O^("J�&�o���NP��.\�|��.?'�a��P��p��H0��v����H,�ÚMH h��Ӄ�nІNhѕ�^�C5�bE�4 �qax(��TW}��Oz��Yg�d�4IqFaV�!�C �]?��4n1�n��e�p�vX�%�W�b@g:qye���MJZ�^tTI�~�i��)R�,��t�/���")��~Q,���F���l�z�������60�rG������`TvԞ]��ZJ�s�"�vE٨�����&�CU���y���Jo�DSL��&װeT�q/dc����8B��qf��l�3!���F�9YN���MY��J^��j�o�,zy���I��=~�˦����nŦ"&��`�	`0��5�n�7�y�� �$t_��V3���
���P���V<!�v�իt�">�"n�ܷ���)d�㸼Q�O�7 �Z�X�/��؆���Gf�L=�#ԛ����R�1T����=B�YY|��oJ�5<*h�v2��3xC����D���OF�p"� �q+�
�Ǧ*���K����"F�*�sn:�����â5�Mk��[;��p�S������ѯ���C/h��X}��t3~�C�C��oL�>�q�)qW���VN��Z\9.Q�:���z�7#���uj��dX5I
��[�v�x�?�0k�0��d���0�Zb_C�9����mi�zn���n|�p�/�qW�(��������Y!��9�hD��7(j��7�	�v�ڨ�:�=�<��J^�iz24�%|���i�JOYc#t��� +�:���4���b�1�p����UA�W?��>����������ӕ��UU���^��F,�k��W�c�@��G A�N&\�2/��q�E,>%��,Z<�Z� .�+I�H퍪���
O���H��G�h{��g�e͋Ja����g�8U���}�v��k���{;׭kk�5���ELJ�X��'<̂/p�fr�;I������ju��?�٩�q��ɑ��f��(U�p�#2-@j�.P�i �ڍ��S=l���=���z�?������C$�¼̓A�i�I�C��[�\���Ja�%��ć��DP��H3�����\�gf����;rKү�QX����3��]�&/�����0�f-���t"@��5�IL	%դ���U�/A�0�T�)������I&h�+��&֘���p��Q�m7B1��Q���s����5���v�~�f���*F��:w��`��]-��oW8�%���H�9���2����9&�<I���pq���Tk$�=��
`��8��2��P�o汚%z4�<�'V ��2YQ#s��Y��e��GJ���>ƏUPYT�m���*7�wËm��upn�`@���Hv�!�x�?�j(��p������ ��G$'�0au��G�Qf�<͑�Wpÿ�/�hhU��|��V�?C�^r܈X���,��s@çXK����@� R��<�}�7H*��zb��K��[UVլ��:b��Չ���-lu!s*'�@��B$F��V:"����e�Oh(������/�EA��]�Ad�|hI\U$E}�w�U
��A��q�curm(Vm45��Ri �]�FE('a\L�J�_;�V,�=Q��a�P[�|���t���GP�of$�	OW$t���
ׂ�tM�,�#��(��<r�͉�#�®A;���A�����oU��]��-��o#����[͑���H�Oki�M�n��>�K"���Q*I=��H���Ǆ́;�/��bҀ�:�6� �A#���]�}j���a�[>�D�L��p<�V���e�Z1C�Ø)���Ǩ�+�:�Ϊ?�OC��	-� � }�&<�:���K���'?U�[l5d�H�lm�� �8�ɉO?Mk3��"4;�i�?�H[��ϵ{W��o>�5@b=<�` \��I�/IA�CPdB��YMo���\ai�A��H�{)�����aN�L���ۻ��#�^�q���W���T �����nއ�� P�+���2�y��z/���&&�)���`D��٭�8��O�lRo�e<��
\>���,8|[���:M��]K��+׌
�>4�I���k|�Fnk�x�}��f����I�{6OmI+?��ah~�����LNC�d��LX�]Kӑ0\��Lƾ`�q@������ٺ��`!�l�S��m"l��0���Ǘ�El�¿z���䦥��m7��B�|�T���>����4���Rp���놕X��H���X���m�K��.D���rg�<�'�-����6��+<c�!T�e�`�B�|��o��L>�����j���&%l��%��*b?�	����G��WY�Mڗ�U��}�nQ� )F�'�?��B���ư���&a-�ɀz�������!O�^�~�p�c�4Z�!��u�P�`#�#��W�wu�9�W�c����[&��=��.p!�� 5NA�Fs�X�,�+$\����âr� �n[חh_��"W�0��p�T[��=�]�&)I�����^�s("0�O�^. uX���!��Mm\�O�<r�}?Ut�x�����Bٸ-&��,��q��m��+�X�M<��F3E�l��q��`
F�v&���=pK�]��l(At���v��ݧ*���t0 �8"��Q�(���)e��d���5��c��R-���M��jm���PV/�7���
�;D[�+���ג� ��%��ٶ6���~ɨV�Jǧ3�p����<jZy��Հv	��RS՘��a��%��w�ȯ�#X=A$K3�'7����Bi�`�t;��ۦ�� �=�N�{��0)O�E:6�'�g��ҭNr4Aep�I�-s��ƕנ�=F�a#��{D�o*��Y����w ���>��U�j�&!MNzLge˭_��Ѷ�s��u���ڎ\��gekM�g`��T���)俴s�;AB�=�g�'�`�a}�\L�����g�us �{qM]�&M)4��;@)!~+�xN��J���Spʹ�҆eR����{����[ǭ��Ɗ�%'�QCl1h�u�r��&E����1�\+��>�T��¼�]��U��ɢ����;
P )��+���PC1a���QA@��PA��PC9c�����jhΧX�?�!4-A�4�A��:+	S�:�qك�����<p�]�!ߥ��h���X�U��D���{���R0�����	�NA������Y��H�ic�VTZC�fѪ^�e�I_RC����1�q�4��w|�=;�3Ź�z]]i���`�6�(<D;��Ed#���](R�)�e����Z:`��Ѹ���'�s�M��c���)қ|f��	���N��L�֍>���W����R@tp �P)�KǾ���nzM�L�nM��9�[̢E>�Ë X��{p��o��6m�|]�Z����ca��(gi�] �Wd � py��B�*��,q��h�]�ɌąP�&�&��=���-��-��3�>G��1NYu�Q�o�c-���J�c���G��5����BiG��{{��:� e)�SYſ4�G��������>�Z�}�J�z�U�_$���b�q��-w/5��&]EGޘ�&���S#���	����l���!��fr�=�@!��ȑ��(CK��x$dI0�-���[B�EN�RB)=�'�z������T��Y���Gq�R}�Hq��
55x��r�lU�>�KvqK�?՞���!i��ZLn0���D���şue�Q�S�W'�͘Ef�/������2Q�����D���t	��z嫂G�m.`����:�SaF��Y�A5>x&4569�]b�"n�B;u'	J��;Eӯ�ܚ`�s��ۿ����(ߝ��}ë�w�\���0!��V�5��xPP-�i����'ל^��fi�b�s�|� D�ȉXiX9����A��}k������X��w�����;0X�GO��y�l8�F ���Mjջ����V������PRLuu;���g��6��ʚ�+	|E�0��N �>ʪ_9R�Oh������Q���~��k&P�ܵ�<��A��%����H�
'[�ҳ7��z�&_FYBNucm����ybd�Jo���wYJ�����+�S��׀y
�$�u36uUȒ��Rf?ٲ���/g�t��U�������[�y���$S$Im�P�.6��?ȫE;f%'��sN�IMs\7U�$����c2'����v&h(.��_�8�P2f�/���tB�e�P��^��x����):�u�5I_!�W�����F��~p~�վg�M!PP��ꣵ/��K9�$0��&��#;�4|z��
�':a�9��©hC�9��z'�q��R��������\�� ��#_�ycڈ��S���,��l��t�W��j|it2�g��p5����*��L���։�*>LL}{��](�vN�3<N�F�pj�ʄ##
���(����J�QK��^��_{�ڋ.��Ns���Q��NtUbV�����u$8����W+k��:h�ɴ΍Pk��&Y�.�?�ߧ]y�<f���0:c{s�Ӷ�v0vS�W_8WM6�b%���?2p����@H��6���������@��Ʀ����d&�'(L�KBv�áW;;�������9�a2�=�C<M�+'nW���AcjK�i�`f��L�<�9~�>՛pn��	�-�U�g�8a���ܪ�RDs�w��B$1|�q?�$����"d!�{!"lB����wu�m�i^d^d��XyL��m�ٯ�#�_9#<�d�>��Z~���R��h\eInP�ơ�J�H�a��W��[�a�<���3�Sx�y#4*���QlKַ55�*y���`�����M�:�W�,��ǕR.Լ6�\|�������}�A"�WA��ǟΩ4c�:7�Z�M��ȧ�����h;� j������qh�Ÿ�W?���=_M�ɠ�����~B�[ݫ����4��y A�����Wܓ���Գ�U�	� ���5Y�;d�A
{���B}�U+��m��Íy�:��R7�p����\h��t�/[qa�_�ǱZ f�8��5����㿪}?׃��-����8�Y*�7Or���o�ۂ?�<P<�I�Z�{�h��}��S�@m����5�5pdH�}�5!P�}X��	o�l5�]��e�w�����+���K�#�!�V}L�N�Ä3	ύ��\������z^-��C`� +�D7��8{��.կP��Fd�
w+�:67_"ҕġ qjj�p5���$�x $~A����-D.ޙ'7Ş
�P?-��Ƨ���C����K��I�aMnU)]o��1C��9�sd�����d��@W94_�$ȹq͋�^��s�/�e�Z|��S3�G]��5�!��gdN�Jh�p3�@E)_X�]/�n(,YY�E�d+��8<�t]�?Rc���5���5�,���(��[�6�n�TґG�'l��L��?���}�J�j�8�r��˻Zb�mb�����-�t�����P�Oe���_��h��]'�ָ����9���3��#MM�?2n��2����ޣ��A��k���v`C���"�7Ф ��Mi�1��ҫ�!Iho�82(��%l.~X�~r�v#<�Q2�ѿ�U���Z-�x��i&�]��~�����~��B�~����:���h�p	o��p��@�R.���_�:mz���?�w�N�.�nV��s:/�Φ eQ朸��Yp���4��Az�a.�˞�y��n�v��g�Q*�ն�X���>��_����r����R���k�ꅫ��R������P͆E�̭f�H�k���ρ`�/�)S���i��5B�j�З5�=��k&���5ja�3���C��B�_d4�����jE��ٟ(����	���@�!�V��1�÷D#��K��*Ħz���.�r����8E�ӣ�m|�ͼ9e�ڋ;�Ŕ7�1O�fw��Y'ڕ�=��~�9���x��{�d�k�eq�)l"��L�e��].�qY1JEa�n�꡾H���43��&��[d�+�y~�t�/~����Y�8�BDiۦ�R7�ͷϾH��6�#�j=D�c�����]����	�}%����.����=Y�SM�/�2{i�6%T�6����ӛ�X�� �Q��@����7�.X�Yi�9��T�����@��y~������J������^n��
��ݜ��B�X��w&F��N�����hzz�����J�t�^g��H�Eq�.�n�7ǵ����b�����Ѝ��󰫱�10tH��-��|Ѿ1E�r�P"2(M6�xe���*iB���=Xx���u���+?�8.X��Q@y��#�@?NO�g�J�1Үr�������{f�F6NV�|�Jz��MӒ \��&���D�.� ������𱤚�zc��^C�4�dr�@"�!ڻiʟ
��m�A�8~�;��s���or8:�5l�RRvX�E��`�M}�.�/��d2VT��aj���Bm���N8�d	�k]Qqm1����"�N��i�`�Le��"�`�ѹ��D�#_y��z|�-a-}� �9a�k��M?C����I"{�|Be�W�c��j��w��j [e��_[�R�E���X��"���L3�T�U�p����W��@��׿�c0~	��*�:#N�:$�,�?h�u����i�O\�mR⚦�jb�䨬_�P暲�-��%�l��3@��֖����K��>�)6�c�n�]Z���,��b��˻y4���Z���7�$�|�Zg�ds���X��7,�XRW(����
#���	��:�Dғl�kN<1�y�~<�'Ժ!w�9�����[n"�W�pp�^��c�UV-|!!d�?�ؗ#Z,�)&z %Yw��&Tl�˗F!���x ��<T-P��
Y��re�����E4��~W.���ι�as���{�c�6]"=���$��Ƹ�)Vk�)�{�9��`��;�g��E[f�1��趐 ��
��q�� p�9k�%�R\�~t�;�/�tL��X~��*�|8R�ŏ{�zU�S��_rrM�t��43���N��b��ʐ<�WM�Ë
�A�m��g����`Q�p2���
�!F�_BI�l�
�"MPp<�K}h�g��%�lv���W��nQV�e�&XI����x�;ѻ>+ADn�ve��ie���FXY`���cJm0�>}���#iv�f/殽��Z�\���_ɑ���wM�s�4�*��7���b�|{���8��O<eqV�G ��4=�&m�X��Le����P��XTbȬ�p�a�#}g9��l/��`���YS��"�`�.p�}�1�� a��H��8SjC�]������3Cc����ĜY
���#�N�kh'�s���C�EC`��ɿ���X��I껻���왵����vd�dn�n~�ty� ���7P��<vҮ�R�μ2|�B�ً[Kf���zА�4a�`>,�(�Gb�qV>[�Szs���Ȫ^+ =����=ۙ:y�>���Ȑ(����~�WS��~}1���
m�'ߥ2	��/�m<'�s�Z�N
�^?�^�sEJ�ܭ(��E5i7��o��?ȓ:�6��*�f�=��]�1�:.��% P<f�9���B�wL�6�����;д�w_k�U ��:��3��������M�H�BB�j&�5bû$����iM������((�Xڛ�H �փ�7��-��J�Do�3��A	?$w��o�*���ѓ��f&��Px��ϭ����T-���笅��(��}V�D��K*5��4�����h��{�=��� �z/�]�4�(ar��0�j	�X$���E�aeN�vR�����I@�=�<�fYi-Ĝ�J����Gl\ �4��H��E]�A��W��ݥ8���B9���17�<;���!?~6�������~BqPξ;�	qV� =��6�ȑ�3D��MmV�g�NT��ϱ��]P�0�u+ S/&�L�l�*�vݙ��c��ޅ`�ѷ&1"�[[7��t",_�-S4���z��������ޟ�z�zp����GhT9^��o���Q��j���ViCT�y��WN�>�t^��g�.5BnIgXY��k�?6��ݿ�^L��"q>)��P�����Wڠ�_���/Y���y�s*/4ps�T:�[o��-�l��=/�;5����yt\�Տ��,�u�Ǖ=<�Jyj�h��er�t3Q�V��t.�&]��S�+��H�9���Ӿ��B%V�j�]�����щf�Å����8�?N�B��!#�9���]ݱ�i��19ٶ&RQ�1(i�Ey�w�����39�T��@��(��W��P��֗Dg�Ɇ����炘쎡C	
�=x�V2DI��\(��5U�ᠼ[�C׉��\q�JE���D�E�r�!�mJ_"�=����^���R���[Ųyt6`]F�%*C�9�d��M�{��HIc�b5z�ĵ���F�U���zY5-��v�Z�����y{=���M	�u�Pe�������9�DFF����떊��*f%@k"E㱿>�K������z��tږ��MjN�����;�9J-����<E ��F��0C�%md��L�eM�Oΰ�lNN�F���c����E��z���gC˼�_�,%��A�` 	�m'6+ zS�O� ��|@ۙb�)ͦ�t�.䛥��>x��Z,�?J�=��@����u�F*�h߃/ǜvrls`�����{J�����Sv�IO�0})�S/�@d>j��|�\���db)g�RlF�r&{���\����'	���ǫ$� ��t�u�k�G�(=߶�K��e}�9_��`(��P�����iT�T�[�m1�����#)��O6ONq�><L8���x��:�����*�@6#��e4�E:鿱������b�-����|�f4��9������66�=�}8�ip�C�j��}~@v��^���-���-d�uA�`˚�yz㺞v��S&θ0�fL46^K���#KO�������� �`��mwy-]��B,�Ӝ'97!Շ��u_.).���$̭���c�Ɏ�r�C��*��+����	~�z����r{:㔄��!�"��ʜ}ItW�-w)�am]�9��fOz)�S���[����ʝQ�|�s̆�:�:	uzLAn�������WC8�kA��>�b��5��G&�3C~�~��ͩ�+ҥp�v �>��ۼ�5���K�y�	q9ơ�F)EF ��OZk4N�JZ�9�,Ls7U$���W  �er[ ��6��2�I>�z����a�~�������B����*�ˇ6��&��p�o{p/z��l�(��G�=9�bQ������`�yz�ɶ���	�]񼸤��n�E�߉�*/*��g���ʏIe�G�
��7&���>�k>&^~pY%e�U�\��E��w�3���ď��d�[-��]�{G1���ŅG@74U���B��ǧDx��8�Z��|��[�@�V��RDϚ����  ��n3�Y�����:`A�3TOBH���Q�OE~+]�P/���U.��P'3�؇8Yn*��ȪL5�l��>E�����_5c�V?�r�� {�e���̲�y��\m��*�*�a��$�ۉ �8}�	?#ԙB=�T�K��r&p4��ɠ��%�%�X�T��t5��%�w k�-�r��Y ��$̶�L�#q9�k��Q�6�����ڳ:�4�����̜}�gs������'|Bn������<�#���� �b���R��W�Qc����	a"ࡱ,L�o��'���cs��/�C^"v�C��D����0�������⛒�2�X��v�cz�ʑ�︣F|�����Oؾlvp@*go�ɝ��J�!1�)�*��$�X��,�S���� L5Ӏ0��������mΛc�����t84?��$��p~��U�T���x9����߾N�x�.�IA�B����<�oڙo��!o׉G)��rGs�J���Q(�YVO��E���y�Hb])=��9�p4����i��!���)n�-}�ިKԒ�N7Q��.e����	�a��酈�Q(>#U���U�؊V��w��?i�]�a�	S.�p���f.��U���⁗&��v�����~9Ӂc3Jl)�A�v�u���yjpW�v=g���v�E�,����ivYqY1��o)<��3�@x��������Z�
����Sd��Z1��M���؞a�iL9�}������#����չZ.b�ܔ:[&y<\�G�b�
���g�>�M� hz5�?�p��g�ݽ�8���k����I�0�/��\�ɍb�<Z����+6���A����.�����Z�{j����鞤�����j��K�K~^'����r�{��ۡ�N-W����U��4�v�?�}�%m�ڈ�9V7<_�OX}����m�՞.�<wI�CFfy��u���:���&�y��˨���
f��p�-�\�7��G/ӵ����7��,j��J6��g�#�pqb.�ͤ�	2Y��SPr��#NP�a>���_�*2[��#E�ǲz��1zQ
�7�j"��?���=�òw�y>$a�H�r��>����2c�X�X�HL忐e��^�d/�S�}tI�QÃ���p;�Dv�&���W�'���}Sk���+��J)�����4�0�Z���۴ ��]g��$���$����]�3S�<�Q��p��W>B]V��4�z�����H�;p��8�m\dV��LBL��Q��ekѷ��s����e2���Z8�Q�mX��;[wඥq��s�hN�$RH�eT%������,ۡ�fD�ܢ��ɘƵ8�]��r$f��W0�N+CG��0%��Eݼ+��M���������z/Xl���+]h�Hmd���p���(&)��=����[��^�,�5�a�:�Hi��ĕ����v�(��mv��6R���2���HU�鎘Q;�Zʗlf�1��)ؾ��D%�GB窺�.ܠבZ��6�լ���}V��2.Y�X���s`���@��{�ɖt�ykBbS��#x�d�!+px�O���E��F�n�֊���*��b�'jc�Ƿ�$��'����Q4
!}�?�3��[�q8W�g{Y��?0䋎�%Zko708�Ϲ��$x$���G���['��A)O�������4��?#3czB?�T�L��Y��������C ��{�?U���z��+֚pZѭ�y�-Ё��@I��u��)����m逃?̂��,��mu��	� ��k��e�	�(M�!�]j�*Y�fW$w�	� ���?jH��Go9do*,��`SBʶ��O�R�:)*̬n��qSEׯ����f �{�]d�X�	О���,���u7i�����L�ӛ�9�&o�"Y��~*�ѪU|��D �ƶ���;&||�,m�v�nb{F�D�2 �Y/�'y��:����i�c���o+�9��\���6#�����kq2y���$AS��؂��'�r�6ԣ8h���و�ls;��=U�n��!{�e��U��U���CwGwH��ЫvWfAm"qᱍ�v��ƾ��,�K���/�%S�j_x"���]<�[l+H�6����ʹִ[�xXK���[��w�{{�81;�=�j<�y��q�����'�vZ�̾�MAby��c=T�ra�I��t�ҩ��_C��)@u���'q�=G%9pI7���Ev�_�u��)�����G��\}�ҸWR ��ʖ��/.VԨ�`~�O��'��ĥ}��$eg^�{t��z�j�
4a��'��'��De�5��,�������Ԯ�22��~�kE�"�V�zG.�����P�f'GR-nđ����2#)��%�m6�bi�w��&�����b�A0��w	/��yyw��u -��t���a���ZK�����qm���ށNdb^����Ζ4F�v�Z�����?Ī�L��J EJ?��wM�i19�x`(H���=o�4[�� :i'8�Ki�z�#wV���%��\�L��<�&���_x��-�	U�oL���t��p�����-���V~��j��^d�u�=Luj��~6���	�҇M�u��m,�f5�'��a��HEû����tVZ��:��/#��Є�"P6=��˕�߄!ɗғM���_ԥ��&
J��Vؤ��m
'
��78S��V��G��6��8-�Wf�f����6h0���3nˏ�_/OJ�X�<dzp�kk�c�5]C�- � ߞ�,�)��A��K�f���i���d��<�2$���[8>ԧ<j"��ڕN$3gd:�4H1p�5:��#j=��;��=�G\9Im�p�z�j<��P��?����b�O4.�=)I������<�A��yS��;��WC��	�Xl�\�M�Ey��n�O��F!�zq]�MО᝕�w�2�ׄ���k��QO
�č��fj!�A�ym�e����$@�%���i����&�Z!��9̐��z#ҳ(Fz$�Z�s�p\rT�+�4Hߩcg8b��(�jwR����vԤqd���5[��}=wFr�"���5���_�E%ܟQ�I	h��H�>۲dE�Uy@��xwf�Y+a#,�xV�Qv-�ST��{Ƕ��т@b��I k�����3�&��4��Q��x�g�t�ZNL�((a�ƅ���BR�u�祆9�Z�)f���df1�|w�pd𣵙����t��{Y,>�B��s�ko��ӣ\���_>�?%��XsR��u�rt����]%����T���u�m4����i%cެ\r���Sեpױw�Vg�<�dIB��3b$Yҹ��p���l�\�7e�Q`f?�L��E-ЍQ�m��V"��-���ө��H$�=T��Naյ�-,��}�--<�6����w:�o�Ld"��D�H�������>f�MÌ�}j3Y����5��sCP����=�u���(K�P���3f%=�+ΓR�A�)�Y�熫�{.!�$�o�.HY�����?Ņ���Ր^;�!�p�����6w��%�g����L?q?�`�c�b��yV�����"�L���#�Cgz��n����]����Io`V{���3G�g*�%"��h��ny��O��g@q
�k�4-:�3u���K+HE4�}�(�~l~fr�4����@(�irHQؽ�G	[$۸r�ԋ�,�۳Z�q]P����0Rώޗ�)d6��{"�vn�m_�	>�X��p�HC�ʤ���[��.�f� ����13^���f�	G�N$�s��k���Qͮy?RT���.Ɏ���@���`���M�r
'-���m\��\w4ك��j�*;#�7���'��0��^���+��\�U��QG�	�N(fx_>y�Q��q�_<jt�����h��_�d��I��}R�'��'hI}��9��&5#s��T,���yb1���L�3�C�
�\�S�
�����ۇ�Jd�Km@����@b^�[��Tz�0T��y�|��4H#����[�`�_���-v����k��^��7�wb��>h�3,K��՝*\w�(���|L��LO��ip��v�c��U���Ҥ��ܦܔ��>h��8C�Vb��q�f\�
db��1�	�/�+F�^�;$#^��H�!�̩�*!��`��Za�]�u�S���	�:�Y��߸n<�T0�a���c�]�g����t ��˱��=�VYN�x}l�]��k�d��� ~ u��Ƥ�&���OS��nRi������>�WĠ��^����d#-P"�F*� ��ڶ�A��D^eq���҂=Gc�;m׍ e��-�'�w*����z,�O4�m��\����D��~6������m�%?~Ma�#��F �ZJ�2_�a�y5���x��$�����?�2Qj�[�W�FR"���X��/���D��#��8h�ب�O���m��z��U�%�/��V����#��t�Fu�c}�e�^�U���l:??2}�8r��G����0��4y�-{bj�U�2��F�Zk',�	f/4�q�H��G]P��h�6����7��0RB�Kʦ\���3x���بc{ƑB��6�;SN��]{"V5!���'є9&���EIff�u݁����2�.f�~�@�N�{}��a��9��0�����;l~����v3(�l!�]��we��c�����Қ��WGS!�c#��ҧ:��@��#|)|���J�5t�^pe=fGޯ2�F��������i�Y�^��D�o�.�."1~�HFJ�~\eH����>��m�R�5<?�k����7��Zx���2H�.�0G�3z����l~t��Y�?Θ��Ur*qD�o�ق�k&�}�81�aJM��0�pFt���e$л~��jp z�ͮ��K�=*�}Acn�p�8�99i��P�R
�T�P�{�f�Ek����.Ϟ���� ��3s����6S@�2�F���}��iȽ�_��ZI8z�C�%���y���o�B��w�쥯؟8y�|�=��s��(���[�����
4��I�g�eE��4L�6I��嚷QN�Ѐc�ص���rJ�.�z�7£К��#��=���t%�=�:��z���44��G�]�,}m>�W_�@-���K���ڹ�������*
~�W�J� ��(E|�2�pb/v��m���!�+�M�Rp�N�E��.�i���B��:�\��_�2Yu$4�Mf�=�:�s����4�^'M~��<��w�����9 T=B] ���JN5� 
�j �����W��iD����4���(2��U'����t��������_���|�v�(d��(�_@��ʭR��nS\�.XXZ6�O9e0�	����]TQb-~�3
l'f�f=�$á:W��B�E1�dDX? 8�Y��'&�o��4 ����k�Ո��Bt� :#��3�w3�Y_�zH+��ף� }+�6u.�g��l]��y�Y~L��_�:W�j�����H���M���?0�F7�����g>\�#�*��m��\��UME�\�C%��"�^ ǂ������Ɗ�x�G���� >_Hw��������N��_�$�&�i�eJ-*rL먡 Xemн�3h�X��u�m�F]yW�^��u"���ګ���l:���B��^n*��D��� ��gT�驅��U?���g�6CCl�� /k��7T�w'���o���Yj�2u=�^s��d2�t�!o ��۱5���fˋ�6cGh��E�)��~���cw��)� ���IH4����R9G���@���lD���4�h���\�ɑ����"��:t1D�O�	�$�������b}ѼS`��w(C��ao�lmK�8ށ�mB����%����y��&{�YR������Ɗ�?���c.d���]���"�ҚD�!=6�9����2q�Ԡ)���9�8���Cf;U26�]4����}	�Qz��<Gġ�Y�w�w*�M#,�r*]����=�*�H�n��`݌��(��'&I�wr��Z�rף�����m!�xsj� C�g~H��6SZi�Ǡ�I��&ldA��S�ay�b����S-�Yz��?,�|�N��ְi�o6�XaJ����B�UzZ~d�,����F'sY�����ڠ�'�ꖋ൯ mG�TLJ�w+mܯ�4� mr�/J�V���k�}���L}*����ա4�\�^g�۫�xy_�2A�bIqMhv0*����1�h}������=�4@4i^`����nDa P_ܑ*I&V�x
Ħ�o����E߇�v��9�sj������������T�P
�.l�m�zT�t$��yE���I�������g�c`N���_���"�$���;$�-a�}����_�W1\�jDV��C���r���4c����B.�X��I��[��j�Е89�"�t�,	�0���!o�J�w�2���i��k�IS��&Y4�y��r�+��ι�e������R�|��c ooc�lVț��Z`�&tj�dZz�6yV�*̡��P�K���Lӗ�4��9�\��92M)P�s�F�<��0��C�Y���{��q?d��w5�����������!3���k��T9�1$�R�TYǞ��Ü�(�؇����3���:4����k�jy�� �+l��k�r�ǧ�&N�q��XͼS��k�u�p�=Z��TGF`��m�-�a�!q��<��"Wic�d\�Ҙ�u�\��ӆ(��ȯ�ċ����u���3�1@��f�P>	S@ِV�h(yE�l�x�i��L/��rTO�e�,]�q#�YS
']�����l�L|��j���|_L����ȫ6��@0i��&'y.�|T[�����i-3�~�8�#�xǂ'w�
�;���%�q&�/��f:��,u�z���n�#��ǟ�Rn�Qﭓ"1;����v⤢VYFD�-�]^����B���jؼ��Y
�}��b�j�8%�:c�h�Y�4T��l��D�^�Q���s���mnc ]7,�acb��:D��~��o�ϑ{x{�{�l(2F&��h�����c��A0I-���v�j��4q�=�ґ�(��ȃ�t����6��`�������v��V?5Zl�����Q���CXՠ���Um��b'*S3�K��le4����șey�x%����߸u�������P��L�R����Φkt�?�80�Fm�N$�*;	�,��G�2�e{u4�c?5T�͛'MJw�Vjy�@���ƣ��5=��'5����Ws0�B�����!�(��A�yc�6W(�����Gx�W��Q�fz���tz�g��|"�=�{K�	�0��/�}<�p<>A3�H"+�J�f�asp��/�t�m�w�� ��^��$t�2���\ f��������K�е���ڢ*�{��_Cu-��>��{����ӵ��4�A
�+Ѵ��P�K<�<�G�ux
箉4|$?Mt	���V�o;�� ���W�-�ͶGЅv��SJ(��6s6LL�����i�+nc�
D�B �~C�@+������ͮ�d�۔�)�e� ��:��:NG��ԥl��,!4�\W�}�.=�����qKY��<I*i����饷��c_N8EI��+柕����H���	�L
�:��2��^>��S�_��yP�1����.�#Nrޙ+h ��W�{�m\Mo�'D��#��;�.'�v:����ɬ�m�[�
�u�U)�i~�d�+�It�(B�j�ذG��&KX��W�`ZE����Is[�Dȷ���7�jL�a	Jg�:�
=Qk�{!�v�"��WiNo��Oc�:�m�Q�����]eѫx�N����@����f粇�P��u�@-�|ӯf��]��X�*�X�hE�'v.Ƣ��p�q�	�'hy��4�%r�wH���bh�xo�YH'�b�#�-	��f��/)�S���2hZ�O�V�#*�)���VӢ��B����l��~8
��,����p��1���V��x��'�l�j��(b��^P�D��iFٟ:��E4�{ߎ&av�)i����G�g��
D�|.��l�a9b��l�J�yI@��zm&����	1I�̡�n����@le�%FzX|����S Q{ۃeV;�"����%��`u����Yd�������U�*�%zf���AM��:W� g�C��f2G��Epd޹����O�Q^��;KM(`���O�?��/����p�Ј;v1�t�I�]�"�Q���x��nfψt��X�//��+Sh�jmN+k7�3`������]��a���껋�?By��3]p��� ����a{�d�)ʑˠwT��9*�o�Ļ����J�9� ��o��(���C�صׁCd�(TM̐�<��p��%X��Ƿ��>��'	�߽*��S� Z��c|�ϐ���]osi��Ε�&�M*��K,�*�I];w��Ճ�f����a�������(o��Bt�5_~���bkJ�hP��G��!f��V������lK�4{=�ʾ(a2h�����`�K�i5���2s��gJ|��`۳�2��u��qN̕#L/Us_k�qS�2�Ԃ�᪸��n�u����`ǣ�ԎFt�{�$;b��CycPt�/l��q�^��%=�����l��a��\�K�����eh]5qtO�}{��ρ,M�.���qV7O�^����dWTd��x�"2���+��X{\y3 ơ����a��D���x��e@A�:Ǜ9�0+��	Q��U�XoڠђH�"��'\�:���;wu�+4ԣA��#>�q�5�A\�L��^��K���ݦ��@���	�i.>�$jG�ׄ�J��f�b�X<	t3t7�/p9re�I�� >���C̤آ6csǈV)�>�S���Yߠ���Ҧ~�v�=��e��]B6v��]jl~8�R	�P��g��9�$P��/M:�;���x��̈́�ò�����*{��XJ"�zbO��QR#+(����-����z*�,��u�	�����W�rpO�Ȣ֞E "�ղ�#��E�x/At�~��[�9C��HWO Y�{��g3i:ZaXD+�^�E
���'�4��<At���J;�ԤL]��/z��	�W����Y�^�,�#��G_�b6DE� {�q��\~U�V���) 	��][�A��AY�rTs�XPL%2�o�=ݣ�W���Pv�ҹG�ר9��jvE��]�/�]���u��XU�u���n��L��:�M��b�/��D�	������|����5�:���}��>����Z`�G3�|�k��e�d>���������.�T��R�|^TH�8' N�:Qg���<wA|<HR�ǋwj�~���A�^���=��x�!�ERI`��p/MV�"�OV-z�o�5�$:�-G��̓M��d�ES�2��8��=����PT���sM��6��g�M �)rc$��
w�7�!S��5''���<���)��z���4b��85b4�Ǥ�/ƾ�h���m.��x��~���u%�!Lsd�<�4�ƛ�6��fI���5t�)_�
���[H�tz��b�H��&�`�1�μI�u�.C���ٳ��1��T{�����ș��U��n�d�ޟ%�Q8H�L�� R�����F�S��i�˻����uP�7�3������",��|8T��:���0����+��$���.�)n��ݿ����B���w��Ͽ�5񺼞(�lY�ɉ����G�x��B�rz6�6�D^�،S�Wl�V		+�Nnd�ٛ�9w�đ�½yQ�s��	�5d����.qa�/�h�O<{P����U�)5"8*+�B��[s/z���O����7�ݍ��+X�)qWZڑ>����p�.3U�w��g_
��3��>,�u��^���g�O�3 ������.Tl���Gֿ�N�z�0��rx&���w�$0��9��*��{@�j��a�|�|���I��p\:b��="��߁J��b6��{3ғ�US����j/r1������q:��\�jF˰t=u�ɥνK���E�;7@�B�xeS{�ݞ0�V[+�?�͌	����G�?�S\���.�'���󭺌Qu��x�`�mw`'B��
���a|���$�zh:^���U�j�S<��}�� !%��;�7���R\�V)d����D�3�I��gA�別�N�� t�]8�)�.v0)��Cm�P�x�o/a�Z��w���*"�E���.lU?����b��SĈ#R��*��dׯ�����e��7�	���-����$G�-+����Z�6�.sO��~�v
<��u�ɹ�x�eK��z�
�;�a�,�/��.2��a6D�I����<��ydE���ZR��}8d���Ur�k-�=���X����v�*''�SWf� ����Tc0��p�x��+ӟJ�# ~���Z���R�9��Uߴ���`����G����$m��`��s�2�
j2�\�	9����ߝ�9o~�?��8�門����Q���n,��Y0�����CZ�^Z��YH�g�k��.��r%���C`�c��1�]��8�T�{�����zu#����C?�P3ؾ�N(���ce�f�٣�f�XaF*�7��
q��6�����
t�KP�|/8���ў+LT�o����O#ѭx�)W�|��Iw#�����nJtNo�4��Cҟ��R7�J�,G�5�V��͆����W�õ�
g�p���gFଷlF�&׃�Hr����T��ᙾ��}57�q��ъ�D�9B��'���ON���1k�2&x��������?�A�X+(��j�Έ��*�+ZL]���R9�B"��X���P����;�*[$\_mM%\�����Y��ʹ���]�9�0�.s9�^vp֐��+T ��0"��Z��k�>	~�+���x:���L^���D��`�>k���:�s�'Н�_��|aX�+"����^YBCE�E7��!طqo���e��IZ����L� �(��Y�7��v��_+�	K�^	!p`�P'��E6��A0�U���9ID�=��Z��9⎍�"Bp�5$b����=��<ŊYBLZRh�'�H{dq���*�W������!:b����y�bC���=4��.n�v-ms+����l�5{-�p|}�4N(azD��%�B�����Gg��<�fx:�
�˯Aj\��V�E'1K�Q�r�k,0to���A0�k��4�e�L��0@��l��3���N1Hpf�{eۚ�׀1fi3��z� >���$�Gv;�v{���ᢹ�q��c����s��bNm! ������Cܨ�$�ǝ�N�5������dl"�Mhx���a0Ȑ2�o!|���wN��v븖(Opb%�:g�~���
��ߵ�i��Col��'2fg��p��33�䟡��hab�UݒoO_/�C�k�/��� 7e�>�~�pw������}/]��?��U֑�b[m�<t�.�m�ԝ�v4-����Q���8Ud���{3ۙ��O��d���0{��pGtb�6�C�l_���s�+���S���@�V�A�xǲŘJgWRQE�&B�Y��l,ޞ��Z��	>�n��Q]
��i����c�L�:o1~Ѭ�Niu��Yep3��f #i��?��`�(hB��N�;܅rOTz��`]o���®4�x�g��~�j�O�𦖊Z��2�]X�g�҃�
�4����k��:"4j\K�L��v˄=��8����8�Q:��74.�kу{�~M�ʾ�%b�n|ff�X�!oIi֠�3������;�.Ȗ� E�/dc�:��	��y��h�p�w��5�^y=��eQ�l��^߁�
�_�& ��9�U��ʲ�:��z�e��[����i�b���9
�@9���rE��IY��5�2^��BR� f����C��^��,2��������� ��/�=�@:h��.��^��w#
s�_`#x�(�5s�#�E�k�CUk�fEq�p�ˇD�р �`�ӎ:�k�����]1���}�^���R@{u$%Up&>�cӪ�M�j�C�}��V Bw��a.R�)G��x)�I@������Q꧉s�p!��I��+����~
�+� &"�"d�!1:G&�e��S��3_	���=���X
¸@����&�n���@�=ڈ�X��o@�	\�k�Tn�`Mj-<{#��ެ� ���J;1W��0�*�Y��ո\4��h����{XjB��+xҡ��<�r	?�-��9���r����-��<n0�M�����$��3,x�2+�<�X1νe��$Y1��ʫ�N��Ӆe�䙒�B�/υS��Os�(�������y�<�6p�#ol̺b����T��` ȯ��T�4��7]L�D��g�s3 �s��Rq������;J����a���Äg�۔� *es~�J��犒��T~��Y��p �"rd�'��lO�E3��n�2�Q�(����q�R>�����Ɔ%^-zZ;���=��ߝAK�E���|œ�z<N��1�~� ��h~=��h�f�������h�S���K�s��(�Pj�����e����?m��s�g�L��!�n8��w3���,�o���M�}�'���R��cxtE���ܬ<|L�r�I�d�:��m~p"j y?�"4�Ƶ��\��->.,�=>ƃ������_rq"������79eG٥����ǉE��$-�m��I�yLX*A�!�������5v�9����4
ť��EVk��K��.�ho�v|�9;2�����Ўs=D ����U�e{)0�%�T��頣�48`�VzVgiC{e�!A.�Ul����.��Fn�'��ToN⅄?�aP��
�R&�T��l�ya��C�}���GkUӈ)a�!��үe�B����p��)�lQr�v���o#gbH�e�/�d3�͞���ʭ+&	TJ �#V+S<�.H�~�
��K%�\AZ��:4l�lFnl}�rªsD��X�bsŲ%9�<���>D�E?U5<�<u�UIE��̡�߰�]�d�^����@��M�d5���Lq�dWRE�҉ҁ�� L�X���/yk_-	�s�k��Z�vؼ��A7�1��l�gLJ��b�)�?�P�����f.�$�Ve2q%�N 9I�3Bi�F\��u����<]/q�,�^�p�����=�!U#����ʛ�]�x����\����U�ⱦ^���Ρ��	Q1���D��D���Nrh*x�f�n|Rwx�c�sdX�#@�(Փ+D*sl���Ӣ�xu���S3��*.��k$��m,]һ>����6�u�D��;�c�y#���g��Hc���!Qڍ�	�����=�#tb�uS���k�����L\�|\�ꋥ�E:8^l����q�(�E�P�'�;�ٖ#SO�O�J	�N�͓�U7�M>=�6�	���2i�~�{���%B+Pj?*)]���<����Σ�n�_���:z���R��8�K�]pvD�����4�f�\�Z��(���?��ؘ������������ݥj��SZ �w��4�S�O�x��:R���"�]�"L��o��@E��#T�=H��#[�?ʪ�7ڗ5\�V���M�w�j�uO�-���g�k�M��ClF�fܮ�9~�ӂ�N�kl��k���k�7]�t��B7=����д�Zl�V��m�7]��}NS������;c~B���V��a�t]�ۺ����Ȇ����Ӗ�ɗf��ߣ���׌�c|\�ϸ_9G|G4|T	����q9wA�P�+!�d[�o_GG��:�k��&��̃9(���]��1�.)�4����0^s*(j!��\l(��v�C��%3Bg+��/��Z�!��|ͭ6�龬Jz�̎�M�Q��&Qi�n����9m��&Z���f�kyf����1B=W�RQ�����Y
c�������8������T����`Ȋ�7���qytY���J��*]��G�9�9��d&'�e��|�Xp�G�G��"W��snkv�%�lWlo���~җ�W߰��4���$X\j�5!�����3�\�;0W �mb䮾-�><���l�l���ꨁ�O�����1l1�9�Ce.PRL�S�n襣�Fʽ�|V��ua+(mcG����4Y ���R<�7���5|F�.G�Ư��0�0�q���Y	�^�=��fa&?N��G=���T���rm�MWˀ�Ƀa=���D�;Ў�ߤ�k���1M��/�2�$�J�c�P�����D)o�	��Z�͔˱E3r���h6��B�S��籧�wy٩2	63��a�����2ik\y�+���Ӈ~ez����M��;;��Y�+��� ���K���q�~J*6��Z�@�s_m� ˣ
'�h|,�k>�Q������q,������n��ĭm}ٹ!*�c�E�4P��O���	�����$��7�g^.&���R���y�kδ�>�G�zp�Tל���Q:���>�IQ5F��ٵ�FG��.�_�XGo�Mt�9�U^��B�7`@�[�1F��oq�]+��Q�Jp��*�.< �������KSΏ�)��*��ʇoB�FTzd�[{B`:��@�@*qr��$-�R	����y1.����fY��yn7D֛�������{xNQ�@Axc$&+���J\E��1�@��L_!R>-�qZ�{��isl�=�z	9~�I�j��`dV���AD/��[My�E+$�JR���A~�P��.d��M���=g׹*��jMj�U����1�$B���r�cb��q�N�猫 }sH�*��X/�'y^e��=�.>�O߮/��A�k�0�WC�?ύ�8�������ϴzj?��~�o�z�͢��O����x���2��(QE8������NMv�n�XQ$�~B�����9�+��U�8&M��i{�I)o�7��7��j1���v���	�o2���%K�R�:��T������Ϡ�e8+�w��ϧ����-��<��Lq�P��a��.ETE���;}u���+�C{��ѝ$Ԑ�����p��(�?�����3��o}Wpnag��lS�3&f�t6ghM ��0��z*yvv<������Q##�k��]~4�ڠ-i����0�zsȕF�C.�i&�$�W7l�)����\#�/��o��3ya��i�W#%�b��CnP/�u
��D����R`n�o�I��ɻ� �Q6��m��<��Ju���dw�-��|99���@)Վ0���'-=����7���y�A�vZ���:�d��	9L�lE?�K�_�_�X�����V�4('��_�x���:����±��L!d���Y�5�O�{ ���9;���+�?#����B��"��s�]3Vx�Q�RZgSD���܅��b�U<D�j\&&	��R����ETU)��ᶿ�L9w���*p�i8v�Dt+��	�!���� �۞�n"ʠnC�I��.DU��m��%N����u��?A�
dy_VC� w�	|���i�����xǗ)��V3��ǰ7%���&��Ysz�iK�$3Γ�N�濢���d�5�zA�ޕ����|�Ucwx�Qe�$��8�
	Q���=��B����.�]�+�-�+��r?\H����ֈc�k�	����\�#h�Lb�5����f���ny���� 7M�-p���AG|���E5~��C ")��U��_�K�\:Sy�`��,ኃ}��9�B!dP�L���>u��t�Qd��y�!��ѳ�s�t��6w�&�!\;֍il� 9%� �/�2j?���וR�C��ACb��L׍ޞ����u�|ٷ�;�e��M�*ur�u�#��Fz-yVi�\3Y�Ѷ=���^t�8�����9i���Z�A470��.��O_��m�x�f�t���o��NgouMB}
Y����jP	��~������l�E�/�	��������"�of<)�W7d_�b�Tbz0��|bWy;Mh����Vfȱ[��pϪ7�w�j6�P�pH�ti��>
��2��fR9x`u�$�`C��B�̃eaS�N �T�ټ�^tv��u�9Ӏd��>�ܯ���:�#(ҝ ��/��0߸���Q��Q�'�4���:n'ڝT-�%��5��>������2jc�L�j\�%/'s��s-��"ŻU�E�1��J@@�ܪ����y�*0�����:g��JD�w@���$�"؊[Ѷ:zAq�ZH_�f�},ڧ��viy�S8�4�����+�����g�`�A��a��J�[��ص? �{"�	p#�*A�4�>�M�԰�T� *<֕׋_Rw�k+��(�\���UW_�b`�,��Dza^,dZ�[��1>|-˼G�,Q�/�XKs��r��]�r,�a-�݀���S �0<i�oZ��6K8y���'"	���l�����2��=cCtၥ�ҫU��şn��+�����3u�e7j��Ks���(�G�~`.3ڵ�K@��Yڙ��F���	hN�S)8��D��z`���
��`n��~m;�쥆��FO
"����;��:�_�,c�]��K�� ����Qb[fcN
��g�;hB�t�����'K�I����ok�ov89�f��C�h5'�����ڗ ���^�O,�i�OE�j��Q��Yf:�.%kʁ�Zߢ��a��������0�_��4�_����	k��(p�~�����!턏�=wg�tݧJ:#��b�,k���4�$#�z5�-����830ފ��P�q;4�Fq<7������f|���a��yb���ok��=�.��,j�M~bw�)D$��;I��y��|ƙD�hش2Ѣ���Ox������Pg�و���F�la>��F�M\��ҚYCw���
q��	2��p���w�o!>�K���D+��S��/�Zr�S���F�����~���*/�qR�8��&��)L��/e]G���n˖�#������ydr��_�1�� �b�q��(<��lh.}|5k/*�ML\"�D�0ť�!�g��Ac|�ˣ׳��"�����Y_�(6�����fg�
��s�/X_�Ү��S�VD	�~�<3�E�r;��m}F�Y�T�Ϳ�2�� ��~�������FUi����a>2#�Be2��4��'}���x�A{:�+/�R��A+ߍ���!�)<����ŧ�����Y��{�h�Up���3� e:���f��,��"�6�M��r�6514=b3�/;u��U[Z1_������6V�. ��c`�L�]kW���L%�2�"%^��y�-⫠�ّ�tB�`�a�]:n��6y��+�p��F�˭�re�E�.�\�%�/N¾�Z��&@ �I���boS�� �����j �С�J֦�&E������(��b!`i�cC�DVZ����DrJ62w	�G�s��r?{������\���8��C�5G�e@���BՊ�3q�U�v�+!S|�y�:�?�+� �� ��knG�p�w�)�!�c�j��6�e!3]�	�{�� ,��tC���i��17��uv�Tp����亮���إ�ؤA��TLg�A��3��вB5�sy60,Z���:�;ѿ�Hu�.�e΃�<��2o�=ݣw�����?��������x�Q��M�K����� �U��G`�����>M�F�Z�r�@k�{[=�~w�͂�8^V�X����C������(��tS�1m�L�(�)Kퟦqѥ�ZKj�yw��tx6b1�|,"ި]R��u����א�<F`���cD���/�Ջ=�¥#҄2�as)�uPg�+��7mh{S�����a���DD�m��D��v4�����Ŧ��#"
q��9�=�����j]��d#`�8�a��]�tK>U�K*|�r�lm���1�B�{}���9*ݝ�٫6��S�lrUK~��z;�]��V^ ];�Hp;�"�L����-���_�������$#�\4@��ћ"��Ū�ˤ%/��{d�� ��Y�˔�������a0aؐ"�mi5���誆�2)�z���E��(���)�ž�P�0���� ��>���{VP\W|0E2���@�=���[t��;x]��T������k�%�V|
��O��Z����X+��,�!_iO�A;:υs�[�uD7�2�H�RT��j��������Y��l
6�3�OS�\DJӻ�2�CL�jr���=�[A*�N��C�����얘z�!\S��CA{>��O�4�)�«��VE�Xk�
��gٰ��֛������S����3m楞 6�$[a�z�9�Ecģ(�p��\bVF��j	gj��[�M��e�*\�NA��]�����+��K�(��wW׫��H���HKy�����pi,[,�Vߪ��$����ZC殘��J"xg����/<��w�ф=��ukO)��ӛ�b�Y} ;[��F��v�@Ǐ�D��)�\_�X�v`������loע�D�J
H`�S�tzG�{���C���H}����%66V4���W>�@�R;\}��(��>Ptu�����A��M�΢r�~�|�JL�� ����Sl������n]ϐ��Ѝ�/�v�B^����|�W�I��~�#%�R!��'�ϪqR���)��A\�G�����꠸.9��&!�4S��餢kW ��|�'�j��=��LX\��<�6��^��p������� ���c������2���.�l	
�܁;ъ�1i�.�f(����Q��&4�s���ʶO�$qYST�r"��'���S��ÃЍ�S�R;�0��<6������9Bc9���=�b�-��O���p.�ha@����`K@�z�l6��~����Q'�κz��M��tp7��85�9Ģ�Q�a������)�]�?�?@�JS�(��V27�)C���¥+Ss�n�qtL����eb$WC��������C_p��ٺ�����U[V4�-	�9x���nAq�w�w^3V�I�[��ɰ��2�Ҡ�A@;��V��~����@���o���W*�
������E��1����>7)ZG:��\hG��Hי,�\�;���kY\	}8*���*#A�k�cʎ��h;�Jo�b�+�dG��11C��C�K]ޖ��,t`�~�% J��".�秫@)��������<��Ayו�V��@�UO����|4��L���)���E^Q\c�In��`�^�$�7|n���^āW
��t���%�9*�
b�gfFZ�*@!��q��E#۱��Zv�]�����O/��żM7���;���+?�;�E���������V��i2���ھ,E��l�F\�6w��2�LEp<�+�g��׾C�Qx�FV�fX���������$���f	�G�g1�y��Y�-���kU�ǩ�1�o�_�:�������B��'��k�\�ǻz��,�Q�;ː�2���ֻ=�q�VM�,u�o�v6�mw��S�	�T-.����.E��/�g{ԡ���[P��A�]i�dI�{k��J?1�۩���R�ǆC�5���NW3�L��H7Fc����]�Iu��48<�w{pI�_�%�b�B$k R���mK�墶0k�S�2ƅ�Y��� =�˒��B2�s;'�N��5d�~&����18郡F��/��s���1)�`cD��׳EL�	®��Hey�-x#2[��5[�x��l���:Jt���~AJ�z<F�@
B�V�u~�3j�� s]C�B���1��nX�-ͷ��7�t����'�l�
?�������Y\%�2SR#F��uI��'�*Yֽ#!guJ�j�L�e_A�\X$�_�&�) �����O[i����� cC�R�54�������g��1������0��XLۈ��b^�b��F��	�;/�DDp�
�m��[��[��o���
�H��7U��6�w�I;�hUU��]A0=蠚E�4�)�=��Y秜	sׁ^I��N��Ff2Ϳg��)�`f*N�_�L�1(��G��^m<�ǔ�����(��O<���R|�p�GHs�s/�!3���PTcf]��g��-��w����-���<�S_�wo�" d1j���v�!J�*@��ꢑ�3�kD8L�EL���h�*'�!H��9�!�+H"t�� ]����ÒF�����Sz�'�|!;���[�1��X��~�}��Q19/"�ܻ�)G���Tqps|� ?��#�A1�~��2쭢X7�]��](����3s��8O'�8��8|�{)����c��ls�+������k��TjNFr��N�[�B��q�w��]0o��n�am>���0�n!�j9����p�9�;��.!y^`2���������k���G!$��_Hb�v�#�L������#$pw���c�?�Ŀ��9�܀c�_v���l@j�zi�4�z�k��p���s��%j���B_��J7�������X�,�t�AtڔD�'l����[��)���?��%�fY7WI��p�#���=�	�B-
�`��g�v�B�����h�s�K����JL���<t����!�3�EnV	05����/nPa��Zڙ�C ��34}�h� ,�}Jj��#�#?4�Q~wHC@f�� ���5�dg�ȴ�i)#V���KqW�2�!
&2:7��H@1�fu��,Y��鈏�7k4,�b2ʧ����m�0�%�/G($3:N�Q/���I|�� �)q�oCf�.�h�
F��*�_I�g�x{{PH��1k6~4�X���e�$������_i������V�Aa�O�};�9I��L2˞�9��]�b����o�����%i'gLv�b�u�R�5�ܱؒ~�yGxb��A�2�͍}��}�.���D�w���n��\�2�%/EP�ڮ��:�3>�: yu����J	��[[�X���&zg�+E�]y7�j����ȧ�Ŀo>0�b}}���g��'�F�b���A��"Qj��f4��ou�,"�����r���։�b�Q�ck
^�W���,06bz<�H3��.�h�&7�:ǳ6�����p��>��!V�7ہS�&Y~�*�� ��lV�D�t&_���ޢ���&φM0G��Uc�)��Ҙ����Y:�����Boc魠���E�0�<?L�A��kj��6���E���ݨ��n�bՑzJ<��s|����v���`t�ǩ�P��n>zU�=-�y��&�i�/#H�Ҹin�^�:������4���iF���z� z!�./��#�p�+��w����T'Ү��$p�9j��h=�Ұp�Ua��#R�kO��{H�z9�E��uI�YJ���y�%�Ad^��~�.w�!b�1���4����������X�)}>�f:��ֲ��V�/�u�WN���= �QTt�>��YH��	�O�����W�]�w�m��J��c�;��X^sX`H�Ԅ��4�d���W�KH���ԩ$�K��{��e��N�wI�*�QBO7�֎�]]*������:�k-vOF�(�K��/����	�>������|���a���5�@�`�4�c�2�W��
��S4���0�N�􉋢�x@��>�&I�@�'JP��w�	�W���i�U�䣬G�=��s^n��O�5��Β��l���S�ɨ�l�@�#��l�3�~��q3�k�����cL���s3�jv@kk��������@����`�|��L��d�ʶv	��6��=����&)yu���Č	k�ʽ=@K���T����0l�+@R�,�c���H/V�2�xkn���2�1�t�N�`��Y�A�pB���}
l),~�2����B�l�R���̬{� ��F�����!\<��y��o t>A�ev�ȹ�#Ԥ���o:nH\�z2��q8_��:�Ҿņ�pz�Vu�ͽ�LR�t��V}�
����d�A���h���VB�%��i90%��$ ��-�"ջɰক��P<R7�3����d2���^�cA{骄�#)��3F��F�X����W�@��=�ЃX�V =�7����^��K��5N@��FG��<ɏ!�����?7�R�#5Z��ּ{�A�
7�J��A��^�q�%����D�(Ao��LjS|:�����	�6����n���e�uH�d�>��)�m�$���J���N�q��ֲ�~~�>޷���\�Az���E�����@y5��^��}c\Oa��YW^�}OY�:e)��)�ƺ��4k3D�H֩���]��38���Z�>��V���,U�Ůܑ
��=/BYI�����A`�UK�������-<��^��|N/Z���Ӄ�k�5J��"�EԵ<W��jDF7�7�:�F(�|=W�;�BЕ�Ҽu���T�6�ct�B\-?��Ab��[����6vB.��O��V���W�{�q,���\����D��ȴHOP�c�,�/E"z���1�3��7���4A���|�a����>C
w�C���A0-_�WE't��R���un�rKF��a�3��Rx!!P�B�֫@.-"�CՋr�8Sp�z�<y�|�i��8=����I��P�9	��W°�<8c� �%%<��4�x�
s`��Պ	� H6ze˽�����/�ǔ���J��_��~���4!�e�p
���'a՞7���=��^��[s���%����֩��BZ���^ˑWo/��Id���b�f���^�J�1�Ŏdr�نֺ=���(��H�����k��zs�"	(�0����3�_C��sJ!Nϵ� xe�W
M9u}eŎr�Y���H��K��Q*��N��r+���*J��-��� $�o�0�pՅ5u��.�WD��X�#��ub/����Ds��щ�c�`�[#4�����|�C����{e�E��(\{上��6LS&�z��H�	�Wԁ��C�f���ģ�z�-vKS�6K�P�Ǫ��KoS�B�X;<�g�.5|��H�,�`_�^m#�ͯE����N�,P��M�$�K��7�;��'b��|gW��\��m}f�(��u7�C�GJ��l����}�֋������%�������ϕm��t]t�AG��f�v�:2L,U��ήF`�%j�Pߔc6����e�[��U��!�eB���Wcz �b�D��,'Sƙ�
���H3���"��)߲	.��8��O�q��"&�fTN�W���`M�N��-X8�30�5�����̙&�6d���)��o�#Enl�� ���*��M/�����,���%χ������aµn3�U������'	�ꕩke:��_pd��)�Z���@�b.8���ѡ˂w��@,"+��{Y^R�m�Z���<��X��j�'�#
�s8��z��;Z4c~��~%bp��5[`�Z��9;��y�=�j�b�<��1�tn�/��A��+I`$e���թEjW~\�5��m*�M�0�|b۟?jnO�֣Z�3|���5�=�iN϶�Z}�oZ!���Q!�Q-/��܏���Y.�SF7%.D$���&r��=��������O+w�*}v�I��� &9��ܠ��:����6.3�l%�	�y�[<
6��Yaǡh n��'���x)�m��J��W��w"^�-O���e��f�r��O �OU�G�+h%h��Lo,�+��OS�j��m���dU�t��f躊�߬-a�ޞ"�|u;���n<MH��������(,�h�S�@1�<	�f�d*ר���d��ֹ��Kѡ��EO�����ҕ���� ��Ҍ�e��[)T����AuO�M$�~N�J���:茔�m4'hB���A>H7u=�b)���Y�<�$��l$�*H�X�`//��.�sW���Dc� ��YG���N	gO��P��������$y�="��nGݾ��;bA�c�S�����\G��G��.�e�W�q�/FuR`K� �̟������%Qd�h�*�R��S� 8�r]cMz��e��tL�\����OhS��~����.mO��&�c<��|�0.[�h����Cf�RM�|-k8�-��~�D/ȥZ��be�;����훥W��d�.s�?����L��Uh+��TeSfx�C�2�9_!�#\�k��.����*��z�."��i��^��1�����J 6l����!�,(��!)0o8�5$��������".���yI7)`�ș��,d�Η�X�p�� ��p< "f�L�i�e=bul�Q��a(k{ޖ/��<2��h�TM&�� �G}w�DlN7S<�ÿ2󎺘��������K��Y���� �S7�ض%�[U,6����	>B��OF9�܊�J��K�5^�r���?6�+���ZP����uݰ����������o��O�a!�;�P#Id��;�⫱�'���Ui5"�΍d?�|�S?�Ϧ"�,���Z0%����:�M�^4P"k��u#���]��O<�0�:���[b�W���0uLX������o��?C��Iփs�NC�!��xnƃ�V�'���}�ڞ��Uިo@E=A�!g
z#��K�4U��Lȇ�Fbbf);�7�L?DW�*�A���/ggm��λX��wV��BS2�Ħ�f+)wc��"}ʬ��FH��x���	��yr�If+�z�m.H[�˂���\g�D�)[u�d�D�����*;���'��]��Ժ���^�8�A��� 
�`
�`d"}����OZ�mߐ�(e]rq���^Q�<rp�����O7J���A�z�`"	�g����f��fv�>��OY��G��6�!�N��+&)��/�� ���1ǥ���
�	�'����Җ4��q�1,�i�v�R �nHU�_���r����,|��G�bf�ouTh���?G�[�Q�z����e������D��u��*�HO�ֽ�Ao�>J�Ȫ�FSٮ�+��=�K���?	�E��L��u��FB����~�0$�����L9��C�8ee+XEy�K�rq�a�O�*�����f��rۣ���0��y@
֠\�����l�5F�2 �L����
�!�V��_t�1׈c~����s��������|���>�.<I�9{��Eݭ�Su�EG'e���;���3K|ϩ��&d�A!<�>Z�x�O�����2T��(�tf�{-V��)EyKm�S�a�+K:X��?������ߓ����D~���$?0o�P>vK��?0sK��a}���j��ƹ�NS��\�$?��5V�|(W�%Inj��i�f��)@�n����'���\G�*����G��������m�*���zx8M����jh�|O	�79�s��\o�m�'x�B(_g�<֤��n�-��iޮ!ۿ�`A�r�~�
4��bAo}�9y<��߶7M���_.��iM_���l����v���NZ�l����eD�/E��Dƪ��A+��z}~֬_��r��zՍ�s��Q��4K��D���;��!T���'�@�
w��)�8��4[����O��n����~|ވ���K�9v��57��Шq1.g���8�1S��
58�߂�U�w����^��{�'���Sջ3i}
{FIU8m�@2}jc>�\u�<�������~P<YDd%D��?��+�^0o~��pJx?����5	|>� ��0��e�irq�8���|�n\�z<U;+���9X�T�U����m����.n�]h,[�2�x��t���i�H��`Ȣ�n��@��m}t"�JK�'�s\5�9*3=�����q����g��gc]���h�(���2�xB�B��PLy�ּ���;��T��ZnFk���L��b���b��ʒ��W�<r*�_*��0�{���B;z=GOJ�Sc������':��:Je��9�+���%���qu���:A�E���+���Y�{��������t�Y�'R�"��32տiRAE�Ч܀C����҄}������ ����!�ظjV�o7�e���W�΂���Ʒ�,��X�Z�u��^8����]a�6�k��kz
��<�s����
��M��}�х1"���,+$׷�2��a:��4��쿪j��H�E���D���$۹�C��BN��M�Y�5��-q�����*e+d�_���(�\��!D`2C�BQS	9����t~C��P{/b#��+o�{<-��ō��0��L
Z[�_�/���o(��9aX@���R?���¶»ya����'M��k��%ě�*ѶQе\
�Sgc;�%�:��TΎ�E)��X! d_�5��Ɨr[�j-ڔjo��׋uy���8�{8��������鷾$�94I>)�f��������0inB�Ŵ��ၔ�0r8�B�3�?�W��q`(	83�k�6.G@0�0D�w��^�&�w�#:��S�Z���<#A���=GAwc�`��W����d�x���qL����7ٞ��1%��t� Y�Z�>Y��j��+�1�=��2���0P��] I�BY2%�JB-z����nG�p1ζ�WjĨ�gw{�S��^����߷�_�Tm���/uF8i��<P�^�C >&!�x��e�ٞ^�2K��.�2~�@�{M�j���*��!a<ЗROץa�ƹ���F���Ӆڇg.�&��x�}+hM�/Z%\��~ �kH�����m�g��=2�E����7g��;�ÃK�N&�pN������M(r,>��c��fωL����濴I-��^`6ԭ�<SLߞLԇ�6m�fdf)B��W{�4m�SJ��tx���cP]/��e?ٱ�Y�>�6�Ts���E�߂�������\x��!�T�:U�O%[:��?�k��q���g��	�4]x���`��ߧ|�����{�#���~��Bzz��Z�Ѧ�0�4-o}�b�ɨ1E~�g�M�*����}i�i]D�ntk�ưF�0�����b �	�����&�]�$��}����;�0#�������?zB�>M�Ի�E5�6 ͷ��7�M-�{�]�r��a�_�2Ϋ'�֣���tڰ/cLg��LL��1����ʃ0��Ȁ%��Ͻ��I��CyK�J,z7&���U�G.�vO�:�G�vR32�@���SZi�wsBÏ�p��K��m���#l���NGC zt���$l�Elr%���[�����R�V�[a�ָ���m:�r��-��=�h.�=H�:�D������݇� R,�
�Z}�N�r�s��-��y�4̝��
,G�h&C��ˉ0�ޥ��׋�A�Īj��ߥl�&��y��Ϋ+���#S֎!U>�Q���\�Q`���[����L�,/qO��\r�)�gR?1��k��C�'��*s�"	�<ɘo=q�q%��@di[J�aG���B����D���\1���O��Ga��Vg����WU��R��S����%;�7R�#��r6A|��l�u�V.�|����M,�_�2��ye.å�LX�YW� ���_l�H3	���O�^羜ρo�[1��7_;b�fw=�Ќ�� ��q̨"T��j{���Rz�`[bl���X]c�Y�����c1�0�*��G$<��8�w���<F�Y�h�������.�\.��Ƞ�9{�d�9��e*a�V,�5����3u�İ��m� i�]��b�0�F��@�>Q@�>[��4�q̡n3��Wi%h�#�l�8�������mHP����o +�����ޫ	Tf��t�CqlooA��Az���Ni��j����e��f��ALO�x��lr�:��0{#m!��Vs�gl��V��F�|y�`���h�ls�*�L���f�����겥n��֜a�F5'-����\`�|�¡�/�|� -�0��F22�v��b?ۅ��E��e�V&�܍ٽ��.�ť.�<uJ�G�ٺ}��xG�=y�"�t�b�����4A��R�KZ���Ǡ�k]�@�#9(�
z�5�S��d*aI\R��(�7��`�rg0�\A4��w�'����&�־!�I��I�]���*:�P�9[���v�+z�P�+�ͷ�ҝ��3Y������`s�%���c��Ce����
��x"�Ę�!aple��������������rv�ZH�k���A�������w=Pa��%��
V��y��jr�pTQ)^�:����5�e΂)O+1J��Ȅ�#�tE��c5� ^m4r�Cޣ�7z�I��ň.V��{�n0	d�Уup��@��ʣ�ʯ����!E����ge�)9�C'�������?k\��kz�r	N�Y����c�F��v��=^�4Fm��<{�ة���Q�];ⱇ�" #�}HK�^���dNi�4�t��7��F�ty(,�i+��,�m����|�%	���.�Up��z�w-�-���/�h���[�f���.�UM�:��z���i�!�p5�K^a�Z����)
wυ �#�K	�}�1���sN	����xY�$Ř�( o� �B^A��. <V9��������,��^� �<,uU��x��>>!���3�Xd�c{�2��`�^A�Z=�P��ޗC�"���*I����ϩ�ߌ�w�*b���.�W�ZK��n�l�ػލ0bM�� R�M�l�4ˑ#gn�ʬ�30�ZE�f���,6u�ot�~W,e�y)�� }�:�&m~}U�H�R��Z迄�/��C:�+����L�§'j�����6%��N�d#��N�a��u�JCTV�|������x�Y"d!�[�Z�UA�_�t���m��#���_%�߰L�k��h}goW
�?�
R�W��ĎsC�� !
�4���2�ɜ�� ~�6��C�q��`�jP+���*��[��!v��,��}���X|��K���rD����8v�O��Q���%܂�g�a('vٲ��SZ薬�۱Z��M�Խ��#��)�(}��Kگ^��<=o+ �@^��T�k�c{�tἦ���L�QI��>�U��ܐ<�587�AQ�OP�����=Ib�YX����p���(͋_�����QwkƧ1m���k`�*�w�iҙ�X��&���2�b�B=��Ǖ.`�/p9��p .�H��*���g�S�
�ۦW��JV /vi
� ������x�n||,<)O�a��Z�˥�`+��ka��n������$Vx
'}?\?	qsi����ܙiҙ�*���q2R7��G�u�2�k�E�A=�Η����+���3�0ƨ��5_~O�7p
vDD.��/��H�����&�����I�&Q��J��Ӆ�@+�T��-�aJ��{>f�oL����H��_���ӓXH��{Y�2X�S V�%B'*
��� W"��@������A?�:wIb�_�pA �)>������<��-�a �.D��v�%*%�� ˴���V2.u&�?��K�C��F�Ǜ�@ N2�������|a0gK4�!��M����17lǧ����l���꙳(���u�2��5&*.�/�/���{���7�� m��`τ���O.O\�闪����~(E�#f�1�����ҕ��"��+�?��]����b1�fޓ=$�Z>$F���8:U��<��A��猪�s��,/��꿪���:�]UJ컵jҍ�S�Iy"���beFn�U3��,I^vW�Yౙe��p���ж.��r�W��S/���rt��[��.�����{=Hް��`t�j
|�J�\\U���N&���h[��ycH1��o��w���>��u�Y�)C�ws�ǧ�V��aX�b�^��G�uz�>)e#>N�W�W�����KzV6�/t��NF���Rc2��!��	�Mc���"������EH�n�lBS�P3�0\w$���CU�_��!x�`�%����M"WNp�Ŷ�1����&��X3縹}���EEƟ�<R�ZV��m��S�⹐�/�����W��<���X� u��KmY4�H��`��������rm���X'&�N(y�]�Wh���Y�¥�Sd�YǨ����`C}�2lsޏ�Bv��5�l�ڿ:����I2V��O��͞*Hr���I�:X^����-i6,�5 �1�sߒ.`I�'�T	�h��e��u˭%�Pۈ)��B��m?��ʞ�'�)xx���Vt~w����@T煏KR_�-���7ރ>��`��]�4JTY�bϰq��*jF����x�����`t�������	Ae	�I�� �yLtߝvB�d��N�r����Vp�G9J����u�Ejʎo&+������{pâ�2��r|�{L���e�bi2�,��.��e�t����r'�s����E�r��no|Ik�Z2��������F�o˔Fm)���g��B��Qʗ��]�/�
���g�#��|�,>�g�^���_
�n�d�7{A|u�3�*S�
���U\���P9њ'7��١�8�%[f� U<�������C8nQА�P�F@�!�ک�!�]�;��F���=`텑�3Wc$vه֠"�Yh,���bQ��c�31��}RT�S2갱�>����:�M�X�.#�3<b��9�ü�ZX��N�k�;��%��j�#f�w�R�x6�3]ߕ1�Qcp�K������ٵ>��7���{-B�w�7��n�y����T!~8��-����!\Q�ś�M���ѽW��Z�T��@�z}�.���x\�^.4*͵R����?at��C�n��<œ�����\cC��xG����Q��ށk3ȶ�9e��W� ��J�/ɈdT��� 55A��R��`�W�	g��3��#�5CM/\ �܃8���2��'t�n���D�=�3x6z7�/	_j��9�b\vg_b�����m^��ȸN�.��<>	�����#W�í�����O��	��t���v�����1Hom��*��4�Zo��LSO0�*�w���q/5�К��.�VbI|�hdҺ�:� R��L����Yf�:hlֵZ���s��̀=�e>�hm
�����!�P�-O�c=�S�v@KMSH�_[~��^^W{��sB��}S���n*�AR�3˺E��H�}e4SN���_�?�`vx���e��FD���6�%�`�ˎ�YR�%5�?���`W�Y�m���I[bE���r�&m��c���nvY�7�q��Y���\;Ͳ���\��Ю�&=�'�'rf7�*{�֙yl��t��d�ԏe12�B�����o]��~I��1=�����Ʌ��4�����Y��B�V0l�'����NJ*���M �m�H"d�vNlP;I�q)"�9�������fċ�.R%B���A����ҁ�ùRj4��{�����ɰ�5��L�܍�{������� vP-c�����ț�}+�H�Bߙ�pL�:" o]T�8(=D���Ώ�rwU=����i?��>$�\�Z�3�)�D�ҵhw�mWi�_���PÙ'�d�ЌT�3�:/H[=Z����K������"<���^z`�5�S����W��Û�.!y���ȴ�� ��*m���|�vV/n�?\h��g�k�D�K[��M�<�A�էώ���q�X;�T:<�B��x�.O�k�'Ǽm[�̴�6a�E�t8h]��^�r�^�lK'��$o�r��K\�MkU��O/�j��8շ���j���:0Έ�D������lP�`I�pz���я�O�ОW�5�9	�K2�v�B����18	��Z����� ��j䏖YwB2�H[�s���8�[�<��b��biG�Sn�v
��ņ�H1���Y���y,[VTj�驀�������6�1}�q��@G9u�\j�h�ع^���3����+�]yü�l󟮗�:�=��]<TX�?"������OR�!Z��Q�@BgS!�B^��㼼��#yfqfk5@�ƿl��+ۆ*�"cD�ـ(eB�չ�=d�5��l'��@��_�x��m�Vځ��qs�2��v�J.bF��M���-�.c��:�9�r�[Rf���i6�������EH�ĺ�y�7�U��ҧB8�ԧ�K�4�zCK�wI�E��r�������guup/�����~#��9T�F5��[�m8`�kS���$)�Ok�S�����L7�	+l]�Ƿ�5�v����*%s(rg��O؜Z���I�S����-M�޿(�OV��I��ݙ6����X�U�E�O���b��K��f}��m�W̦y����#>�1�X�!:��5�Z�hU��ۄV�Ρ��k%+��&�u ���vɧ�?ҊL�		���
�1�Ay�+�L�*!+�p�z-�La���`���(��gb8�~��� �|�}K ��-Xg5#L�z
���0z��c��ԓǶ�PQ��v5��3�i�lӲ����K�:v�C�6(i���@�33vj�7Rô�+k��\V��~=���:-�¥v|�)���i/��K��cC����ud�h�R6;���V��n/��z��=�Qh|�88�=]���L��piw*[�x۳l�@ej�O~���߂��8�mW��� *�'�L$`�*{�z;�i�������soQ�^3RbO	u�a�p����������� +��*_��4��]]��\Z��U:�E��A ���c	��T�����kh�����/B��6V��Ohj(����}����'��|�9e@.O^.��ZI�a�)������SĮ,��@��)�ZT�pm+��'2�'�3�M0���+z�Uԁgh�Ș�{s�|0�[W!$�YSh&y�<练�t�l���o�� ��J�QP��%�5�eG����S���t� M^�ʸk��W����������4��3�`�8Y���Q���`x����>����[xQ�φϪ��1����f�#<���o��gKW���7^5ɳk0%8�뾼���mn�&3z5 9m8�y�����z���ȭ~BY2,�l9�FB�;�Tˁ*��f�5~g�k�/qV,}��i΄Y�������3�T���[q�"�^���h�&"k"�x^����Ft���6V�;z'HY����N��!Z"Z
PT���w1_҅��#��M�Sf��QA��PpH=x1^�6)+�����?�Ẍ́)=�R`�p������0��c��%���58���1�z���Xf��n���@��[fC�.wa��J���9E��%ScqO��sb�VfF���[=�r�/���S��C��d5E�b�@�ˌz4u1h}��7���=�􁊫:��n!�7��	x�Т�&Dސ	�\��Y�C���I����'����
:Bv�J�Xڊ����>za�:��|>L�׮~�v�ABP^�ScMR{�[��n��y���#�|�h���T[�[M=֔t�-eUw?� H��|t���H���ڽl�LW96�@��+ËJ,�=^�ȤF�(	�b�;��lྦ�����S����3<�'�Z4�$r��Ym���OHl�>]����oԀA��N���o�E��nB|Y�Z���oa|���x�Y,بc���k>�IJ�u��������"�l��eSx�RI��e��V9C��^�g���8a6C(�T%���Ϲh��=DR�3�+������krҪK.2�:���\���"��VE�(��Xv��l�iᜤ�{�߈٘������I["�m���IMn!oʍ_ ނp��#螾g]z|}0���z�����bnݲS�E�B���*�x�w0%�����4,�/���_��J.�\��yB$���z�ܻ���h�J][X4�߻LK_W�v �Ӝ1qE����M��,f�2e�.��``���-�E�[q�N旪6��j-���A�\��?B8�	d0��pD0㋘]�%r�Zu��˅�_��ڮ����x�7Z�ڂ�v`��v�C{�;���
����t��ӝ����fvSѢ�3�˨�nG.���%Zg-j�.ԣ�bG~0ּ� ��C����U#:f/��C�����D���J�7_�T��ى[Xb�k�4���Elm;�/=����E�|g�#����crb;�GQ�ڔ]un�o�F g�рj��$��j(P�DD~)ø`�#�k�u]�$a�<+��y��NԾؗT�2;�!��XMP��/���G�����g:b�J�s�^�{%�H����D���o#���̔W��~:
-�Z1��S���ƻ�wG��m�A��8��ˌf�������r��:���]�d��G$p�L��L��+����͔zk,(aaH�6�z���y�5?�e��\�g�k/��C�n?��?H��!���54,1M��}?<:�%�3qr�I�I	�9�=���b(4'��
+[*6��>9/�Ѧ����,����q�c������7q�|
~֍�f�˥�04V�wٌ��VJ�CL�d�,�w�����X�?F�Ⱥ�%j
�y<�d�+�k�����F���*`���`�huF>�G�f �$/���� w���y8-N�D��I�>�0p�S�΂LFarx"��(�F�H��u��-ݵ� ˸�2*��0��iv���5W��_n������7C9 ���7;Wf�\F`z)��`�t|I�O��p�4������O^],��H�3�C4���̊(���k��` �J>��5�^�2)w�Sp����.��㣴?�*�di��:J�[������s��`q@�j��� <ć9�:;�%'*��bx� ��wX36׼��3��h`��N����s!��N}�c� ?�-���p������oN�<N6�XrY�)GY'��]2�A%�mY��E��p�]�,���q˩�@E�ig��1��R��a��e��b���z	
�>�mMg���x���(�H�3tfS�����*����&�h{�+tz��;M�⠖(&��Am�����N6��AwK�td�R�����[�i���ט�jJ[��ўjxP������"���tt()Uw_�k�P�+�n�o�/��ܩe	�W��^D6۪��$��k��pS�`m�.��.	�2OkBjt:�表��E���4A��֒�ejL��ۘ�1��o�C�"�oo=�K�����������٠�ڱ�ܪ�껎Q�p|�� �����q5��x��ag�,Xk�@�]�?����x};��]��Ҋb��z����.o'0L �,w�L�����:%}��a&kL�� ��e:���;<ڜC}��g�\�i�:�r�x�T���g����YCH����o�n*XuP,�t��FQ-+R�~��˹8�� �y7w�mݑ`�MYrnE�T�c�L��W�����^��,���S��� �c&,����8�H���c��3AƊ������-h>���,�U���CEj~�Y�T��v��]�����4v��/+���V��4]�����~�O��w&��@~�� �_��	Z���R�C�r=�I����)0��S��#�Զ[$���$��K7�ɻ 2封��Ϣ��D�,�_xK�5��X��?��|}^i*V�C|��iW$L�N5S��h��;��Kd���t	r����EWŌYp i	ͣTT�烘�S�y�5��g�4N���*P]'#�[A,�}��&u���W�N���?���G���Qw(���g��N��P����~�xn����h�����E ��X�P�� ,����c���°��9��ʾY�t|I�P�U��'<E���c��V�x�d囱��.��	eb7�N"�G>3�lۯj�'�b<�?	���=n��:�GdV����[��E����Cai�P"�#eY��h#t=��U�/��DE/�w7�h���JN\��=�*���y�)B�=����
ͷ7P0���Q��d�E�{0xӦx�x�X�7��|��`w�v����jbЏ5l��yB�{�b)ɡ*חc�ʹ�1�eW��K�_23