��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ諝@*���gh�F ߄/R�b4*�P�ˌ{s��.5�3�_5"�5NYA9Jw��rU�I���[[I���)�E�9�i E3h,����Z� P��3k9?$�����R�W`�O�y�S��H�@PM�5Fa���(�d��ӬqxE�H��u�]�;V��Q�hǻ�����2J�Z>L�N����Zi��t��=�� ������i9��?{T5��e������}o�'���������`)��'���9�w�!���&?"v�*/fR�7��
�]�^݆����Zϣ(�� �Ih�{@�'R��V�僃u��]�c��H����=�ʷ�8�ler���-w�|�
�]�B����o�p�n���U��B~�^j�^�~V?�8U|��5����"Sx���"H;�D�?��	Ooxv�O΄c�7|h��Uo���� ��Y�w8��!�*��
�\ �I��v �9��/�2X/Zѷ�ҷ��ݬ\�/�g������� rA�,v�y/���8�JO/n<
&S���L�m�j8ϵ��2�S+b��+�����X���`����n?�w�l��pJT�)�d
O&���&9�V�Z�3	�b�y�`��7�f��Q�`[����w�w f�W|Y� �������X~�S:�pܨ��oD�#���+v��#i�����S�=����I���k4V8H��{.F�}�Ǉ|=��� DS��8���>H��3�@�&��P3�~)A~d�9��)Kd��4H��w��c)����B1�2�5\�F��b�@κ�y�D��n�4ʹ8�03 ͭݛ}�[��ׂ���x��k���]�s�iK�x�1
��,6r��US;��H��Bu )�q�lUYtf���Sey��>���B�8�30Zl�7pWL<\�:�'���e�]!s��?��H�C�Da+J�M�"65��/�w�����/p�������ݲC��w1ӜuU���n|�aV�n�2˹��$�<�M�A:���hC�J7G5��H�Xp�l��zhK��ޕ�6������g/�+H���Jo����@)�Q�&z���s�&��&q�1Z1�ap�C���suU���ݾ�MFE��yY`�T2�rC���7�/{H~x���bY	x�Ta��%�<�K��_��n�� kX���;� �ẗ!ﳓ�uy�e!S�V�U<�(=P�8�>�!>c�J���X��t�d�Z�KMs�V����"���9�FO��s��	l�wg�ƄG�����+�W"�N �R<F��%��`1���Df_�����L:�b�mfS3��n�q!� �ū����Ύ�0�M�+%A��W�?F�;b���5�cpO~���jC|e{#�ۓF���7kQf0������]���a�Q�Yz��.���."Y4��Uoy��zQ����m�u��=2�$���*`��|89%�%&z�k$����f���i���T���~2g�t��wf���M�*f2��YmVŭ��E���i �� �+(��M�uE�x;(�&|b�N/锱B9+A�"��+���s"�0�x�P5�N�~�i�-�Y<�^�Yy9�Ax�����Tj��Ц�_���b���: &�T;P��j��6����֠$���fFh�F��ĄT��F2y��2��{��ㅩ��ϾٛQI��a�fV�F�{��m��-yqG�/��:L?#�Ȯ �*�Rxb,O�u��eIݟ?:K�����,r�vʧ:(儢�r�C
���<aY�C6��)�[,dd�
��4���IVgQi�9^�:���il���ڦ�8;$a�@��Y��� -�i���BǕ���=b����L���I�:N˹X�#�g��i�߁o��3珱;��@�O���˃\�o=��#%&h�k�J~���
ef����yG��~�12�O�Tuk35;��)B���;U�QV�k�W��\a�9�,ldVu�!��Aq��������6h�5u3�q�NG�X��i����2寨:Qكl(I���H1����1��D�w3(C+��)�,u÷s�킇|����*e���JQ>N�)�R;&P���
s�!�	�[c̰2 sz��0U+�U�����ob���;�CӰN��>�,I����깂c �ο����@�0������NX�gl�JU�w����TȂ���2?܂�C�q_�L�,����x�[��_Iv�}"N�}O(%��a�N��$�v���ԉ˟I���uhWj���EZ�K��,s����?7 "p��u�;�r�33Y��0,��PF�cM��s�cGM7�S��i����N�V��&��}�PE�u�#sJ�>0�+,x��Z�tZ��$�J�l ��l�x��$�}���ځ���a� �4�W�qvAy��N���Dy���#�}�8�+�ϵ��]�+��3�*/�Z��.�hD��>�@���)�]#�:�Jk�4�M�A��Sa�8z}�wG�f�>���'��=c�#[ (��^N�s#	d7�ј���@Z�m�h3��s�N�O*j*@s�{��WV���2 +ʈ�4�iHM�ܖ��aV��#�����j�9(�08P�D����+I �n������<F���w��>Z�^;.є���E�ۗB�_>HW�/��v$-���d	��[�w�1�Ж��7#�����)<j�TS	�4�%���t���WxO�DQ]u���X��;)��:�n�.��%����a)%ue�m[-��ìl�L^"_�Ip��yQ%���9�̸ӟ����k����T4��z�N�K1��S�]f�����.�/��E]X	������~%\�����|}��Y��l���=�_�:��;m�Ⱦ��U�h���$"^���H���~y�r�*���b�]��uǾ���� ���/w�'�>`}�6�!/:͛:>u�;����z�t�~MHD��n�LdP�vt����*��N5 ۊx�%���[P��l�>�)�iM��c�u�.0S�n4A���Һo7zW����n���^e��ՀIE��,�I�
�-�p5 ������Z�u  K0sE��(e�йTu��8�?��8ԣ��	N�j�B$�?�I�'[9���T6"q��EV�E �gzrϘڮ\�c{��=��9�"��	í?��U�d�X�tsx��A�(1�Ot�v���5ZI5��+7Ǔ����J�Z�KP��HK�W^��hZ<mN�e�����7Jc2s�_}"��ڡ��,DZݷș<6z��$��>ɾ5�bI�h���6[<H�"�&V:<������B
-f�Ul0//G�s*k�
��M����m�.�N��+g�����-��Bq�yT�u�X��Pxe6�	��8������I�[4�9rN�"Qx�:�� ��CD�v��|Ӝ 
��%ŘH��?��y�.����hh�gzi^���f���]���1�A�{��AdN"��D��>����#���$�q� v���Q��(aj����\y�m��*��{�@�oܒ>F�?׸��@�Sa���>�@���A!�*h��mX��v��U��~�x�Y�����U��̊j'k6��M�Iz8s3�;F���q節ye��:��d1DEt����}Ɖ�SW�������$h�����Xڬ=�9vl�� �Z ��a�J{Gz�>��A!M�q����R����=�q���m~��!~�߬G�5��Ɂs<�j�cK10
�����ʩV%۳�䈒� ��8��H���-Zx�~�-��u�<�o�b���Es��5o��?����>&!>�P�|�}��֖B�
�D^�kT�Z4��ɀ6�'z�{��B��|d]ZU�����y���f�����7O7�56i���WU�U�=0��wל�)H��P��I��,�D��a�<��
���v�1�0��6W@��6~c:x�+�vP�~\��*��A�?�-�r�_ �u���y���	��!_lp뱙;���_K{|�������R�k�8�u<[�,-���s�N�S����2��s����̅O{چ����}��i��H��T-�I�͞��=p�cf~Q*�f�H��u�^�N4E��s�3�Y�����4��WdAl�����[���ɇ�~@��b�)%y].4�*	�)`��wн�b��`��gC�u!��u�wޓ��Jk�4+���j}�C�̧s�ߐ�#�Nnpv��!��Rܻh���쏩�e�+�[�\"��\`)c|���w*�y�爫��8|�{	8*g [���%(�y�1�0���H�l�|Qi�V�w�|K�[��P%��;�w�EV��sk�`�)���mQ3�����wp'��kQaȤ�ב��%�`aS
��QV��ߗӨM�4R���t����-��F{��la�{N�e�f�Gn��AF�Q�$�j��P�N����m;T�hB��ɀ�2�I^�5qx�K��t.cĵ���rH	�B��J�	�J�>�Y�~٤\�� j�#R���$�*�������S����H�'
=�P.���ʮ�����1i��*�)�
_��b�^��%f�{n0��m��F&�pO��$�-��E(e�ܿg�����F�F�<%��$��EqfОGR�� M��=:<����<5�T�*s����ϓp�.ޠd_ɬ�ߔ @9�-��ƵS���1�9ߘ��u���	$��l��𢃾6%���1*d+�K�bG�Z�ڄ� ���hC��Q#�V�U��J^6�����:�^�:e5��8��A)��_��a���cx��@����ȣ�+�rK-�U�2���sW:�"'��2�x�M෋�e6�rP���(�>3݂�B���5z�k����fS�/)�ʠ�,�,D����F�4���#�;����~�xm�KWXN!Ʋ9���Թ�'d��Uf� �7�H��ܹ�X{h$t�[%7��J�����'���F��=��)���c+��Ix<������y�z4���N4�s�]{���L+��CBi�z�'��A����6Shw��o��#�C�w�=�VJq:R��x��TQ�ŁN��;�P��O=� ����5��J��P~�bu�DG�=��E���"K��8 `%
Pu�
��L��-k.{=y��8�Y�9٠�ARy���A���D�I@����i׷ә�%^!��u<��|��s[��6�cx9�
��/L��M/�&q�0i��+�GR���"0m�0-̎4X���8���CW.thbsD��k���g��/.$k턶�,���^�w�=�����x�F�i����"��%���:bM�}=_��S���
�j���up��Q�xG�5��Z��{��O�-x3u�۪�EVE���t�d��.����.̭EL�	AΑT*V=�����	�g�G�N�П�s�ݿ_�L�*LBY�UT�%OWD��x�.�Rq��� v�#�m�|��sÜ�+�����h���K���J]�G=r^��ήi�(�n2n��6�b�,t���I��N_$\��\g�1f_pד��֗ژ�}��
"'	yEPn��뢯霱 痑���Ku��$�k��<��4��׊!w��_B������F�y#�n�I=)�� x���8���ه���Eo�tWٞ��� {�AĳV �q�I �+���j��e��TL�PzY�'����M#��^Ʀ�"�Q�brm�P�_l���2bfu8D�`W"��
q��W�]�i��Mx/�4/MNn���=��C״Σ�NS��
7��/��#�4Z��I"�A{�~_v��Dz�[U������B��sМ�c��9gZ�&����{m�`�i�>H��.K���y�������K��['~ �d!:��q��8/ �������Z�L��t�ٙ���G��j<ol���̍D$��H*kx�N��7��F�'1S��h�48CŒf	(|&�>��4���Ę��`R�V��myW���gy�$�������ӭh6y���f�r;�_=�khu*�֡s��7�$�G�7r�P���K�뮾�~�6����<CdI��׬yR�]ӛ�N���I��ݵt��j2|wE�_�
����T�d�!x��� d���(�C&��Z2폇Ȑ��k�s����n#�*�)Y	�a(RIA�a|3����]#�xSP�3�2��Չj�^S�����11SrԦب�_��Ĥ����
��Q����/8�k,���3JZ�$�^eݛG���d���=w�A�PzG&��Gk�Ė4'Q�|�
�ȻA���@�����#�s�]�������oY�mTͱ�������!�la�ԧ{8��$�R�V�F��R�����N��"���������7Ϭ�R��M}�M�e�:Hc�����p�[�Je<�F���A��]8�(ֵ�L��4Bн�?�U�����
7e$��03�V���)��\䲭�/R��FSZEO��\�鸒-Y�ᬹr;�ykc��Ԁ��Ә���n/��8.&�s �:m��¯w�X6ß��eف�''2��'�a~���H�.e�kh���"
�9g����=��5`��6�%ֽ���ғ_�O��m���EQ�f�w�]��x�k#H���Q2h��5�����1�\����u�����S#+�kܴ��~<Z年�+�2b-���y�[�Yoz��xJ�K�_(�.�ZG�]�}�����	����Y��I�b�Ӂ�����R��3g��m�y�c��[3h����ӯ�( �t�Y��Qx���}|J�"U��� )*��>̩~���!�?�3u�t6�8ռK��-?���ţk*T5��t���m��献���dD�t�>���Y]e�iyJ���������$��%}hǎ��ԽC��	T6� ��ae_�`��p��e�O����TL��P0+����F�A�BH�|�e��h+(k0"� �3��n�\C^_����H���ר�@����|>���.�ڛo�"�Z�i�t^�@s��ӿM�=�t�V'���Ff�Q%|�`������R�!�q�6X)y�cM4M���� ��+�ķ��u�RE�%��Yd�7dm*z,�p��R}gP�f>��l����ǎ����:��h]1^��=��/�au6���8i��h���	Z�l� �r7��騪�ƾ��`c�E��sLt=2���0����a��
I�@�	9̗�]�
�bdP{��� CF���Zv��WJ��+v	>wk,��("۫၃09�ؐF����0dA���4��!@�#�����V�R�61��nb����dEm�K�^�6��Y��y��I����&���S2�mMw������p��w��
����֏�͗�^J�1)��"�Nr	�8�h �^$
{�}�H&s(�8)��`�>����Ǧ����+�n����p��my��qEh�1:����_^Ă�F�j8j�f:�A�ܡ}� �|��k� �Mz+/��%ZfۓUaY�M�,���G>���T�V�S�r���� ۘ����rJ�@�5GcKy,~��#�^��~>�WKn�L���'�pQ�A�dU�qr��v'X��=WKI�7�ؘ"��4?���!Q��P	6Rv��䍁�ہ�f�n���s��٠�0��=U-����bt���B,Ɏ�7Ye�"8��d�ܠ��-�k��7�O5�v�a#���r�o�pq�5�TdĩwHȃ��0S���O���VR>�睸���w�����_�m�3"�\`���Gb>�4��5v�ܝ&#=���	��d_����0rwl��jW7��?��dd�y�vf��!.���u�OɁ�o�)t,Yx�_*�4Y�� <�N�Kݰ�� V��-YmX	⪭ޫ-��3"<#�.,:�.NQ�o�BI���Jx����e*V/�>K����E�`��^9�UT�#��r�QC��a��DH��5��[�z3�%�kRW�T�r!W/m�N\��Z�0��:B1T�u-�����R��>�M��J����Fm}�Aݳ��=�Q�W�J�Ԣ%p}�yP��j�:,���0�
\M��{ܹ�WBF�iQ���hjN���,�H]��v�[=Ӹ�ۈ�a�L�?�I�'��O��+����gpO�H:�� L��T�;�n�=GV͞�'��d�I#]a-�W�%?Ly�B��n��f���K�(�?kd7����O�u�גb�G����w�����}�%x�p�p��j��E�:��ʧ���>5w���������@��=����/���N�G.u�b��������v�ݥ̐�֨L�f0���X��߼^W���~��dc"Q��:	�N���6���k�.��ZW�|��k�$��cm��ѡ~P���r������m�7�r���*xH8vk�n���	�|IE�)�֕!��\m�� ���1JY�O}���^��%yя�DEv4L��Т�}�;|*?��7/�����.0LN����|�U:���1�ɦ�ujo����3���f��	Z���x���R�A�S�o��FI*Җ�\���C6�{(�VE'\�k�߫.`��e`���9�F����b�8<��t�[�gD�o��e���k4`��;^��>�t��(�� >���sx2|��L���_����W���� �����1�����˙zJ�1��"6O��Afl4?��(W%��K�*��c/(p!eg�)d�[w��.�X�n����V��l0m9��pó4�hl�^;5[�U����eh�	q�����g.Y��u0_ZM��1�,(��2��^{���<I�ݔ�2����
}�[#l�KZ������`6�@z!�J�ϫO��K��R�/��6���2#��h�l�Ϡ���W����t�\F!�+�~o�}?���ߍ���Y�,}�f�!�o�=�Gg�E�tŔ{�L�qX����ʹ�LQ�vÀ	X
��°��CLO�YQA�"7Cӷ�yA�Iܩ^�� T�2�2�f�.Ǉ0�� S�.�,�\�[�7\s�ׅpz*�S �������BWN��:�;���Nx�Ғ{L ��^�t��~ъ�Y�v^��O���۪�tHA�-3��k�U,��H���IC0i%�*��ƞs5����y9�x��C�E.�!�|� �مf���N`8�cP�ǑP�`�f��Ϥ����Q�4�~,�9;��Z$�n'&N )��Erz雨��  �(���Eh�w�x�\!!X�� H��	�)�� ǅ�X��.R(�ۆ���rY��@i��yt�3�+ӥ_����	��%x��Wp|:�n���6.3�:r|[���{ڮ���g�-�~y.�g��}5�mp��V5��-�/�ꫀ�������F����N1V��J^�HH4��VD�02Rq�^|]7�J'2���%r�;(�q�c׏��pI�B�!��2�;aT����K�2���J<�xGNL��Xu��&zWE����V�R|��|޼_����4J�I�K��VF�6P����vSm)D|�^Y$���nH���1���j<�'A(-�3k��Y=b�Se1���-��k�Z�7��D���=$���%�����ǶN&CCVg�C���+�����I�ߞ�9�I���A���l��C��Iq�j7��T��eN���?m݆�A��16��$5�*�s�(L���;`=��P�6#�*5 �	��q����`�n�-zV�̛��e��\�����O�Iⷪ�0���:���0p�("���	� V���������z�;���C�b�
�tV�onF�<�����ۋw�WC�B`v�g��Q�8|x���B��oI�����[D����>�_�^:�υ��,��Ǭτ��j��O�� e����=� �)�Rl� �ubv�WP0����]kPR9'֎�?�et��;T��ֆ �����X�k\g�S��_���%�2��x[�P78f��Jښ��if�J6���>����/n^á%�y���)��{���+�3��5�o�]LD�ܓ5ܳ(��P�5ICS^��<x��n6I���'�m��gT2,j����M���[\�������%��bJ=���~_]���~�-��ώ��@�x��A�1o��cTt}:��$ܪ���	�(i���cnW�����ߪ��I'Cr�U ͉���i�a����e!W�d{�a&�5���S��������D}���<����/Hֳ����,����[��ȇ�}�:Z|�z�dj��Տ�Z� t��:S�3�9��%�j�s�� vF�z�vk��p�8��������-���3�r!7N�۝�{	��5�T��qo.��x�z2��2��k��H�#�>�I)�:"����~|F/@4'�,��7Kي�_��R�jt�ё��3#|}��.8u���� �}e�#�H*?�R��¨����c����Z0	�6\qY�O��h��@�fv��t���EB�>V�`6���&�ȼ��1�W�o+�p�4׌�D��=��y�nHGj<*q���ȍ��c���Ŏ���ք�!s?;�v�,�yp��3V�LS;/����<��#/ͩ�.^�Pi���}�l�͎��\'U���^D���0�0^��߳�!�}����t��U��a�l�P�ٳ�#�؜l�n���䩰�~�*g7�Z)��ˎ���؍i�#!�e-�@�P�Ctsr<��o���o���ޚй�d��׵�ٔ��\�;��5*�,pM�œt�6F�`XD�C���X�L;b|��ۊ�&e����j�4���<��G��{��)��I��t���vۺ��n7�p
��+�krp������}#)-�!r�@q���4���y�8,
�)��8���C3�`��Ε.;M��N��r��?L�Z�Q�I��|8�d�'HI��c�uE��
���e�4�����C��V��&��K*����?Bkj��Ń����H�:��MjVP���Z��-�cq�#�PU`E�R^߉ʹ��3 x#8�Ut(��D¡wn�P��5�fms��ku�~;�'؂A��+��!4_�"ƪm��I���4�n��g���}��Su3,���dАC��	�
�X��\P.����T����G����2�.��{��
�'��%�J0�UrfS�,^�r��"���� !ȵ��K��j�e��B