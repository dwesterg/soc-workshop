��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8¢�}E0�Ķ��V@�~y�x�1M.�=���}�g�.(���T��O�6��<(&{�;a��=Z�����h6}��w6,��F�="W�l�r�L�lCU�|�`�v����y�6�7�xV��^,��^y���љ.��\� �����Q�����1`���!Y'���m"�.�JBFxSW������e'H�յ�{���يB��y����)m�*�[��L�˜N��9�����Cͪ�)�.f:&�W�M�/��,��%R2��Ѩ��{=���W؇�>����>����E��C���B
,�+�VF4�=U�lw6О��A�c��< ��|�|=�������/�JeP�`�#��p�jY�0���9{�$���/��Ș�Q]�U\��߸�\������nP���X�:O3� o�2�_��jY�i-#N/��_.�%D�Ī�ɮ]<;�wfe���}�נAb�L�2��>�������T�� �9w]���X�P��E$x��|��~�u�Y��@#�oWQ189ʰD�(��r�]��4��{�}U�XN)��O��N���$�s������1�ý@�$]q)6O�!�!%��6�q���$~F��DVot	ZB��L�/)0bT)v��ʹ��m#G-q��?�����6�]h��H�pd/}�s3�5|F�*�jjQ.ΙyTr�^�g�2&t1��=ѽ�vF5�䫃]��`E�AU�D^A|�<�0����_�����L���Ԩ26_S�:a���k���u)�O]�Tl_(��p�B��1�V������Z\�4��0��EE%�Y��Z�sE�f#DՁ�Yz�D�|���_�Y+���=S�v���d��K}S%��1��x���Ӕ���=�^'�I�Gb���5i��[��>�)�a�"�ӪŨGUج��X��m�<ĉ58��M�2���{�	�d������_j�L��E�L5��؍xQ^ٿT?����$�7��/'���G��Gu��9}�����I�Xϓ�{'�pd�^I����W���L�v�j�����ʔ���ة����%S�lT�ύ
�{n��:�3�r�yk;ć%�\�5��7N�l2��{�=���z	���&oT�J� �P�;�s� :Z~�Y�a��`hӍv�xW|x�\�'��u�������߂[U�h
}HO����h4y�M����@(�;�T�~nhx*�eY��&x�o���bn��
�P�X�w8+OGO�;<�e�����O>��9Ăhc(�r��k6�u/�v�<���s�C)G�\�gݹl�r�?q�{��F7�[N�/�F� �k����aj�?d�_� `� ֘������3Atsv�50�a�{:	�_wt�r=�4X����0�'	/z�;m�e�W4��o4��hY��O\�(���R����ў*m�b���g����>tz02 ��}�wy�t� �~���	q�D:G���Pn���J����φܔ��}	i�4��d � c��.��f�UN�Ν�v��6�S�]w�8.�(C��(Eo�myQ4�Kb�
@V<��L#�X���c]�-Ţ�;<Cg8r�}hs�X+��5Iċ6$?(Mcv`s+�H]u}G�$����`´ߔDi��$W�!p�Th��oW��$F�b`d)-Ԡ��V��&{r{PG�TWt��/�M̤��q��vCPA���/ޖ&X&�j�I-�4QErZ�=%�p�fj�dmw������� 9j�����~�OW������:�t�*v|+��U˸�I�R1���(~l����;
��$JĠA�5�����t�K��X���*�pGzG�Z)y�H`��^h�*t5#�Qff���^���o'Z�>5��U	��s�������{m���-��D�]�n|E1��	�"�'��?���@h.=T����5��$��fJ`e���9N,S��@ͷIK�deL�����]|�Ūc�U�S�qJ�`�E�\�Z��t�Y�{9MA.�S��t�9��D7�"mDOO��0#a�Y7:�F�eg����sx��s.HMP���Z����O�¿W<� ��N�G�n�7j���5Z� �w�m�����=u��K^bE� ���o�Z�ܭE"�\����5g��E��;+U�p�H<Ax:jA�?�ն�+�d��(��Cp!���\��+��%|�af�8�����l�ÓKq������5�	���ضOYL���x>^��f�zQ�k!J�c��as����N3��A��ʒr}~Z������f¬�+'I�::4��m���3y�4�/Ǟ��KN3�,*rEu��=��s�9UO|��C�F/V�m��ΓZXf`'�w{�h�/Vzԭi�����Zbx����
��?�l�Q��N��V�z�_~<S}bj`��PL=��� ��c�	��7�45e����】���2I~Q���@$#���:Q��l�a�ۗ�6ъ\3f<Ću֮�Ք�4j��W%�A6��s����p�2Ʒ=��WF�Q�)ɖs��(�N�D�l_��h�rbq�u_�B��4���i�rR��Զ[����r���U�P�����E�����������HC��� �x���=L&H����3Y��|�!ț��	#cA�y�ir;x<t�Ow��R�>��jG<3
A��@���AN����%"��b��$���Q0Řpx�H�fM���bӣp�o|hs�Fa~g���;�FbE�EO�Qo�gH�]��7>>����8�@��c�&�`i*���^[i��a�}ZS�e�k�U?����ˁ����
Ly�Sܷ�d_,�qw�B������t�-�l'�e��M�q���WZvi��Lv쐁~���%Hf�QaX��_���л��P7<���AZ\B�v���^�G�(nlMr+�����r~:̜_O��c�u%�����Z�JsQ�K����B,	 ���ȹcE甆�C��Z���D^�5�2�W���"��s��
�F�P�G�%n ԫԗ�#��L�8V�]�����B�L��u���m܄v��/|�I�q��Z"��d�Ty��.sP���?�3<��s\�˅�"���.���(���TS�!�3RT����ٗ�],u����7fS3Z.u9f�.�i2,���2�����{�g�f#�ۭ@�'�=@�(����"Ǘd�� �F�F����FJ9���O�&��x|gO�e��� 3�}��0�}�[��B�_H#M3�{bcq5>7�� p��=�D��b�Z�	���_�4���]�n�9�y�vϮi:vN(sPxD��uE�gQ�����)���I�@7(Q8h���3�Ow7�y��)}R;
��C<������O^��tY��F��Yr�sg��1ol�Y�~ł>X�����߹7�KĻU:��]����'�21����<դ������_��Bq���ł���H�����P5U��v��Bw@��ؔ��ftH��%uKX�b��������}ᡵx{�gy�F��P��zV�p>���)���1s��e�X���?>�֡пV�D��L֢����@�:x�Mg�e�Iy3����T;�_�'�SC3�f(�i���)^f�o��=؝�Z�T4������d>�ڀ����1.,dAgg��&��d�?��(Pv�Y���L�r͖U:���ʒ嚝ށʈyKl~c�;H�sk؜~Y_�����aHm)�g�"x@Е��ǳj��N�Ja�o#a�El7��t��}����X�J׆�|�h"��I��V<c�b��2����=�vr%�V"��|������c���e�7+ҸX�fߣ�����ElN)�L�q��S ��B�;��Cw�m��W�<`�$�K��|�A`F�K���A�Uf&�8��}�p�$G?��D//Q|�L��#��Y��{t������F��sB:���Zy�ʝ,۔��"Z�Ne����2����-e3?��_�l_��[���8�r�v��L�,|�������@L=��i�sL�^D%� C;hb��V������Ga@��ʋt'����o���G��F��'�J/�F�G.�uYW�Z����~H�];�A"ǚ����0s�� ���R���d��)](ۭѦNS��i�e5��v_�%��
���>��Q�醬`mZ1U�����d�;dK�Э�BT�a� �n+KŜw���Is���V�p��.C���,R�_
ő�7��S�o$�c�f�<�ﶚ&��]��Sv�~�.�!i�P���WJu�a" �7��%!0k	q��I���*{ΐy{u��,�5�I��Y��{u��Wp�t�����fG��0�ڒ�/\d�V���"���@J�1 �=i�0����1��+8�>zv>�K~U�����,��5�����B�����`;,V>/��%W������m�����5Mu��ڶ���8Xax�`�ؔ�=%��9!��ܡf�2�Í�o+�����`fB1�9p��	�xe�m�ȳ����NI�Gr�?�#�Z���]��?a4�c�?�h��k��K(òOg�rg��~I":�#)�47f����S�����`���A��댧�b�;L=if[˶�bC>��]� ~�uJ�І�qW#r�<	Y]�DrnJ������!筓�%)el���s3��\����&Yw��*����
	�	�ryx��3pa�����A�ˠ=���1�K��U}��<H�~u��;N�H�
k���ʽ2�����ğ��!W�'�|.XA�s��~e3)y�3� ����uQaV������-�/�E�vo�j�@�u�T����7�S��.(Xh,sv⬲g���O"!�*��lB
D�i���5m�s^�+����r�]��&���o?qZ(f�o���zM��?y��� �w�i3!��<�A]������x&\�>g��J"t�ӵ3Hk�ީ�͘���l����W�x��S��w9f�#�ܦ	�'���Ii�Q�2�����f�q�h�Nt�ϔ��1'�5�(#��/萿s5DgU�x