��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQo�qlj�����1�̀ޚc��F�^6+��w��Nh@���S �(����V	�K���ܮ�w����f:�2׷~O�xH���>;d�N�،(���x=ޫƢ�����:e]bڣ���"��gHf~�:��e�����)���?}��I^���v�`?C�Bi�&� Oz����S���>=��Fx�]��h� F�x��6��88)�f��Y�����m��B�х��X�K������h���D×��#�O���5���1c��}���_?�ؑ)�n!l0[�lx��ieH���v��@ɣ�z8�,�ک� ��_��΁�I�����O-ԥD/A�΃\��Ԥ�u�*k���x�\;P�沏�mRE��p3�h�3�2�x����6���._]>u�� G�138���E{����$=��If�b�E��h3�)����r|Wy�h�ޕ�)5�T�}��I���j����㶯��"�c8�"w:Ʒz��Ыw@��?��+i�K��W�cq�v�����2���/%���F�A%UZK���S���!�|��햆QG��Б�+�rQ�*���8	BZ �sHt��ϩ �rB��c�#��4��Ǽ��r���T��2�#��}H�TU��h�g��6P���3%��V��f�:��GX�+[&U�"��2x�\1"���5��W�yG���J����c�����O2$=��٥{z�A/5G� C��_�ra���,���!z2�$%�o|$�$���[0�}�Ӵ\B�ʇ��~��i	õdb��A�[-E��S�v� ��n$���A���(~��Bz��=eFη�ۡ�5�K��C��i5�����N4{�B�[ᢜ/�?Zj�1�3,�]�PV�n�JoT�V�d���[/p���ē��n�7�*E4!�������( �!�v���J^��jݑ�(�F��k�b�<��eg�,�U��6�~c��[�]�=��4o��0~\�4�?�&��r�=�ݪ�E@^C{�	2" �L��B[�a���g�~d� �ݼx�p���NWok�5��TaW칆r���?�|e�w��da�U	Z�}2\]	��r�����;(�1e��94�h���19qHŗd��kt
x��!�m/O@#��h��=G��z35�5���Y�ͬgV7��d��M~agR�����l�RP�됬w��:�#�6+�7��F�1A��'�ҏS�D�f:�iG/�Ǩ�]����l�4F"�O�U��)�,F�����@�A����'���^�x��I��bǕ��R_)�uE1�ta��.lZZh'��S���-ބSE���9z�{�`�,��{���{���J��H���A*[op����8=�1����l$�G Eo��g+Yc'��.��u+�ٽ��f�X�t�#���(�Z3{K��P��$m���j��_��ϗ�h�f5�Lw�����n�!��zY�A�s�m�I:C�tr��k�	���D����i2�=��0A�|`C��7i��&f�m�~�@'3&i���x6U�5�-���T���8I�@��0�E
o�*�ט��,�a�O؊�"~! �g��t�~�SA$���W6�E���?�)�?�+����S�Z*,28�t���Qׁ6
q���2���	�L��7m�2<uq{Q@����8����Q�J��jl�$zuc�(��A �}�m��t�%�j��h �^Bxn�h��9�P䗏6�/��g�MA��} �XO��oIŽ9�H��������Ͷ^����6QE��r	d�I-�D/���E��n�^�p��4�r����@�:"���� ��g��_"�����,}���*��DD\�}0��-�s�|'����=�'/�|�4���xM;�����t�d/�w����X���k5��_���<!�� ���1�V�N'��˨�m`����Ti�m8�^-�y�n��5�G�:?���$�����EyȌ�b��?o����*\���D}�ns .�T����Xb�霤��8�N^]��~8�G'z���eVi����)�����r��5�K�>�`��W_����o!P�,Ic	~�"BE��S�kj1��^菴f:�RT��b���C[I�j�W
j�4��[����9r�����2�[�ÿ3[T`)mpm(�����R�R��NC���]ڭ��b����FKq���72��n���>�RpUcǁt��♃�>;<��p]�);@ȠY-�'||B6���_û�����/(�@DR?���/�|�/Q�G�O��k`]��l��\���5	DLA���Fɦ>u�����