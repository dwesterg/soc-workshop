��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd_���}���dlX$gx `ڒ��Pi��×4DY��\P���1B�\{@���X���]ia�72Ι��k'���z��K�o}r*r{��1bKB� �>F_h!ժ"�V����C�H����3��t����V�~-����35��^=��J�����Փwح�^��I8⊐�&�Q��/4N��1�i� ���$�f�:��ۈNY�44]`m{��������+�.R9,M�S�]�k��k 7��=e��~��jd�l�B&���d9��Y�C�rB0���`�4|=���@φV�;%�:(����<,L�Nw�Y�c�P��6���~��{� 2�UxWjt�2Zg��j:�a(���u����)�lΘfۼ����#Ȇ�U���H�<���;��� SР�iV����$C�v�!/T�RC��8�jyЈ�?���.�������ѫ)3�W���2^ǅ�J��c��!i���*N��
Q���}�4�4=������������ʍ�n:`~����A���Bӂ@�ҠA-f�Ԃ�v��rD\��֋U����SN���������]QO��2uv<���U��uZaNgo�l0�]=�b�\���N�����>��H�����խ�G��
�j@K�gʙ�������Z�}'���iw���%�	g�G�,\�jA���	�k��X���5]T�*�"eja��4K���d�raZ
��n�!�<
��gm�|r_�ߛl�������j֐=I�t��];��sx���1S7i8���|��IW��[,�>8&	x�䋕|������`��J���-���<���0�_9�G��w�����sEq'1O��5��R$�p�O�㍼�]��1�Xu�y_6��
�~���o�l��J�hhr���}�wD���O#p�lyw���~ڪ~��L�aJ$Q$��Y|�޼�#����K�~���ZÝ^by�����S;Z��M'�R��buz�C�O6N��S8��=8!1͙��^n����nBs�ֶ���P�(��oNRჼ_���y�n�/�gl}�ʬC좹�=պ76W�%���1��D&�x�w�؛/ꦙ��^E	<������Ӆn����o3c��O	j<H�a@6�^�\B$��l�X��A��Bm�{$B��*ȵ�7cw]�)U,�1�=��,9����,&��]P�cj�,�k;u���yp�Ҳ��q�pQR����.�z:r�.������y[���i�C��ۊ�����RH	��TiI���8�µ�\���WS�p�ν<�(��F�Ψ����#M�h90}q�"��ā[Zи��9B��Ap��8Lvc����3�e,��m�P�����	o���w���]/tF;���]�h4����T�h-��p�p���'�b���u|[P���K�X��9*V��0;Tm���I��B��]<���I[x�PY�9c1�bي38G�"���v�NÒ\"Gny���u߇����|pT�`�m��G�"Rz�Z S�%��;U?�.�vA6ۢ�9��k�L7K�`%/��#j��Vl�?��n�a+�Xe�g�BbP��|t��h78������|y�6�|7�+��\4�N��ܣzI��0���H��k���\��[�+z�%Yo�%(U���"�d97���. ��>wf�-]ͷ������]�<�LEZ��qWO��>	iZ��cFGܷ
.�����%�l���bj����G�����$�9��<�迨��
̄�½|F���V�S�����-�,[�J�ˀs�Jɰa��>�>�2y3e�JY�3��S�'���8�k�@ˣ^��n�£z�����.|P/�쫶�	�=��uv
~s}c"��F��c@)m�6*M0'�M��l�7CN�ȽN7�P���N�BWD7�Y�;ؒpYӍ�o�n�+]��	�;���RF��]|J+}�d,���e�`��P[Q���8�)2��I���-���a0̑h\�m�N:A.�Ηt�����l��y�ƙ�+z�b⾯�a(=>$2w����S�Qm��_dҧ�q-�܅�R��iWY�6�|�mN�=z�k��E�_{��S��L�|���+��X|������P7���/	�����b�b g}��&" q���I�Sl����� �p�� ��9�!Ni��w��'S��>FM�u"$`�]����(�Nt��B����Ȼo�G�3���t���#�3��~B�����>��U.�*C����EW:�f���|5���H��1����/�*�F��X��C���Swe}���`J$3o�[^���O��Z�+,��Nj���� ��:VVV�����h�e$�F��&P@��)?��-bw'�a�N7�!nC���\��O`"ȃ%;V��S������y�+����N2ϖ����/]⭳���D~Ywᠵ5��%3D��Ҕ�{�ן��F6�����y�5K���y6����"�v���0�6��dm*��
�Y4�~��}������x���T�ڔL0=,a@ �y=�c�y��;V����]L��uʉ��x,ƅ3���W��	���+H�
�̤�_��'�q�Eg�w�|�9�Qf�=�'V����M,$�zX]�	���*Rd6��*�!{%̬k�������Mp�<bec�p�3!	��1[@�Q�M����Y�Q>-��Wt�mİh��3�ԴBq��<6�M�lƒ�a'�аG��it�U�z�=SD�B���Z�� ��[.�DZ?Yj�� �l��'8�\9J�R��|+	���|���j��y��dξ2���c��?=�rAd���87�S�'��U��s�lUN0z(�kD�hao$���b�5��/�r�h-���a���Ԓ7&�R�Շ�\���U���+��FF�A4�	MS��6�Y�'��G����x���q��}��x^��&j��Mj�4Ni���h�`S֠h��!���fS��?$�Ab��%dE����{R!n����i�r5�2��Yu�΃�U��U!�,\c�,�W�m�v���F�H<c\s^r��~���&��H-JX#�ӷ�����C�J��(b����q��T����c5]z�K�1:��B����U�U�B��6�쮚�M�kΆ/!���W�0�/���h��&��`�9��V���I�R��J�h�Y�o`" &2s�����^�k���ǽvUo?���q�z
u�����Ծ�� -gD� "��v�:	������=�\2�3Iܚ՞�E�C䘹���QqiS~ş$N�,�Lg���d�x�."���=-��4��Z�3H%�zl'/�J,�;��m2�=�u����2�Tj���z܁���BdZ��oh^G��m܂��.W�>Hxp�۷	�b�P�픹ÆH
pݏ�^�8]�^��2�1��i%y��ۼ^N"7�'\�Ϙ�=�
8E���3��{b-䎭T �����j��I�r�{���(�;� AC�<С>����!�;1{�4^�uhD}����2���x�h�t��E��.�~�����AS�GՕ�j<H�hQ0PV*��\��e����Ǹ��ezLH�q��6�i���~��/�σlaӚ<1���<ڗ*�.��k7�@�}���Mo�?q��ǫ�h��b��� .����Y�&����b��Μ�i��2�!yR��d\�q�&>xŢ+ѐ���-j8�(����w	���5��FS�1���N�r��Ǚ>~;��@��H�s`�N/���ϼA�����nU �J'f��Z�k�j�.PF�?�|�3�N��(V]s�����a�Z����>���qRa�`e�I�,y�SH�أ�ɚ�@��}t�$oulJ+(�#']���>]O|���|�ںN7�pq㓥Ǐ0␳UDX���k������z]E�ݛ�v������!�'B����5�)���+:��r�6����ӕ�zZ���R�m�F5״N�����Ւ���~F��ƥ:��p���zK1\��A[ ���c�Ke�Y=]�����WQ�n
5/\k�K�~�J۵�p��f+?��jT���Y�=kR�'��D@���U�`9���|�݊q�������ԩ�U�%�,AY^q��c3R��*�$D�e��_�1�B�Sp˱�fr�,�����3�.��܁�Y�r�<���X�\j^*v��(�Y�����}�!ᛨtNz,2�