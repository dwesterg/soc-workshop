��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M��i~�������8NQ��b�.�sӭ���厸��g�y�aU�'��4�a�(��@��џm'>��/�aRQz݃��0�g���~Ǩ@K���^
x�4�W0��1��*����v^��|��v�#(�0s0B;�w�h\tܾ�7��hPz;�~m7���+$&��#�>7���VH�6��/~�l�I�4��.���ߴڝ!��,�$\�v-�6���Ud(����z}��l��G3W���v,U��l����x�k`S���"���H$ȩb��M����q,_y��C� J\�UoB�.r�_��8P��$kv��a��[�˧�ߚz����_�ްr�(�L�޻��6�;L�HSHՆ��F�VI�O� � ��%uO��1B�� ����{ҥq�L��Sk=HaT�:_\�����]CM�#;�H����:L�2�Q|<��,2�\��e�1��eh��Vo1��\�x��m"YH�2�᛼��B�����J��Q�������.COV}����ҝ��N1��	��a���*ZWUWѧ��<�tU ��3N>����'ϣ�k0C��U���>���D3�B*����tdBJ��TyZ���T�������{����Ӂ ����"	v�Mm���"�q�2�� ����-UHSL��s9V��d��5� S�����Se��x�-�g�?FP�zpD������{ ��ŧ��¤PG�T��ּt4B��r�lK�M��S|��"��[};>	C�<�Ѓ�Ĵ�G�m��/{~��wfX�H����M@|> �R�@K��ae��r[�@�T�����=C�ɔ�/���i8���D��oF ��Ak�<���q��<rx����^�;O���y�� �*f���
˕j���צ$*�h��z������K��%E������&���i���l٣n	yW��6��A�U���6C�$��aiK�|�㏦�	��}u���ȫ�a��9��7�e
�����W*�"�.)y����a�g1jƥ���������u�������/+S�,M\XuZ��g��.To'zH��4�t���
1�SH vNVO�0gB���Yum1C.*z����E�l(��B2ݖE�Nfw��7r���G`���:�=[��~>��)��\38���L\U��mғF��JF1�ֈ��}���������Ug��@ �Y����"Ȭ1y&gO|�*�N�_��oF���Uع�Y;���V`�)��u�?W�U�
��f�"��B
��
#JlN� �yb�I�v=�~ol������;��K�m���26@ �N���9�՜�������ч�E�����8^���ߏ��x����䂯z��ɉT��	��Y����/ƫ�*^�� �d���ݍ�`f�@��*�>ʰP�@�� �hN�@��ډ�.��D�%`���#iVϯ}����A�;TE�qu~Ս_�k+�,]��C�_J�D���_�_b'R�Ο���Z�lGD�������J`r	��3�"�҄�&�n��&xSŘo{�b�_u�f/.N��J1�\���Ϧ8󨕬;}�m�lZlh�ؙ7TUM�E,�-qv�Y5��,�A7���<� ��H�"r�N���@�יNuTw�^��i
�;�$�pإS���d������n�"՟�oOx�� D�yH{��/*���ZW�k�Ÿ�[C��?m���Vr��T�x��Pa�O���$��9����'�׍��iQ6L�R��_�/Vg�#ٝ�=��<��3�Et���Q�IU!���j:�{�E1�&ٶ
,��'IO�2a��!�D�D�2��N��s�����㸴��3d/K�q���/Ŧ��^@*̢?��j����N�.փQ��T���m��Mm᣶�D(�E�������<c5�eJPQ��Լ�lhs�=�E���׳��U��F/bu
<bcb͹�g�cI�g#�p��I>�i�8�dkTE��TȲj��6�Gi�pGb���r�zf��W���=nAݴ�D(`�/�A�� h�'\�&4]�����Z�"-]j�����\�c����֭솻h��Ñ�N�_m�|�uWO�V��O��
*\�/�#����K�t�ܞ