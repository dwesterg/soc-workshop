��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0w�N���Z�@���8�z�W�꒪Y\�X��m1�9e�\�YOb���h�6���LY�[�^���q@��5�a�r|�81� 
�$g.���sێ�+��w<Q!z$�?Lđ�(�:��� n|-ú�E�YA)�'�n�\���K](��6�K��	��Wf�E>]���k�d�!2�]�{���։gF~�+����O`�������� �����<��)I�Ȟ�X���a97��h�#�t�ݿ��~by�4�@o�va�������v&�5�C�T�F�ԅFհ��Z���M�'���Ǥ��|Fž�+�(L�����u7�8x���q�{l �� �L�k�0��a>tF�n�Xmd�����Ƈ�fQZ���OM+GT���]��K �U�pp�R~\���U�-e�|�+�gMƙ�/��D=N�^^��H�:]�곾���[���n�'|���M��L�.��?���6��!:�4k��ԎJ�_0<j��^��?�H�Jv@f��B��6��*eх֝�u-|e�HXz��B����crU������%8�h�����D_e�Xz\o���</�Gg�-#`��Y�C##YJ��s&���8�u4Ukwo̦-��h�4,pIc�b�,}�.��d����ɢ�^�E���W¨௾Y�I��]�jS5�I�}g�+�����/s9���P�ض���X6B �L���ՙ�^K2h����QǺ"��]%��"�*��N��<�2�&~t�8��PdI�
H��|��7��Bw�����^�n�w�c�SW���:d�z��m��x�Y�O(����:���� �͹����b���f?k7&xx�KZc�� ���'��}��
�>֙*��p$~`66�+}�{�j���'�H�2�#�܀$vF�y��H��x�'G
3�#*��/AW���T�<��/�|_��ԩ��9h�3m�,���s'@�e�v:[+;�ԍ��K�{�{$�&���v���Ld�Y��81E֊|~J'uv���VQ��]]\w��,�Wm��������&���4֬�K���*�t��)�37��V;���68ɿ��(�t�(RB�V�Q� �Nؿ���C>8���D��hmJ�ݷ�CA�VnCV��9��^��n�9^�E���W��	�y�S��{�S���J⠺(.1�BH�H�hZ݅��Y?������^�L�pni炘���O��2�B�l���i�6��`Ƿ)�YG�O��M��a�e]E���5��&`|���~r~��Nz'�S"����\������1�)�+���8p����[L5��E�@s��/Z T+��A�矠� �P�Iȏ ��.�<��K��@C`���9t˧���4޹imG|���JA�!y�K�EM�(�2�Gy�;d`�t��m�Љ�hFT�n��Y��(�'�n��H# oS������hG�鵃+�e��V�u8h�(597��J�b�0��:�k2�T�U�&ѤK��e0,C�2ד���-�����=lw�-��k�-�J4�<�[U@���X-G������f�P�N����!J���f�����g�����̰#E�e�-��nea��鱛W���7���PC�?w���o��>�i0/P]�4�_%"׮�e���^U��y,��usy6�W�@��D�>vc��љ�z���S���O�o �b�N19Xws��+��Qr{F2$�w��'&`�����`B��Aɾ}�)$��2l\{�y�E�%Y]�{��S�*��)3�J��&�"�*�͡˼V�c��;�^�=�-H�:~#�����z��a!�N�v��kv��Eޠ7��DX�Qr3>Y2t���eh!��-�l�8v�ڝ�@��
���n���b����J��Oӿё_��(u�)B	�fj	��"�=�cҗ���׆���`Z�T��l��m|�S�>WAg��u/9�~2";n#훚!G�|����RY���L�"�.�UoKI�b��6��ν�ii:��˰VE1��ߢ�x��N���B'{L�C�$�<|�j�	�}iX}�ь?��8 C!��.W�a�*�9B4���v	�k�?��x����UvP�θ�R��4�]�� 7S�����V.�;HxF<e:��y������3ĸI,�;����R(�����'��qF�[��ʎ>K�_���N��-
�m�QPWpn� ����K2�LI�
�?;��)�N��9:��9�5�i�$�t�%+�\jG�Ҽ�vK�M��5��ȸ���8{�]���G4��a� 3��@+QP+�M���\k�-�ف�Sj3�w-���Zrj��M�suW�g��8L���
����P�w�P����o�#��Wp Z��I����%M�h�Ҳ��"�ћ�3�_V�K����@�V7��Z�N��3Q�|E�F��9�}����E�G��p�q��$K�>.�"�>�ў��YޡH���(�)�}$�ض+���%����Z���P��(�c+B?-���"cA��А'�B����[�Tq2�0�>B����W׋?���X��2��	�~�No��7F��ɥխ/-#�H0�ȅF<�};r�wĵml��f�;n5c�G(�K/������'����p#�r@��,��e�p����-����U�ULY���Q��ھZ\6P����� '�1����:X�0�x�A��ͤ�"�;�g�5��#����$aO;��O��aP����w�š��JA7����{�S�'W��a��E<��8��U|H�źctTd5��DP $N��@Z�{��W�zH����� ��$?oo��잆^N;��T��E������b�&��|i�-����ߩ{��2v�F�j!�'[���ts8�_03�x5<�k�g����2j�ӾH��`T�g0}��a�H�9�T�s4��XRr��п�m�3	���N��8�*�
ui�n�f�K�_ӫ|F�Wm�t�T7�����{[�QH�`�Ug����\LX+�Pa�F�k��v�S��_�d��a��"=iJ�Oק�&��!�������>5V:nd�R���p�K��+��ͣ�4���?�G2��iH�'���kԮ�����q3���o��L�t�"-�j��7F�?8���L�zRB�o������3^��e��3ʩ��f��݌i�'фDD2�a���uyO�;���&�Eg��