��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0�H�0q|x�F�Z,2�6���̘7ш�)�7{<j/){��$�Y8`��,�U�^�4ԗ~�#m�Dڂ=FX��>_ߕ��+�X�cd[m��(m�L:�ȍD��Ӫ}+烀��c�I��f�����ۏ� V����ʦ�B����Kq�pL��@�	Q� cǁ�2�Bw��d�*De�&;��^��5��΅��9��@E-)j�W��8�vf\�@�����s�6��uN�p�Z1���a؆R�Na]U��0-E���������7�K��Ĺp��yÚ��s�X�+07�����gj���%��C�l\n-�)yT��((o��`�m�+26&	^�f?�s�7~�(c~����`/v��k�$b��G`~� �=
��ݍ���������IH���Z~�"��e��-WE����b/m][iHSVHy���-���h����b�u�$��t�e(��cB.�z�&=��&��T��l>+D�ȁ�z�����:��b7U�?��A��p�T"���[	g��Zh�I[ui���V$6B��?-%	볁����e��ԭT�6�#
ɗ�+S��ڙ!��
~
p:�r��!�[ ����\�p9�/s��6�E�s��4C�v��,��T�P�c�Ԧ�."��q���փM �~�V�ɚj���!��UBS���I-ʇ��j�m��-��YvBf˒��Ma��g���KWʤ�9���M-/�b,���-[$@���{]gA��T��a$1�#9���a��#_Zt�&�>���ag��Ry�$^ܙO�s�E������huR�/�]�¡���Op����)3�_��-�$� �����:p?��3�k���<���5g�S]=�	V���{�<e,�5�k"�+�����b5t=�B�9t`Az��y�)�����ʖ��������fÓ78�Z�Ͽ��r����v)�,�/h��) �!�������:6���$j/S�#y�����9�-A��WfL�>�*�ۋX��5V��[�F>��O̕�V����}v#o�"G}�r1u�"��Wzև?)S��� 11��I.��BIt 5N�,����.]�����(�Ȼ�c�v���׶�5m	���a>q.m��W��?!S��3��`tC��� ߦʂ6t� �3ՁR�P�M����b��y�0���*s�	���3F����QR ��fL�8�H��>�n?	0�Xa�ե�Ƈ
���rK�Z�a����M[�ݯ$X�fI�.`���#rm[�Q�_� ��~�P11id�cƢ�_�e�������涆4a|�!.J��A�~�H�4PO�������3+�ԾH��4e{6�ߧ�?�>�*@������PŚW���Ő��Y���7�~jJ����jؓv_?	�~c ��|, � �N-.�#5SWk�F�+O����yD���ox��~�Ð����{�T�5����h�k'�],���@<���B��_\���L�T�L,��5��eO���"��Eⰰ�\
x�V�m���!"��q������+Gw>��g��*�{�B�;1UT5�PΡ��h���0H���Uz�kʽt�E}�8�e��ʇ��s�\s(Q�*mf��#B.n@�8�Obȁ�jr���}ߔ0J#I�$Ep�#y�� �a���'���«C3��^$k�N�D�-"�}������0'L�Ky5������6��#e���Ű�����ԯ�6����N�T�q6�rt-o�2�9�.����J�bx	3���c��lD)�W	ޱ%���.H:�X9�.�~�����\���1��3n>�I���r���z⋙76>*ɴ�H��4i�S��y<9�υ��V��#5�&�L����Q [ZA�F���1-��Pk:O'< <��?��I�>K3�EJ�1y�I� �n�@�\���sX]�C�fŮ�p�ǝ�����T;�9y�PW��������^�u��ܴ�~�;&�����5xf�p��֕/`�}�Z^_�e���c��3������ `��*,~P� �w��`��0����j�(n<�F����� 5�Q��5f�6e�uҐ�����\&�/��dǯ���_
�
�;Y`w�g�U�O�]L��p���)�@��а�"��c|�ӈ�V���=m@����3��2R��5�3N^�_[�������77���cc�j��u��Xz'�$�_��8�?'\h��u�׬����l���u��3��n?��["�U�^�E�pp�'�`���+	���O�q�49�dVY�
$��.G��
<�"hT���MD�!
��������H8Qz��Ey{������,��l}��H+n�{=j�1�����ex��[ �j�����~�=�����pQbL��+k�	�3{�e�(�I�}6']��{�um��8�ۙ#���j��p��7Y�ܛ^�@"}�@�k2�dtV�@�ri\]�8�i)a��8���Ɯ*u�ru�R��E'��Y,jqI�� H��L?n���.:p~��>;=��n�J_HZ�k�TO�	J��?Xq�K��۞��3(8��ee�L��el����?��;�{R�0^X�]��*`��w���^�Vu/� ����_?�Ql��h��.W���ʎU1f�;U�ٿ}�Ȥ�Vy����X?Ĩ<g{� (�Qp��BK���Kc����>��E�F0B4��O�c����m�!�(�`��W�D��W"A�3�faו&Ҿߧ���E*!��yi���tGqy���vQ��"��k�\�tޕ��|�y��?4/��XSR�6�p�	w����0�Zf2e��F����)'�����
d'�����)�U$�ZQ�y�.����	�%E��ת_�º$��4��Hᾀ�}W_���vЫ#<����|kǱ�Ť�[" s��-0�0ô�͙?�u}S����c8�L��Ƶ���D���	5�R�s�.����y������:�y2�H!�u��̼��I�$�ŰR�����!�J_H�����×5�t��d���j����֢��$����"�]u,�T�u�~��J���6��w��8J\_��?�jq�HAz"��F,!sw^㋠��>$���baJ��|��6�I���>�2��f��3�P0��zl$񾙗���C�F��>�;dRZ�⨲M�M�tG]ѳ��6�������)��q�a��-�w=� ��7\"An�*kE8q��F��t�:��
���WP(/�_�.w�9g����*A��=/ɷ�ݩ,�;&�AH"�@��)��B�)@�-e�����Ӱ��ae�S�f[Y!3D��L��`Qq��D�|7�.���T�[V��J#� �����Pb��'
�r���mv1�m�"/L@N��Q$NF�f\�Ľ�My�%�&��V��DٛJ��Z���. `�D`6&�t�L����Kq27h/v��퇧u��� =RS��{/��O�)R�X�}�:����k�P���(2��(�Ի|�PJ�^����w��Bepp���}��s�|�t��/��6M�/���n���玉�PL%��k��w�¶�΀�u�I���<*�<��'��Ov��h֏	���V�x�ě�Q��w�sq�8��j��5�Ł�1��H��K��愃�%u�5�j+@&iч�,�����@))�X��]�Ox���YV�	m�!�Uo1�6$�mЩ�؂�C�ݜ�{r\���5hh��$��hK4��.�힥�NS"U�q�N����l�U͟�l�n������n���<�J6�����9X�j_nRq��|P�z ��N���7X^p�d�)�e��},į����c)
O&v)�|�O�ȕ���M]gEoHq����0����G�qa�>�h}f���e��P�s���:o�=��ϸ�^��x1���BIE�)~�R�-s���r�~"���������є׉��fj�ESr�47���Mf��g�STo]�����W���L���5"y1�4"��l�Ն��:�i��G�}؃��foǈ*�`�3`�I���{:����Om]�d�J?h��"��'tN+�@Q�e�Īa��Fs)֜���,~��3�f ���R���P�cxb-�O��,�;�C�F�|'��1'Q���0@�}��_W�5$	ԡ�JTüS��/��w��|܍Fc^CS���%z���t%�8�����_���t���4�
ù{��<R9x�7��G�mbp�5BV�*�ߏF�:eMv�$�K�� ���j�Ğ��l8�����Jrt�}V��'
6,Ԭ'��l��.("}���~p�_f.��9�-b��ZF�5̔�z��[�@��nEJ�6�q��T��xJ0�H`�X�m������sfi�t��Ө|m���p� X�����_6���s @'���Ѐ;R��v��=�W���U�oB�N-t��u�mIA��7RG�jץ3,��3�a�0�3�p,�ʹe��	q2�}��l\D��ry`�x2�ٳ�㼴E\�Wf�(O
1R�ч�,:�&L�'@%�i��ɽ�_R$jZ9�OZ���[�?�i�t�"��-��;G�u�H�{!�{ì���6!y��Q�sZs7Or-'\���h�V�}*�X����?A1�� �Q.�^���M�`u���x�:���z܊]�h���>&g�+Ò�:����&=��ҭX.�y[\̍����㔐Q�,s����V�=�e�
����}Z(�EI]�PK��Y��7줂M���E�aM�q&E�d}��/0� �w0��l��#a�D���2E��Om�
U��--4���@�w�Wr�Toj��\���`�o]�#CuGƃ�!	��ڲ�^W���j=�9��'��A�ůVm���u�Q?y�r�<�MD��x}�!�ر-����5gRovs}Ö��Hp�F$��mfs��B��A��OF,�yC��۸�1AER%꫟�&W��?ҵ���(^�,�K��h��Śwѹ����ƨ�H2XD����@���d��S��;LN�ؔ^�a�'�q����%�OFtNU*��呔�����bn�tD%$f"�c��'�Ō&�4\�����p��m������������ �����>I�_���š%����+�n	�KE�sP�DY~J�/��S@n���Z*����1dԏ�g�DXނ�"RK�g�Èg�,(�,�=�����G(�a�S�������\���k�d���>��I���F7��sЯ�`�°�%m'����~�̍���:k�?���{x6zY��螉��ȕ��$g�j�hN.v��z:Ӕ bB  Bw$d���/��H9�W��9����~IB�0���3�q�P8��46���������ܿ��)A�,-fV8p�C'�jQ�`N�no-{ͼnw�UƇ��bN�|��l�E��*d���+�t�O!���TwΗO�C��g��������`׍�}N�]O)#Sg�'��!o���^6�y�y������|P�Ͼ�m��c#YL�/����n���!�`�Ȁs��V�P� �5>3Qf�kǻ�z&P/�BQ�@�b2��;���%=e������_&+mJ���٭�=��E�Ef_��NE�$�0�q����Lv���Y�����[K�<�PA,�Ϸ@52����m�ɔ��L4Pda�n�[�s7�6֗��X������K�Ǚ�oY�� ���xO[����|�DW=��ݮ/��@Z�7뱰���*����
˱��دB��H#x�����ٜ�s���%��F<HE��/׮���A�<SE���^7?�`��f�"�C!o���܃k���1�.��]�ҫ+�?��D�Y�VB��pS�>}�#��[�8^�����;"�dn*�q�(B������U�o�W���|`I�@UP��Åc�ci�@m� �d�����y�����s0Sh��$D�L�$�{Z|���#��Kb��1�[x�jJ5R������q^cC�=c���B��pm��_[��Ir�� t�b�pW"(�O�sX\ѥ�!΃��Q��'񯌗8l*�d�c�{(f$� Y����"�
��m�ߺ�ƣb�7����07\)��5��3hM���w�R���]� >
L�F�]�������[�����%"�GS����7-D��v�(!�.Ss���ؿ�	�n����������� P}cN�m�˫�XEFܠE��u�<z�ٲ�R�$�wu3m��P�S�0Nh�N��S]���B�]��ǅ�'4w;MU�<�U9B�He����Io$���h#E�o)�u���d�Ә��6�i���!���qQ��J�\�P$=[��;�рp�er�@�0��[j����T?4�른Q����5�e�$Մ�u�%����:�<`�ES�ǡ��R�vw_�3'���+��KUk#���zo�r���-TI�q��i�5�{�,�����1�Ɩ�L���.!}�(��a����Z��h�T�"P�C�� _�]pى�6^RG�Y�V�j�֔����� r��ftxĔ��V��D�
��̐t8CK��V�Px?���Q�R��0�`���lt�l�`�k8a�MW��Ʌf0Ɖ��v�`�k�u��$������m�Ex��bf�b��a��V��+��o�R����\���wDY�?1cԵ��ۺB�o��$�@rJ�"5^�;C�<�v�9�F��3Ls�f�Ey���}7>�DeeC>,_��w�?�;Z��+��6��wL])!���ά� p��M&K�5���'\2BW��� <��;�,���t��V/K�oiH���j�t�k23��=�)](�U&�������#��2���o(��[?~�{9���(�j]t�X]��o�˯3�\X��(�$90��������k���o/7���\W?���:�Z�sU�����G{ w��c�V�O��#�>�V���ZB|�^�)(�����=X#+ګ��5�����duX���C7Ƽ̵I�f1�i��U	E!x�������^(a��l��`v��)����E�ԅ���v�=Rd���\���r��t��y-��K;�h� �~Ӟ�0�WU��7�E�;��Va��7s?�����GS��.�z����v����!Km� �x�C�8�
�5���Y���g<ST�Ɍ�Nl�x��U�J��g�A:�c�y;a�(���u��e���s^������*ha)����A�+�R���t4-�B�]�t��,UҜ6���1l]v{
���͑�BԾq諶C�&#�/�u���b����\U���L�^���% 6��x��<����*�?l IQ%��/���;1�6��۝�ښ�@D���sSYӹ��lY�BE�����_�1ն�����"��M� �"��u�}�,ߔpsЇuҍv�4g;+��&�>�!�0�M��ya��.���Ѳ��!P���\c��r�$&�#�֨Æ�D@�P�KP�R��9㯠0��{�lӸ�V��߇C9\$���2�'Y��7�D��1��B"G��]�07�(-=���rP���F���p�N7�����$+t�Q����
H�K�BѮJ��C��v�ם,�t+f���h��ڕ�K��Z���|`��aooKp�Ta1\���8¤?�1�9�	G%bȭ1cC����ƌ�Qb��cnR���a���Z�bQ6�$5�\v0�x�ad����!��� vl�Em��ge.�3��A?z�A��Ϊ4�ֿ�hsU� ;R��%[��"/v}�<�����BH��~�U�܊#�]8��"�`��Eh����=X��?Xe�l��)X߈B?��`|M���I�P�-]cӹ{5���1^d�8���)�����6ݣ��3iZ��O�vn���Q��,�9�a��2�������R�9\z�
��"B�j������Qh�� ��k���o �;�s�;Z�����*�̳�b)w�h�����5��Y�!�}�/<ֲ��}�Zp2&9�-tH|�2�T�A5�E�F�T��k�'�(T/�U$+X�K1KG)�Bg��qV��2Z�V�U�v����&s���N�;�e��O��(�^�W����Mι������,.?^����2q�1��C�J_V��� ���.D��6I�fQ�rW�u%��k �wA���� ��D�r��O�&^��ֆ-�潃�*o�d�5h�I�z�����n,��kMOD@�G"<G��~�Xҷ=Ϻ��i:��"�l1��P�F��n������V�'`��h;���_�ބH_��w.�gl������N���"d?|ٍN���}&[�T��+Q�����{ �C�t���X�O3�D��2��L��2(�i��՚�,!�u�|V�bgD��� ��Q�rMNM�X^���*�����2ZWJ��1/��a��X�ﷁ_i�
O��ȫ�,1���heC��d@�&�&�n�X\ψ.�](�םIL�_��n|���+mZ���f�D�n�^��,V�9���d�.�0?�"�͔��q�J�}��$�l���Y	AM&﮺��pȭ4�C��Ұ�d'ǝ�-f�`���f�e�ߎpl�@2Ǝ~|�I���2*�ny2��ѥ�z*/��Z���2ܖ��덁<�`s��N��8�O�^j�.��+Bܒ�L�j�0�������(�x9��n�f@5����ig������f���B���rw�tF�-�I���B{�4!�῱�-�I.��#�Z���4ѵVw���*j(�!9g3p�7"�L?ZD�_h 2n�E+#i7t�
[~���W<�J_a�XvJ��Q�=�k��/Y���u��-	lė���ɼ;XS���[%{�]��@��K�$�����0�����<�G����/g�8��$���jzo �E�� F��9�Uz��������B��'B�4I2�[�i��)��\�����9��\-�n����s���Î�#�jT��s�޸{ɜ{����񶲵�t"���;�~�W6�.$��oR1�h�VK��c�uhN�����Ě�ὔ5����˱�9ә��]'C`q��V�*єS�sb�Pu�[���o�<�8�$��
�_�O\�`�,{��H,"3.=�po�����y���M+98G�a��bFH�^����H��W*�U }��v5���N�jH77R�Ps��m92������sn-;���X��ugtD�k^��n�Iߵ�,�I���{+m�*����1%�"8�RH��V�I��7��=9��n�B��Q��#����=,��[�P� kuԤ�}w��̀-�x6d7hk�z�sd_=�^�Nv�p:�����yƦOjD���%�≠��V�7�6nXH�!�[�,Y4T�4l�k�3��]�s��}i��1�S���\y�hZ�h0<�8�f��VT�s_Xhy��:Y"���y�3���P��@X�������T)�Ǔ~tw�+��{���u�� +��jd�ѓ�j�+|ƕЗ�ǋ�K� �;$+Έݖ���V��V?�(�Qb�v��M���4�LnT���Mv�v�3�˜���ɿ�c��4%ŉIx��	�u�a����ZR�[ӹ�L8>^���g
l�����[ϟ����/�XS��'A�;��+ޥl���
[m_��V����Pm3�xIjY��4H�\O��j�� 7�=Ί�Niߜ&���|��ԛ���W�%��N����\}��
�4�+�˕�#���6S���A����2�5��H��i4j����T�2g8{��j�ڣ�U�;�X*hl	7�!F� J5�O��7��ͦ-�J������2�˻��p~?_��}r�� J���|���c�[Ӟa��w)�M�`	+n���C�=��`~���ђ�`���e�^���qvvײ�j�̮�=d�^�W���SHb�TPJ��6�0���f��>�'�Bg{����iЎ	"�z��v&bo��wP���K�9
e�Z�Aqxm��r|T
�T�
]-A�b�E�SU�:j�hށ{԰u��OYAiS�{�?koD�=�����.��=3^��(-�= Ý��5����y1H
�W���>�/���;�>ofp!�=-�`WR~�e�~���5�.���#e/E@�*}�glI2���}E��^+!�:��j�I��Z��4�ѼB�^���	֞���_z�G�2E��y�cz����=,���!��0� �l���yh6����D�8����R�z��$Ĳ���nKB���~��_�/,A,?���LxQ��2��C��1U��Z�>Z_�Z72
	Q�Ǥ�'%�@h��S=��A��n~#�}� �ϥ���'$R~�Ṱ��6���E��J[v;T�x��4��{�E�
�&�d�B�I�e;�4 ����c�0��:;pW��,�;���>P�L��p��T�E
��ٕA�=�&�Z���H6���ǩ0��}�EO�O�����_dL�$��_?)ǒ�ʱ����ѷ��?HyW�W��KA��OYԗ�׸ΧݞنP��{��b^1V�%2 �Uv�*��h�f!_�/k֫���0<Zrs��/~K��=d�Ӕ�L�lE����E]7?�� �Y���~��?6B&X+��+���6��Z=���!���-��=�
x�xDSB�Z�@ǵrG�ڪ���Ƶ�nT!���CN!e�(� ���<qw�lد���K���j�͢N0)ӊ��|�����7�/c��F��Ǯ���:� ��pJ���8�[<���W?����� 7Ez����Q͢�ݻ�c�e�	��z@Q��$G1�-<=g6��a��{ ��u8f���Gj~�o�$�"4!=z�H397�:V�o�̽��M���@m.�̫18��㍛��D��HVZƙ��� �Hލ`W�����\��~��~B͜��7q:�ԟ��S��V0��%�=� _�S��U��͋�Eb�U��y[:��������x/c9a�H��ڠ�*ݍh���0�孧�ό���$��*3�ҒB݁X�Q����L��A� �6��Br�l��(�~��z�F��s5���9[��4�v,���l1,<+�=�3���=W)tC���U�����)��`���Nk��F
�ܲ�"�R
�|7������PT}1� �6Dq��T��B���}Z���p*�?�����t�;�i������0�0*`�#%�9�'u�B6�߳���&*�����>=S�mSEQ��W�����XQ&b���)��f+#�YÙ.�A��$�������������rd�r��h����u�+ʣ;c��[��V�I���+���j���P�ELʺ�wW��S��/��]h4^=���07��~\�40a0MvC�/L��;�T0�N�{[x���v��V,�J����7���!w�:���L���r��$�*����ϵk@���.Z3�E���:#�|��qM�E�\9k��)�׶S�b$�e�M|:�%�����x��O�����?��-+b(���m)ʧ�`����ɍ���"fh�O��$��ts��c* �w6�G_U������K�2A�?
�d:�Y[&�fݰ4�j����9�D^ρ%�Q#�;������n@��i����"�����?#�.Wo��7S��6�̽�Ґ�PZÉ�.��myeХlpFw���̪'�XU�E?���"!�����?of���ϔJ?��B6��|>�O�e|Ӣm�F�ı�8IW������h���T^��B�����ݞzi�rko\AN1�;m3:�g��%M��)v�m�ʲ[���v��E����W��		�h^��'Vi�y,����U�Y��x��s1m̕�z�	\gge)��0�7.�.�G��,z�K��0<��db�������!�&ecfv�I�*��z��N�{/��/�f��w����x'41V��h����Կ	��y�h�=.��������Mr ��@Y7����}���S�iʛ&�YMYMe�x<�
},<�Wek�в4�H�꾉`���e}��c3�r䅼(9�'��c ��sv�,R�`$n�V��� ��������&� ¿u��H�m�Y������b�.�g�,2��DL����SAq�k��3uf�!�w�يJ�ZG�':��d����vſ��	���q�aY.��,rp(��܉Q��{����g٭䷗W��`Q�Gem�r�<yb}�B)��uh��E��B�:U(����Ar73�%sx�.]AZ�k�O󗫗'Ͱ��-�����!d?�$В�o֙�s֑�F1Mt��$�J�	�Dj^�u2DW0��~�$�\���?�䧨�LW�����WoP'�c�Z�M�Y��W-�lŹ���#�-�é�$P��jrbH����0zc����kcpm��zy=H�6:�Zo���gл�e&ˇDHU���qkE�
�5�� ��{�N)\�s�|��a�����m�o5R ���	�a��-l�(��+:�d*�V�'���Y\�G1���c5����6ʨP5a.�V��B����n�;���EA��1�bX��G[��W�Q@�]X���h�-��D���o�i�����*K����=�����Lr۶7F�q�)b_��k1F$8{]��Rm���u�F�����[����7c��]8��x����\K2i߆�קJ��$d��?w��C������a0�I�Hԙ�6��߸G~3S�����}e\R���XM��}#�^"��3��u�:р�ѩ�\d ���H�5^b��C7���E�s���0:Dx�w�[���2[ݴWtaz��]��-����0����� ү�4�"�Sst��}�3�~q֢�ї�TaК���`E���/�Ћ<�K�`�� ��?�~U�V�D^��P}ϰ΢yc�%S�D�m|��w�w\;��ɍ6i�O�8�}J>�P��\w��Q���>N;0#�Y�mh����y&�d.�0"[��	p�c�槰�H�'+ŕ�}OM���<��C��������؛۷�\!I�'ͣ��@�\u�������5�2���w� ��f>ܪCݤÕv\6�$���/K��tIu6N�^ 5���y4���~�w�sӿD�YD�T3C�/W�(DFr�:�_�QJ~@�l��a��鶱)+�_&ϻV-�LX���?��|�;�b��#l��1d�!��LD� �#�[ε���-5�|Z�����9R�.9���@ڵ���O�e���= v���c����ۈ���s�Eߘu�q��tr�ӿ�C3���tb�#k��ؼ�������ϝ}����9ڐ�*�]����X�58���ӿ'Cy=�;l�9�K��l˺n��c��۬ɺ'_�WM���oc�$j��[�p���rRB�}�}u*���2�O��e�*�+W��.`��p�(.��Z�����q��[s�֐��<!CY}��S���`l�i^ʇ�ͧm��`e���O	֗�Лnk��G@	���l6{s��U����U��IQ ���&�P�]���Ti�5َ���@ɦ�Ă�{5��3�@���G5��W��4?Co�M+��&��lq ɻҕ�f��*▁�)厜Ph5R
���8p����Q������ھڭ�ʘ���p#��11�J�P�Un���;��0b٨伏�T���?��wX���ie*=Ns�h��#S0�����:�(��1	�,��I�D�;�l��ɪ@�Og�hv��hL4ttB�C*��x��l-���{�{(!�F��)&��N^Ù���2�%���x�ɗ)�/�'���%��-�l�,C���z��b�r�x��r鯠ȝ~K�n����4�'�ŀƂ��%��͚1{�1Y|(گI��f	���XO4��&$�0����1����"�l�d��R�����-���������B@����b��,S����b�e����Mpe�>������Q�:��!���ղ�Ŕ,_l�b�Zi,p�L��U��4Fk�L�.\騚A���׻��ɝ���8U��n}�'��d����bOT������6_�f95+u�ȸi���	[�3�l7�����qH79ot�v�ו�/��q��`/Z=�w�&����8�\N!�Ϧ;�I�C�E��1������s_�~5�]�j�l>ƛ*/��0Ќ(U�ɜo�
S�"��z���a��avmz`�}@���m����M�g�؜/We9p�)F^N���%alg3ez��ͤ�h���o��ug��)�Nf��KK&��L����r�c]R��޼�C/�� �h��?��=c�v筒ԧp�e�=/A����y=a4JIVK�h���ek�=?�I�N�Aj�J�5d� L��'@�?R@�n3@������.�f���Ts��Z�xo�;�wI�7',i���Z[�޲����B)���ii7"��Rw��	�0ؑ5�5��<b��2ד%�X���'�-k���͟�6L��=�	�>@b{x�t�	f��V�����h!�ߝ�Q!�ŏʏ!�6J-�ȼUPp��|�3�)���qS��ܘ	�1W��c�[�����1�>%���\����~�ә`Ȝ:G�Fa�Ý�n��I%`Fy�^���M�x�F�S8	j�\��0�����Bݥx�-��lWnjn~�<tR'�_�m�� �'��oR?	M�3:�V[�җ(��F��@!)6G�i֪s�8DI
X�����(uMf�Dz[,�
�9Tm�H�i̽�7��J�ǵ����|ܑ�~LC~���g���T���]��ہL�U�Db��/M�p�ۛ�D�9~�fZ]P�_�ޭČM;)�q����9�
}��Ca�k�$�g�"�$Þ�`�$����t�>\��ji@ A�IPE��޵Ӆ�a޼���d�Ռ��b����qh��l���&5����Ԕd1Ģ��K�"K8`p�/�i
*>5�A�����W�g����o[�'��xO	�8k�R�4���!�F��	'�J�#t%	*�zw����xET5G���DR�F.n9{�a4��K�M1���ѓ2>�� �Eׄ d[0�d^���ne�#ה	����ny����f�AE�<
�/ {Xd�X ��y�x�	|���2?�s�86q3�qS�uJN;��@���s'�*.��G����褋��J%}� �x�< �����0�eZ�/fsH���W���|�R����2�Br����N6 �I�ݔ���mՉ����Ki���� }���`�8�9ʀ;Q�}���-Jn"k
��U�dH�^o�E �2!=F#ߏA��S�c�y����W]�]į������D;��@��&3�;1u��:Z��A�X���b/�,�	�����y��J��]#_�U��0Z�xR�d�Ń���pn�����K�!t=�u|�x1P�q�W�ALK�C.��%���ܱ��0��o�2߶�P��:y��y����S��#�$!�XSS�	�ր�)�fOreYn�a�Y���҉���I���Џ��L�F:a�&����ŏe�4O���b;�ۏ��60,���خf7zU���In��5���9(9��٘ǃ��p�E�'ɍ�}w�W��at����M��0u02r��F crX6��=��{>��2��}^t� ?�GR#Yl�G��E�M&H՘E
p[��閵�0��q��ˎ�W|dY(��>Xsg8�b�?r�{o���T��kM�E�AW	����-��$��JċD�>���ٽc���,(���`��i�T�t}�)_�Xu[9p�u­����jQdXf�Z�]s�U@�D"GZ��ˑ�����M� jA�7נ�hkg.q ���q����'g�� �`��J��T��>r�_��M�u��:��z:!e�_��w)>��K�3sݪfk"�`�U�y�V
jd/ J'�=��	ʵ{�ʵ�P��U%�!��9���q熤	܁"@�q�ܵ�S����:����n���$Ѡ']�}���G�Au�&�ƭ'r�AYC��j��@^}qf����(3���꒥��M,��1ba��Xi~����ʙ��y-� �E��jĚ�\�[��-�/�ĭ�ˬ=��&7SP���@f*c7���;AT���j.I:�*r�z�4�|<�ߑ��`�����Z="  9�3h3�[�gP�j�H�i�gy1���h��^\g?>;1bi��C�����J/��(k�L�6q�j�q�2��.ㆲ�W�б	΀iMv�[j�x'{��N��T:�f���+�Pj�]�*A�N�h�<1O�Ğ��U��/
La�7�X����+N-Ȳє,yW�.��Q�}���r�ZN����"����mId��%�5�r][+������:�.R.�74��L���|rK��H�3]�LT�B�>���FZ�nL޲��I#���(�JYp��"�$#$"��-o�9��������ê��.%�hrM��G��xp���y-+PR{5��;�g�Ŵ�ܱv1We��������B��=cbE�����'c��Wc��ߵ�?8�w0�%w:��2�/��Y�.ߓ��~�y��b�0�(�B��+ܗ,]k/ȨX���_�^���^��TE(�!��z�M���j<`��caC&M.��G���=�p�/���ɥ����D����\I�������j��T���[G�_�\UQP)IA`᯲U:~I�yd>8C>�>��I�����Q���mÉ�?JV�o;s݆�a�i���
�	��E�l��V�Kp��F��n����!�6����k9nG�u�H�*�+*���JOU(�kh0"�?͡ڭ}xg&��U��V#ԍ<S	���A��π�J.�"�I��2��M��/���5���F��� N!~�������X&X�l��{ـF[L��d9�w
L��XR�/.U'ז��\{�g ��_���}8�����|p�0�� ~�&�Tn��z�8��?�C��)3��ʧ�Ts� ʌ��Q�[n|�)�Fy�fU��l��!�����$g)"?��j�O�T���-���*�Aڙ�cR�x;�U�H����Τ�mj��Z��B.{�#�l���D���dܭ�#�.������/^���L��q"[���k�nh3���A��t�]kGJ| ���P+�G�[<�}/�T[?	F-�CPA�k�MD峢\���R��x������dJ��d�!�ú2�Zvm�����6���t�	ʵ�W���/�b]�7���%A��5���9x]x���s�`����H�+J#�;�ʬ��).���������v@
�]��-�5<m��3��l�;OY��U}��v[MQȎ�p��>IW11w��>��K�l���$�N �7��˖�0�Vq�Z�m���I7JV+ ���&�Ś.m�����B��N��A���>��6J����	��?�^�TF�h���YR
g̶7<'@fO �����1�:�����;�TT&�MDk�LY�x����2�Є�'�1�O���-[6ȋcqմ�ŏ��<�P��u$�b�x�ﭠx��F��pH��D������I�����l?��F{�D�]�*�]�#ti����n񋸁F��q���f�)�&Зy���j�P�0p%j.��x��-�q[p:����� �/Xc��&)�g��zC����[��9��϶)��uu�]̒�S�U<x��"�veN(2gb�ѪMM� �5�n`��◥��k* ��X�s2�F[��==چu�m�S��RǼB�Tii����-���t��!T��*��3&���Bm��q�����O�ޱ��I\���F*�����S3��g4���?����F?\c�8M�P�x�v�
��p�,Pa��Q�� ��W?ܾ\D�0�2ӏ��[�꿪 �!ep_��|��"���2ybt0�!��ɤ�Jb}��;��%��3'a�t���AB��Rԉg��ə��S��'���/_M2UR*r]gj��$7nBc4���O�zJ�����%箩��]0aS|x������v�V�G��)n���ȣ��1Zr[+�ev�p���Zd�S6XJ�y(">A��j�8��/��ؑ7��?��kE�\�'��>>Y1���V��]��E�ql��c/�#9{�JZ�֡�ꈲ�_������bP���T�O���PA��'LDY��hc���罾B�ߐ/���iv���:bV�i8}��qI���9�3L"4T�&p��Y�ܮs����&쾇����=�IMz�LR�p��aP��P��W�^��,'N�?��8s�]�J��u~���א
y��p��:��T���Ǒ+�;,���3Ӓ�8=z�]��'(��D���ӿ9�AwX�Snm,/ҥ�o.�V�Bf]좮pQY��k��y� |�KB�3ȉH����Q0G�(n��"��d�l����)��hm����%����Ҷc{��4��K���X���j�0�8�8n�=�{�En��,�N��}gh3�э�N'U'�Qo�C����[Ga�����u�$�<Xa��L�-��R��>2K��x�d���RCo�1x�V�O�mu�l�\���[�ڐ"=S���|���$�.��c�E�L��(�,�x<D��z?$�%�稽��mI�H輤~�FJm���A��D���2˒���tYu�A���;-���T��;Re���xh]uӝ�/����p�Vx�jT��gf��Wѥ[}֝F"q�hx�����"�1J�\�Ӿ ��M��l{����*Y�&	^:S��/�9]����O�����U�b���&�$f�>A�O9V��#>:o0��9�^����X釂�pz�D�^�s��l��)1����bl����ء���.M�"l���_ƌer�p��b���5���S�I���ҖA�y�ё9u��aS�X���c>f�Wj�7*��+�
�W�ب�躴����h��u2���o@Y��������ЩO?����c�.:�Z�k_���m��.�#8���o�@���
9�<{EQ�u�)ސ��R^PlI�n��
{�Q��o�Q��W�x�4_ȧuR�vs���vjbC)5j�^)���:A�Z Z�)�$F\��E�mG~�'˓Z���3����U~���f�y�����	��s�eq�m�ɳ���������Z=����z�:�V��3�sy����d>�cA�w��o~;JQ���@t'�Vqt�f/0�l��v��Q�f���VT�t,�־�~1�d��,=���W�I�r
���P�X;�_���w��-[3߷��	A�B�r
G�7�XB18j���$bY1����=(�wl�Ya��l��-����s~��+"�FɹY���H.M�c�S��!<Ex �$�亨��k�H͒I�R$��:>ߌ�"��P�3�izQm��	xX���g��B�d���t����T�_P���ww����7��x*T.����5�vً\�Q-��]o���݌y
��:�=$�PĤ<"��j� ��L�te8o���y��_�)r���z�!�1�6���2�{�"ĭAt{��L��'
�߃V!{��/�4�T��Ef27�4�J���+���s;Ih�>L33O�T�[�[�n>}�TB����U��%-~d �I��A��F.��
�ۆ9�̘[�_�Q���8��`J��I���ߢ,ji}Q��H��ʎ)��~���/%����WyR��J-&���V�p]4/���M��uϨY�]!7NI�6ʁ�oq�I�m��'�4�9,@�"1E��D"�ڟ8�ݸ=�buI��ϨnmlB��6+�H�ħ�/ԥ�)M�|j�����AP�[A�.1jT5߹ح�{xS�b��*��6\cI���m7f=bj���E)�&��渔��F�̬�����T���ƿ�U��$D��%���-W��L��`}*(�0p�[���}^Ш?��V�.dqي�=��ks-��cDK�ܽ`c���߭"��2��J1]�d�m�>��T�����.��Ƹ��T��u�n�ϫa�@fF�U���$���goR ֘M�YK�^p���Z�>��Mk��P=��UT��4~�J;.�J�ޝ�P�ӥh�@��Mt�i� '}���𸧸�U������G���]�n�C w�t����3r)�+ض�<
2�0|���6v�P����4��9^m/ч�t��u`���A�,�ca:s��"1�� M�!�!�j$�)`ޏ��>�N�O}��+��VXP�mβ�2ӒR4��9��H�LtP��&E������W�0Z}c�(1�Cyq�]&O�g�y+C�Mh[����G(�jB{,��f�+�.�-�]���B���M�������;���	�EIa���%��:�EչL���@�M�wȵ���9�Y�ưlw/��S>nɦt�W���U�2[ z�k^���_�~�1e>��hPzd� �ɡir6�0���*q����G�8��1D��h\q�~�8��f���{���i똴�qw���PAD�*�ٴ�6s�b3u�G9l֮��e���Ħ�����;)�:���4��ÝƮɟV�:�^�;�����1��/�#��Z��d#�����4ߨm�f����ʾ��+0���z�w�����6�����q�LXj��C��M��|���My�t��7u�$,Aq����J��K8�ٛ�{�L��>m��U�
h���Xө�����^N��s��ט7��^zk��[m� (��"��|�S�e�.���*uD�(�5�ǽjk�j�Z�1�� Һ3��#�\�դ4�i��X?���a���OEr_N�Ɓ{B��$0?�Y�ʳH�{NWD��ř�-�b(���ɖ0c,��Mͷ:⻈��o� d��@��H{�ƍ�ߍ����bbOӰƕ��d�_��ts���Aw����Pp��0����#�V��~9��@�S��_�	�����HW��챗�<[��&u���bC)�|�����6R�Y�;<#��RhI��UT|�" ���i�8|E�76d������H�x��V_���0�/����`HƊ���`	���U���Q���i��*̈́��%�?���u�A��H�Tl��6��^�9���y���T	�a3���2�[uzmY�Σ����m�8��g�Wb	��y�Ǘl0~�=�0�8�t��}+�w�e�J�^c弄w��v�X���)�w�m�r��[��������N���栦첀<Ç��U�n�NkΑH�H�{W�a2�NOT�Z�(q[Q�� �h��g�
PD��!��Ϛ
���1��za�7��x)�v����$̢��cr��Jv�I��Z�*3 ��_�d D|�E���N���U)����mv�R.�l�&��h��-w�RB,	H�v���<j�ֈ;B?�	�ݩ�O�j)���ډ���`D�> ��R�?�"�)��U=�h!�?Mc�6�*���H��m��c��{YJ��f�iXi��":���^��K���L�j	�H�5j/#�{j#ƌ�����A#�!a0�ד5OtO}���f�&�)c�� �g��7��
҂)1_��K.���s�a��Q#�K���o�D%lH��)ڮw}�p�����/�EH���޵p��X�³��H��B��U�w��x3���G4P剔~�[nH�,e�ㄝ*ꗦ����|��J ���;���Sk���"�3~W�h�{����Y�?�[�a'�6d��E.�����H��q�֞��ɂ�:؟_�qB���'��CL��{����׳s�ɸ�hNh$�[��ۧL���.�0�� �4���&�)��Q
�Pt�������"^���q$�5��0�{�&�G���п8�A�L�Ǽ��`�?�׎�����a�[�5ZmlCΦ�b��._����'�a���#\p�3_(E�JO��g�Z����������G�ѹ!a�Xy��ŗ}B_eZU�W ��Pj@�$��f��J���X�۽�XQo�6���TeF�1���^H�����Z�!�B�{�/������ u@���E�۰�D@ϴ0�,H�.O.j��@��]?��)����ӕ�!�/�N����Q�v/u�8[��3� �~� `����7���q������X��l_f�/	�	�1���<����h��/At�J�� 6�Q�b�3�;��q��eO����{��j��]���7�d(<��>��g����E��خy2��X�av���ư\���q��������C��yAYT�Mw�N��Fէ��O�7̟j���&B�Ze�Ϭ�I�>�5ri�q�{��6����h8iI^�<�`4��'"�(�ƈj��zm`�h�E���I��bpdy����J'?�ƭ������|�M50���X������)##$\�~1�z}7��tsm@X~���(t�Y�n&֊��;8���L����:T��.���de,ŭ�{:<w�	�#�_��w����}�ʹj�R��F֦ɇ��T���	T�w�iNN�L�4����EqV�'����� �7�a�[T���m4�m��]�	JLNI��z��[��.��0|�
�o�U!˰��fҰ�}Ϋ�8�LP��/�K��-`y��ܠ{b���v�TU��U��)^��:h;mQ��[[?�.s��ͣP�8��
ہSWIM^���
FO��"��CWl
n�6K5���l��DAΘ����2ǒ_��ʿD5�dkMϼ��p�i3��\T�˜�������p.�P����;�*�X�}Kw���� ��h&`����ӎ�؄oK?g
���
10�,�k�Ն
�>�T^#-�Ø�1�U���aed��9��$�.K�
�Nl@W6��#��Ӫ3�A@R���_ðV�s�R��x@v��� �U���e#�U��Ki~�=D����!��[��S^xU����P�#�N2 �k����MG��My��x)���W�QwN>bV���A�,c��I��<8�t��
�>�c��%�șoDո�L7*>S��Kb�(媧���i<ұ��$���(���㗈�2J�Q)%3;�7O�Sp��qk�����	���t�t�ڊ�cp��;Y�`	5�:
A�
�#��-/�{Kb��IZ��0.�hI����Ms�h`_�9��6�<N�>*3�-����=%H��ñ]�n��
sK|����:`{��?�%���4�.)�!cVq�U���6�P�\�����"<-@���Ʉ222��R�$�ǡgk&�r١5sh\��$=Y�e��񳽯�H�/5�.�>r�ލ�}�8�K��<li��w��]D**�p9��ɑ�ʆ����ز�O�=���xΉ輦�B�r�8d>��%�s�-��
y�Tl]���2��!��w����@R�/� ���B":��q��D
�xzN_X��{�er[� �{��/&�kלk��R�w1z �J,L��QBe�r�f��@A���OC�����D����m���,!�o�B���VQ�E���]s�}�E�1_�x�ǧ:��Ӹ
]��������F:�O�p�����3�$PW]	>��*�f��ap���(��!N�)��v�|֚L��*�]^9�(��g+[M��{-��A�s@L�L�ΠC��f���D8�9޺�usb���o��5�¢�iB}W��_㐮UI�H��Ӓ�4b��h�8=4t �z��k�&�|���Џ��AZ��;ʏ�2)�2��(����@|^]�T���4��p�j��3V�V	��o}�Xa�4�*W�O(�� �.&_�@�`n�ik�^h�k��e�x^�%�ŭ��XS���X��'��߆Rr\ ˠK -��!#'���M�!J��d�o�!�Nti	��ůۗ.t�YL7�*��@y�18����g�4��o)"�ܮT��&��I@z��Fm�):�8Wğ!F�e�ٸ�b{y���Eo���&�Ȏ�j�\�I��� j
ޞ9TE��I��I�:�K�Kǌ�T��~J:���QF1������9�}b@�K�s�:1j�ʧ��K�W�R�ǞǪx�C��k�T��T�7�:{���U���*w"ٝ!\�H>[5�	��[>��@ڸw�*����֮_�p9���^_���$�,�N.:�Y�����ʫN��k1��͙'����o�L��R��ya�tSQ��CcT%��s{N��F�z �73����?;�%��br�A�?r��Sp��H]���B�=<X�ή�ۈ�i>ן���'�rTOd~���;=��P�M�X��b�����gUq�Z�%����������g�{��9�I�X�M4�Cf���Q�&��0��`��b��c��O�uӽ��X����B�~�b�W��-���ntnC�	�Na�^�-�����G��6���S}g�jH�!}n�6���BZb����8M4���r����3^��)0��,m����N=!P�k��N��!_ݭ�uA\泍�ܴ��H��۱R�]R?@؉@��ٍ��sE���5^*\��1J�qUu@�l��n���?�{��`}�_�)��̠�!{�k+Fۼ�i�T�.�(�0B3Ԏؚ�c	��]
=��X���t6�ʰ���m-	I���3؆=�.E4�㹆e\�r���r
���_��Q��1�����I�g�r}����;z_Gy��ĳ"^�d8mӱWFw�Rw4�mv���Rr*'t+^��I����5E���ʴ(����[E����t�#!�ʹ��BelF[�S�(Jlf�\3Q�*;��v�)�t����+(r�aռ��)G#�(O�G�*��V�lc&�̷��,-�Ybc�v+.b��4�'��d��ʌm&�kgۅ��KU���Bף�x�U�4�Ϙ4��wb��ЂmY}Q�؟P)���ljǈH�o�0/�n�C��=�.����M�����2Q~B�͚�jM�q$6��eBK�R��n�N�3&�V�m`Ьkg�5=�z��iy�s���JP���0� e� t���Q�\�?;�p)���U>(�������0�19swQp�G�P��ݫwӗ`�Tq���ߕ@�WQ�g6�;�&���X1��U��|�r�����ùWǜ�$�W��2��,>�>DA�0����7���?��U���F������{=�`3I�*9g%a|�"7'5��M�É�?�;؟0�*����� 2	.~����.�4���c�(\�'�NdO�_QȯN���>��HJGU7��
�*��+PAs�!d!5��o�U���ܡA��?I����!�l���E���c�${ȋ5-�ߜ�0�p��8?R���}O���~[�:��@u�zP}�{jIk'8ݒ�Ƞs�]Aر� b\f��>�9�B^�e0�[�3�8t��F��z$7���C�d����M����q'���T�����d���k��=w~�	
�2�ji�y6�Qy�A&@lѯ�*�P��
�T���0����d��Oe�Ł��!�̞��"�Ki�_�}����]�����9Yʾߘ�7R?,;A�A�}��Ky���~�n5B�9ƃ���U���N�{ItT,�C���É��"X��s��C!'}lb��H\��}Q�#�� 	�����`�������$"Q¨_�y��S� �YPtU�:����U�K3�$�JK�(��8�A;�ې$Qr)����?{hg�	X��96�aP�$	���E����Q^��T�U�v����@��헄�A���Xv�� ��i��3�e��*�nG��c	bH|�MJ��N��z "XMU�I�����������)](M�<���q����1~Vg�!����"i\E|�4p�������@m���{�q�*je"c}p1��7:�&,�C���1?b��Pꃧ�ح�"����l�����O�z^Cڗ&�3*R�mjyD��V= �Eg��G��k>���\T�4�H16��&v��[��֙,�;E86(`�io��Fj����R��T��-�m�B�	ʭ62���������؁u%�b��#¸�Ѝ�'Y9����u�ٱ$& }��{�
�}O$�U�����[�"	��秘KU��V��\c��@ާQ�TL�h����ə?���HKA]uV�Roaק�o�P,8l�8��Zqo2��=�NI�)��b�.�Fc�-P���_���d9����&�?�`����s���<��μd�E\M3�Q �'��[���L��5oY��j'�j���r9��+��C�HI��WV�r6ƙ��w�T�ʳv�	dII-�$?PJ�ʣoZ%]v���[�M�[x^��{M�ny������731�bD�����M�2�� �v3���j/�����Cjma�K��D��΃�@�$v �S>��g|�g\^^9�B1I g�kEiӰd��!�:�g�{���%��o⺄�̱.��Y�s2~��Sew�6I��b��M�=�A/��^���@����e�F�L�Q�i�'�LY¨��X�oU� �RQ���!� jTfČ1�QJd��;���Io����x�w�p�/�)�e�V�s�DF�r��Bݛƍ��I��#="mߠn��������ȵo��o�x���F��7$]+�	�Ց���;�/��S+�f�� �b��յ]y��w�~5S���<�:��9�}ċ�5w$���(��s( ��Z�*���!�AGWL]�����N���0f|��Ů遍����lB�a���U(�k� �0yb6	Ə*�]cYr�u�+�u1�P�C�`b�3�C/�[�2tK���%=B"��ɣA�x��h#=6������'%�����>O�g������:r���&������\���(�[m�1Bk�Pl��!����ky�B�+���#4Ʃ>�7�������+a�p=Ib�]%��rci�xF�"���j��(c����^X^�硜ژ4��oW5��G� ���nf{.�@d^���L�*-0�ϧ�u$�����U3�H�=�(i��	���փÚ��эLG�#z��pi	H^�&'K���J,,9ʀ��q2��Lz��2��i�!Ǿ�Ѻ�J��1P�5EU(F(��#�`�^���j�J�/��.��2�}$�q�R�C'E>�Sg������c�3ǆ6�ɰ��'wAß���7��D��X�A]�v����1I��7K��C�!��[_�<Z�^j��7A�(��a��g��+��/uH���.$�T�:/X�.E*#J�}cgTQ&z�D<Xa�k��t�8���X�C�f��L���a�f�y�/��/�3oq�M�°����j�E�"b}$��7�`uJ�绁?���dH�����O�4�p���	�$��������Z��@Av$�,F����q���>߈����l���c/�pФr���s�v�$�pI�mo^`�(�	MG f���ż;Ԫ���0�?w���
p�wH�%�,3��w�aie_��#�[��ךkt�`g2��,
+ѓ���Q���
�j�pϠ��@����彻r�ޘ�G��g!�����>���Ō4 2��/C�i$�4�9~5��n&"��p�+������O������\/_b�_�2��Pav�.��@]���?
 ���7h���`�L�C�q圹�F6�慧�|�/ֱ�U��·n�p(�k�z*���";�a�c x�u���ta���7C���y)���E�솼e`�d1�\���l >*�Z�T�9W� ��ӱ��y�X���(��M��wu*L��D-�o�!	ޔ
6�+l�=��q�M���@��̈`|;����O��]B��_�T��ƍ�?��O�k���\Y�OyM.�g@�gP%/qx\Á����+�<��b�w��|Pb�ӎ��{mSʎ�Ż7�㖚Y'�g~9-*8��F��l���|W�������{��N�
��$�{X�c�m�͔�L}g��G�3��С�����z�-�u��e������v���K�	��m�7��*�ww�-�+m���� ~���}+���i����j��]U��JːѧX9�S�/�0��pԠ2�s��3��$�	9���3��O��j�O���#�3Y��r6 �M�򻍛/9b��	RIճ��UP�������	��F�P؂O(LH4q�%�@���}В_s_��7m�ě�qx�S��+�?��Kn�Ŝ~[Hn����[��
��+�����v����kW�Х�,��\B���5�����|Q�xF"�MB��E[��=�Y�|���$	Q��쑇��*��%�Ȏ>I�B+�_+�
�EB�<k~���λR-��lȯ�|S��,8���b�nCF��Ǖbp�\7�H������x��AG���Ӊ�RKW�3�\u���Y7�OLv)^�w�R�TuVo9��ܜY��X	�$&NYq�,x���Im�T�����3jU���te��co���G�!b�B�M�����k��=��?s����j�Ó).I'm�%�FTaA2��g5� �Ȫ����5NZ�G��-!s�oU�)q{��]"�2�/x�4V�f ���v�8�{����@3S�(���jkL�.
�h�E�g}b<�5�����?2F���i�2��� @ �?�F:lB���~���W��$?�
���r/���7��x�&�` 0�8x12�H^�r�S��5@`REV���]��@O��e��R��Ҹ�E��,�~p�g�X��� 	��炒rs�h.���d��H�J�i��[�d�A���k9���Z��(P<:U!���-Z�WP"��V�M��`'�Ċ}ю���-��E��CS{4A���6���H�i�c�g�K���w��Pj���Y����}��+p�,��?K���w�h.��ޘd�>.2�0;]g���S���:#<���Sl#yqB}��%t�����b����[��)����o!��n��U�`;w�2��
�S��@�)��@=w���F&ه�΀w�)J��p�[
Ŝ	�")g�O��((qF.dF�u1�Rn�;�7.�!�ki���?�sۡz��8HK�
aE<z��3�e4>gm	�t@Y�n6e���ށ��E��~yP��3}\X'jo�vP���O�^��<�kJ�yg�B�Ӎ��7>UH��fJeΰ����	��i&��2�B���:���}�)%��"hx8KUb�$-
�+5�hݛ�=,Kyv��z/��nї1oֆ
�D'l��(x4�
e��嬭j2A0��p�!9q�jΡ����ShK��&p�ci���0u�Ư�MC1��n���g��5��W�Vײ���3�zL}z1S��'�<s���;Z�:�=��q�`Mj�DTi?��o�N�v198ZH��{9��W�t-���6�	Vlug~���$�����Z���
H�$�Z_�"/�}�2Mc�6�����u�D�a�C$+n��m��vw�h��L��x����%���p�I6SXc�����lꀆ�S��~�TJ�vXkJ]V���u���ڌ)�t&H��7,  �܆�p�ŖB������K��@T��ְD����u��vl���6�6�z�-2��U�U���n���(�Æg���*k��z$��b��@�W���c���+cv>��Vי� A6k��5 d5,)F=���Ʉ�.H3O��Dd��%���k1�D
>w��%�+�������?E���,��:RE���.� Y��Sl��[��Lpo;.��p��4rנ4�8�W� g��K��&U93R�����*��MI�gh�yq֢1�۪�����>�s�X�u�}XG��v�A����B���l�iݮ'>udjn���mUJ,���O0�1k��b&�@#Q����	��� �4 �M�U��Hk���F��e7;�uX����S�S!�ߦ\UY�g:��
�x�]^��=\�!�ŞT]��iW��| ���#��CƄ�~�j��uSO��t�&߆I����F"Lx>y�堮�}���q��u�n����G1�v�B��
ϰ��B\z��e �X��9���cH-�ɘz�e��H�*_�{�a�;q	�\�5Ri�z��J����g�"/	�M�s����@φ�x>oT��AR?�|�{I�F�0x#�\ @��R�ԲSt�ӫD��C;ǗfCU\�A3t��yN��r�y.���9*����5�4�7����� ��¨�wP6j�f�y�$��n�}�84mvG�x��w8�-�NԘ/�(�]I�F�5�]8P{�` /���o>������O�鹸��n7��*��Q-�J��.Ĺ���Ǐa�B8n%������W?�^ ���*�O���&�@M��F�EF���8��7R�&� 5�? �;>S��|��T��\�u �JL{�ҔM�s:�M�X"~�eue��|���s ���<�_	�$3�
��|�#�:��ɯ��aD��R���E�(���Y�uZ�/�}|N�h��#�tƃݠ�2���Э�A��0��	�����*����� @ψ�/s� ��,��2�����x��'0֓]�J�S��u�n��A8�]��y�s��ܯ,�F
N�zJ2�|PeUv���6 M��66�x�K9]�Gs�v(uo�	`�jn���	���=��	��x-A�WHܔ�����4�`l!\1�Ӊ  o BJ�k���4@vm�U������ቅA(_yx�(���5]�ܲ��,p(�b�-��J<LVnf�dű�5��clG����-_O��T��QX��h�=i�:��[�l�*�W`o�MK?m��ZΣp@Sɧ���%��NW�$�Ѩֶ/�vSm=o��GϫC)�p��U(��*s�/םm�D��#���G��3q��!�4����lo��$�Є��09jr����@��ߚ(��h�OQ�;w�f����6YۺOb��E��U�<_���:\�Y��* �� fRb0���F���C�0��gO���HTۚy��% ���Eᴿ�-/e.>P�jÊe+��d�鯈5�%����J*b�B�Ή́�)���y��|�)u��~l;�{U\�1:��2=@`.�ka��t5t�I@H���+|��aej��@�1�y?����@��Ue�c��m�R[��g�k���V�H�C��"a�R�hi0�t��P+<�c@�X#e��6b����hz&������%k�I�20L��ITj���*���N��Kw�wSsDە�J;�m"K�߀=VOw��c�񗴥�XC�h�Ha>�*�U����e$�gV誘U�KT��UH�v�BS��$���������wqW�D'NM�<�vI�������߉9�I"X�U~��&
�iX5��������@�E��l��io&����&����^h3�P���n	��K�RKw�M�|Z�z#j˱z�	s�;o�}�E`��(5��c4�������?ɶ��24Ѧ�(�����>��L{����FUڻ/R�7u�k�$�_��D4�w����&5�`%d$��]GA�5V��Q}T���z��:T��'���Cq�����K���z��~�aY�o�|�ű�\Bx	���+R�y���k��%kV�X*rQ� ��r����m�R6�_/ZyEYD��^�g����@S9�c�l=PɨG��>	&����_*G7��[|�P[?��Z{��K˥_�:jF�d�L2��iR�Y�Q̝�k��Ku߿8�x~��.�jJ~5VE�,&RU2�VO���a�����4)w��%���^ۨ<�S`KbA�v�r&$���/x���1�u�k��y�����p�"�qs�Z}
���AD���޵sZ[�|�Y�������l���!�!˧���1��H_��OpWa��-Ġr+J�6�J�Jx]
!Ř��/@��u�o����0<����}l����M�c�����Eţ��n!��C�5�I(@UW��p�>�X����F��s\+�Q��8��K����خ��Yӈ��Ge��~R3x �'��u�t8����k����(1X��a���Y�)�3�$f�(����QnT`�#��(����#6��)����:7Tf�[�g9E�'O	�]����%r��5��⮀�v֥yv�Ft�����	�f��ư��Pކ����*BF�.�������{�:�UZ�(��!�ۖ���Ų+_mI��Q�նǔ@�:������E��-f�ҙ����d'�������]T*���Q�;��2n?��@"Eq�M"]S����Cu�Me�CL�>��P�e�@��n�N�&�\���	צ���,��B�4�$_�@?k/h�eG�Ĝ&��K�#T~��8�ӱ�/���N�Uj�|-ت5|�ڜj�O�69�EUڭ���0�9��em�Lr?Sm�'F�e��j�?�2T�+�٫�#�]��(؉����ӡˇ��_d������U����F\��5�Ap55g��P�
4�q荺6x<;���ԋ,a��lI)܃yt�$;�9�J(��\�p�,(ڎ�
�V�DY���O̜��`�TIj'�:�W:^6H�X�"��qu4(�7�o[Y�b1΂!Ĩt�4�)���Z�^�9q+�k(4�mU Jo��-E=�\�<�~)�z����*n8M��C�~nq%��&�
{{���F(Q׃+D|�7/l-&�X20���Gm�P�t�f�T�q]����9eF������i;Bg$����s�:M����9ńzA����E�f����a�m�3���g������Tl���=^t���R{�7;��4�ͼw�0g&YԸ�o�7�S���{;��c+��5֕jϝ���;~�n�z4��(r�=B[L��Y�b�Y�Ȕ3�{��k�%_e�b��@�n���d��*�C���NV��a����{�؅�#"�L#�Q����3l����,�����lJٟ��#N�N��d��c�q�8�����p����j����py�T R��]�R�]q�h_�87��K9D+ċ
��x�6,Ȳ%�>�?���}�˭�F�F��5S_�G�	�8n
��r���]T-$4�U��D�%~�z��sL�#l� ��#4�G���`�Tk��-m�5���Z� 0��93�c�t��\��{���~�
��[�v%���͠H����2�s�:D�!]rV'%&/FiW����{�_��0a��Qт��Z��Y���g��\�f|��A����0*^���ߝ�zt���v�CVoM����8B@���ޟ}��
Xu��ι�Z� X�g��`��e�;̯o7�~������
W<��� Z��ג@�h�l�������}���zx�;L�P �� ���F�-��y��H��^F�?��G��������l c�S�H�m�v;�p���ž���1N��SG������{�dNL7X0���6P�����L��;��>�^{ڑ^�7\L�������C�z���дj\�I8/�4�
�2�.%^W��%^~� ?���"�Ox��6ꪋ\�OSG6�vn�ݻ�-ׇ����{��vC��������AIɳ&�b+V���q�6-�7�SV.|9����#�#��5�v��B��Y����\�ȼ����Z'��+`c��j-b*l�_d��c���B �KD��~���%�b �K ![� �x��z�Df���m��A�V�@=�/�o�/���`
�76��C$K�n.��o�U܇�\�2�g�Hh6�.=�TR�jM#JSp,G4'C�S���M�̥��"����2�n+�u�i㻓_b�1�WW\�A�a�
��"����׽&o�p�Dn{䙍��vD���Io�@��ƿ�<e�W�+K,�!��7c돮|�u���#{w��Qi��0�]S�\n��n1-�!�+e��̳�VY���ߖ��~���35}Q�ā��n#�1��/+�|2��l�.�wZD[@�R<�Ő���Mx�k;._�M���J��]Y;=�O�m�OΒT߯���OƑ:��v_�#�=M��U�gԽ։�Ձ�(�$���U���A�_�]C�L��Y��y�7�p�ƛ��{"�$��>#^3����l ��h��Zp�����4v��2X��S��[1.����

��6K��n1i��ar�v�Z�������=M/UGo1�I8�5J�@��t���i�ӥ#LYG*�y,�)�za�U�>��f�>�nTa1.�"�M�g�m�2�q6�+��3ɤpZ�+b��$.����G�� 2�X�����B	S)��7�v��(��Ŧ��~���N���R�̍<d�1� �?jMD���F&W,v�k%���w��Y�M�FN�25=�!4ύ���ײ��'�+_�4���/�mN�JO�R&,����`g}-����Ә@�j��~���YIɢ���hJ	�:��=_�N�P��B�����V�y�X�$�3�$��>�q�i�ٵp���U�j ��ᱱ@7Q�L��A{X�Xv����|&͎���4`qA�#����:{�6�L��>^�GX��*�C�{i�ݯ�/QD���,˨Z�B}�/7d�L�2���'�*�=Vۼg_SeC���:�D�%/�|]%��s<S�.@��y�T��]^So�G��
#P�p�fǸ���.c�Sf{���l���e��&�v�vZ:e�K�s碾�'ƫ�ѫ�L?#���v�y��E��;PA%�Ϋ��)��u�kV
U�U�X���/4�)�]iA[�a]|H!�,�٦�ve��q�ҴU�eE��G)>x�8]��ko�j�4X�6���\M�ܫz��L��T_���U�#j��1&����
�/�4�v�������^�r4%�*�f�(#l«n������\ut��@��'�l\���B�C扨�l����H�o�c�O�J�c�!=�y�Yl�gg�Հ��N���g0��2�k���؁*,ަs�<�'ιI�$`�8w��4���4��5nx�g�ſ��<M��8�d�O�3A!�WTZ����W�O�z7��q]�#5�u	�9����y<:�>P���6��'�D]g�FE<Ѱ�$u���r���+�o{�0�nu�|���cF~|m���"��"�&�������]Xl�e �s'��qv)ّ6���U�����V{�v���R~��������"����Om�}]�w�D�5P��h�{S��4fK���AH�T�3�����>��|F�.�67yG��q�Ɂ�'���r�a���;Vǂ7\���������(-�<C�l��M�#D2�� � J�������25�G0�e�1+@�gͬ��b$Nu)�֛��Ժ�=��2��C��Ip�e++u�.���ޟ<8LA3��ȹ�Z����>��܊�+�O{���
O�vQ�o�Q�Ŭ�փ0���0��EI�c����q�_�1�j�h��q�I9x�I7\T����њ|*	6�?l[�W�RAS����$.}u��T����Z��F����vy��W9>�ǒ�9��[uu��� ��<��M��˕�!Ӏ��#�j��
a�-�(+�!bP��q�I.}("�SJ�Fƛ��g�͖7+ �x���? +2��U������Y���8���`��L���bی�>��}r�ʼ���&��0%!3�y�
�)�=��0�����=Y�����0���W�ϰC~�3e�Կx��>���_�c�q�э�uv�N�|�B��)�IW�~H2Otӌa�B
Z=�\rz��»(� �x�7��f_|��z�	^��eīqPv;�����LyЖa����J)Z�����Rf��-+`H�'|K/�� ��zsɆ��y�kI�8M^۟a��Pz���{��V��4r�a�Lek�&�"��Ex�}�S]p���W�9�ts��_9�H`E�5��&!O�	2c���'�4���Wl;x��Λ�q�,����	Mi!i�-��؈�QFlש���Hm)��B�i�d���н�T������PFd�}���Ό�/��dT!�O�Ы�q\!RjʉAoEbP�<['����A�I��ω%�>���Ƀ{������i�iN�[C�6G!�֝�b���%%"����,�8�ֿO���t���b���6�2%�xw��w�f���H�#hߖ�I��7s�,��>} A���0oay+��cI�Ǿ����>P2F�^hR��,���Gv���$�.k�8��#@�Ǻj}��:���l�z�hȥm��V3����[�#�7�Ɵ����8Z�)a�q��{����T�rC�Fv��ExԡQs�����z�
-�|_Y^�^p,/w��{=� ��t�4&0O惫#�����NQ8�fJB�r������~�W������L��/��9�ڪ%qem<�vu�BƟ��Ra�b��d��Ds�+')ù+K�Ѧ`�*j9�A�)Å�@��x~2�b�/��B��RI�B<2ߋ���H5��zX���w0z��l0����G<�S�im��#����U������!��3�R9�o+�`�m���̏���y�&�
|��}�ý� �5�;������75���o�Q�g5}�v~P��Cw�I��D y�3���m>�1�A�Y]�J��I;/�L;N^�>���T*e|�W�~���
6y�."�I-=Ժ���C��\�憷����`
�ah��<�~'2�ctɀК�?�b��7��9��S�bSx[i�I�]�?ͼ�7K�l_�A,Z[�n�  ,sR[�=;��wëIZl��t���w��3�P��������AQ$��	}�f�n��lR����b�JWkK���Q�z�g�~SdT�HV���{��Y�s�_?�4��cB9�:k���ro5�n�{d�s����
� �nDa�α��qH8�Tz��{���/T���@<sV��,zd��]8}ҁOE|yy����=7n@�f��_v�G��S�x��c���g=xU�$���=b���"����܅��)A �=��0��a�$:�-�����V5�ۢ�*׹jf�g�I���(0��?'�����i�7��ӡ~d�Ě�.?�H=@p�����xy�$�.[F��UJu�p�9=��C����p��N�Pq�Z��b��p�l�V]Q�t`�='[]��I�\W1��|�*,�	�ZXN�7�� �ե�����t�7n����ըdU�τ��<{7�,$i�~�����%����T|��$�\��m��ҡt�9��F� �{�ŏ�=�'%{�H�D�+�z��˚�+�fS~o���wp�����'z,w%=w�a�S������z5�p[<�������_�(?疵=*B.�e�C�Pd�@����>��-���G� N%����3Y0u�
R0T-��@��V��
�#^H��]l;\��6Q(W�,~O_�!}�-\��R[��������P&V](���Mc^�@Ԩ!�&��s��mt��>i �t����J�6���,hK7�/D�)r}���Ib_��������ہ�o'��Ky�c����,��D�9�	#�*3c!�h�� �9>�/[a�e,��02["2�Twn�T(Xg>ܗ���{�b�+WVdz��(_�A�o^���$1Ӓ�	{A1�*Y�/�Q����T�rlπ�?�m�b�]�s��œ����m���g��VVbߟ�6��ŏt�R�w}7���r���0�����K|�*cy�fԮ}�z��ަ*�T�:�Ò�A�')2v2c�����cs�!42C�ƒ�Vw�N�&�3e�Eb�2W2:��:Ȅ�I,�'�����_y#��pz��܃pQpc�>�ܵ�y��ֆ2���$��Dx����x}�ۅ[�k��3m��O���*�@��V>�ȹ�U�)C��D��g=������LLp6��Q�$q���>�;�j@�fu�ݘW��H�~rԘ�g�U��4�7ry�#���vt��v�LV��i���|�KDB���V�bg��.9��5ɼ{G�\a}�*���I>����-/HjȺ�`%�I��b��P��}{�2��(=�����z:?�69��RXe��/4;�`� �~s�
e|�Q�4�"3��i�E?��)���-?5��7��u����У�L��QG������e�U��ϥ>�1p�y��L���h�k@��"ԓ�w fB33w?񌴵�>Y�i8�好!�!<����]��l}�쯀�������g�KUi��ȏ��U{��k򖷠�����]sg n����y4@����X8�0C��s��=B[�"@*�#�ݍZ�Zw��Ζg�������Y�׌����۵���h��_�$�z1H��V�(��%pv�sM��t�J����#����am�&:��� ��C�6oն����X�5�ƴ%��S,�}#N�k'$ڪ���˵uѫ,�F��L�Lr���	�vm��#n�D�B����Q��/B�m�o����G�î��⺶��_g��/��C)%�J%[�'qr]�\��oߵL�k��f�K��$�0�-�
+!$��j�5��Ӎ�*S:��B��sv1��GY�P��k1Қ�4����V�Y�L��_޵���g���%
���蒼�����m3M����M�'Tnd�����%� �z�ſ�R-�[x;u��XMϐ�h�A<z��H��K"w9�iiG��K,�@�Žβ��B3t�G�i��U�>�
�
�Rw
�S��~�����e3�%Uf��T����"�T�=�e�i�Q�`�M
G/+C�]��X��f�=ȯ��=S���5���ŒY�
� 2w�c��C��:X�hܡ�������/g���#��ͻ�*�O��`�M2ϫ�E@C�y���k+��� ��n�o��*���#[�SO�R46���G��1|����{ �~����i���TkF�K#��9M��u%�r̃�I���1u�����4Ha����HaZ�74(��BL`�׳�~esTc�����!�rmָ����T�DNF)��c�c̺�U'�������x��@��#�c4%F
o(�	��.=��Y�:�߁�� �*+<{Kq�����K>�8j�Z��tdA��X;�d����̀(G_j���{x�h��Z��T-�8��TWq_!U�aZ0ңJ��s�f�	3E؂���li1�8V"��޲b����e�w�
QN<"4z�$��΀;Vc�16*��(9�V ���!O���1X	e�A�?�c�2;��ᬼ�8.���.<}z9�PɮW����5�k8��tX�G�[�0m2��Y�WI�A.ٲ�[�ǃii뤜)�;���k���儰ι�iH��5�D2eEa�����}���{q��L�:Mm}5�7��z��d5DV�E��N׬rC������+W�]�Įv��d�Դ�>��g�����W,�KϽъlZ���{�w={$-͢!�@���ȯ��h��uO�)ÃqVA�4j�v���J g[ sS[6�O0l��4H��s���X����b/s�4F����H��M��YS�� ���ϴTA��9s>wkc^����vs�	��d��j�\�+_;F��*$�Z�����͌�'��������]jpfi7�ײ�ſߨO�@/ج8˅�̵	�!u5Y�b�0j��9�ԘJ�I�?I8+�{�`���	��d�G\�P\1D�Y~T�{�>8�ۜa(�w�7��,A�^����VI���r���;GV�%V��i�|�7aN����RrP�����#qۤF�YP�T�8���d��Zd��rXM�������sf�Z	veU������{o��ޑs@�c��.9�t͇�gC���*m�J�`o�~�K����,[�#K,I�����k.D}v���F�:	HSJ)���������"�/�Z���ʚ�N�y�[�re�5�	�a5(Ō���0�U���� .qk��2��o�鈋��&����So��at<�8�-�>6�L���J��¤Ɇ`�[���Z��Pa���������[�X���}�f˯VqƲ�'^���Z��4z����VQ�K��Tn=:�Ԑ��>,��Q�:���c�>��_!vSsc�:�'���^ ��r�'�rj��Q�|D�B�}-����dHNZL�`�ǯ�X�<�Є,2q=״�*�9��˶�P�)ꚈSOe��������ۊZ��W�NR�Խ_�C���襀�(�6������|zk��+�����Џ�瀫$�hLA��T��I ���h�9,H	����Y&�+0&�d�yѽ2�h�4�?ְ��r��qA����Y̝��fA9>��M'�O/�"�"
t������C����z]/��?�C��?��d���ā��}�F�>��)�:΁��[��vm2-{��]��OJ��S���T����Ţ̢�ĻW��F^䕨d�d��u����^�o��B�)��(\?����\.��d7*E�C��z��Uli.��g�EU��w!���!b���1�����-�嫊b�G�8o8:��6�{g?��&��?�bQ���A���R����-�j� =U��ff;�K٧[@�����5:�Aq��c�Q�Wi=h��<Y�"��q��4�[8���f��i;
Nq���ɮV����+a�����Sں��G�hO��4i���Xa��$w��&eo����=��	|�㺎 tօ�	5�:��p�w��l.��ޕQ�m�Gݓ�r��Ǎ՜���(�n�~�Q�E�?�X��L0T��O�̭ ���t�U"}]�xK.D T����c3b�+)>���&U�����*��y\�-��I�k�'� ֱi�I�n�8ɲl��٫�:<��'��A%�pG+Zs�#:в� �ݪTL��X��^~�q�I0��J*)��Qh �rM��
�e?����
k(�Q1j�`WMFApO-QS73��a+X��z�7�>T;�FϺ��+?d��OO�T�!�#��,��+�S��+��a� �d�_t��QzCǃ��0���_1�hټ�6��$��,#�~���O�/� ��M�0����s ��s�-5$^IS����V̂�a���ӑ̊�H�Nzͫ�12���&�S�vEA�ǽ	SK�nowyҥ5� AS�1��'��v�+����}�o"\p�	=p��%�S�W5�����|*,�Ґ�_w
O�>�e����m�(�4K�~΢#u�=�Ǭjw԰θ}�A���U=�k��GK>�aͽL�Ts�-Mfl�1�����6����x^(J���!
)��8�I`ς�帷�J��+� P�_8�ȍ/���!`����;�c*�¾�=���M�t4Q���ʠ�?�h~��x�W��!��pB+^S���2y���@�p�{/�ƚq8�VP��F|lC8O��{����|����Z����$���&���lwd���-�B�mN-f�\�ј.�bD3<q{���: $U#ïn�w��0��X���s������C);�N0@��
'1�y����s�&�<c>ݯtJbr2W�X�i���?Wp�7x?��WV�OM{���sXu���6�)SPM�O�y:3h�Q6v/�]J{e29�)0ø�]�����K�4��X�X��dzV��0�����`�:�Ry���
E�-&7O����y<_���Q��BR7wҋJ�Fv�"�]2:���̳���+U.g���n�C�<�tz���ɽ��Ū,���Ų5|}6�= ԍ�]oM|L�Q��eX���1��+*����й�=�s�ZrY��./���'|�H@�}i�t?�vB��)`uC\6x�r5��l}��ښzX{-;#u H�%*� �Lx��	��C1Ȗ���:�<��*"?�Nս�d�#��_<�^�3~*�C�Ya���X�K���n�p�(�CJ�i���#�z�����:�8\5�iH�m���c%!k��F��e��^��ƫe�y�Tc�^b�v�)4����s�)�{cK�/�y��<��!��s���$ؑ �ӳ�W��}�� K�fF����Ǖ���e�dPPe�E\:6ř�����?��Ħ��Pq�c�\̡�ݞ�'q�QV�@�v7��:���^!��xfs�\W�c����!<<X "�Z�S'������K|����4$����V2�#MP �>׃�KZ:����7����)������8�-�&Cd�~ͤ�>{��(��b�~	"�k�.=�Jx�LhJZ���)2���]�*}y*i�o��A����,@��;���w�c��̕�g#�#�٭ȷEG ;��Ն:�pG��ׂ;"�������$*)خG�Vz��Z�г�l�E����=��������7}y�I�I2�eKw�uX"OWA�ڃ)�z���9ʱ{�QK�蚑ґ�)��: )ʐj�"]Ǆ蓗��3�3�u�;u~���Mo�o���|�ח\��6��#sx���^��>xր��J"cՊ�!� 	(%�/-���SL��]m/Y��d@��Z�j�� ����(BOΩc�Y��A��fp�<ok'���H��H�o��ǣd���
3D�ldum$>˫�>
�t�+i�7D
�u�����?��n�I��z1���
����!1�d��Bdf؏L[��qlk���*�DK�[ZU�C稸�]O��l�`H���ˮ%�`*��p���rP)��[G��
��d���,ѮH�V%�#KP�����)� L$��Jr�'
�e�?/�Hؠ8�-��:����މ]t�u�ҋ��M�:gSs��衍iӻWK*>�Ѫ�B�<y	��l�)���M{�9{���S�]y���G}��\=b?F�1� ��l�ޏOsV,|�՘�;�,��H4�_`��)88����t�\�燫��6G�M��m:�+���귳{3ic3���<4fK���4���{ւ��h��X�r !!��'Oj���	���B�"҈��^"�w�l�&��d�y6��NO� s�]� O�k� ��]6i�d����bG��7��My�=%p�}I��?�ϸÉ�;���S;�3Y6��-:YlL�a*fv䃒��!���Px��~a��!>���3���T�b.�V�K��u.5�G+��t-� ��!0�x}�nn��+�Ȣ|yIU����_��8 ����"��S�/Q�UT595��_�ϱ�m�d)4��߶��&�Ī�̃�:���s��G,S}�nK�?���Њ&�gbʁ���.S�h���wQ�9�U�7�^,/��l?�3n�6�����^�m�l�Tc��4�Y�8�d�K
f<p!��v�<�8K(��J���j곉%B����J#���T�ĖX�\'oF�j+Á��H��dT|�R�:4{�]�S���J���� %�T��~ULG�J�u���˥>�"�6'$��ĵT����ʖ٧�J�Q��������CT�?-aC^e�e��t=V��=����'��i�׽����[=:�1!!UmΡ1��>��=�}���= ��{�q�KsIk�ԹB��xSE�o��q�sB(�3'f1]��J^	��1�򬃢\�-Y��RNacgh���U���jP���w���D$>|1.lw�]BH~���˭O G��e q��7r&�nە�� 4K�� KT��ȗ�u2���L�w'�>f��T�����.S[4��y�(A��OT���Ĝ�	�uj��g/��Sf: 
��+3� )��r�٠�� =�W-;���٪[��cuL��I�
��Я������L�_��W�ʉ�4��V�n~e"yZ������dS�&W�6��nV��q��0E��{-��gL@[~�C�n�N��H*ghc���P6K�r{�z�0_�Ƞ8Tj�M+W�Ad]8C~Aof�tp�a��ٝ�P�I��żME��w�3&!M��w����?! ^�,SO�	֓Z���`;��Ț�	���Tv$�'I��.G���x�o��� {ω5ڊ}��u����_�Jz��~�O��	F�u�qy՟�s��[^���I��a���C�6i%ċ��#l�H���lm����2˂� d����iZ�ar��x�o����M�C���b)j����7���w^^�/Z�!�%�ͪ��Z釧�KiD�q�;�&�Y�tc��{�#��u�9c�\�F	���|ܼ�(0�ƹ\̀����������A:"��58۞rڔu�"�����AEx������}0i\	��!�`_q,��310���'�S��^H�K�u1��η:��8��JP�\lV�tR$mB���po��a���ϸl>�3�����w�|�:���a29�P��0�­�dM��CX.��v��ꁭh�6��%�;u� ?>�H�f�TÎ�_�5&<^O�5Kў��~�U�OWtb�U��j�&'^!���@�N�h��D�
�!�����> ����[���"��N���V-J�s���k��%�~.2�¬�	꺼� �:�G�[�%�'%����B� e�~T~�V�VIQizx���$�?u�E�v	�MV�u�w��N�ˏ���1��m�B�r��/�n���N�Y�{mMz^�;�v�����U����޻�_����m�wAY���w���W�[U�;\<�3��CŒ
�/$��gx=b�yb�N$�2`�w��[\8w����Uă���'��{�0�7�0�jm�bFx��c�^�+�@?���,;�P��$�:Y�Wx�@]�=��m��𐠯3p���o��(���.�}��Y^��㌧�Xsv��@P��x<�d@���*�[,7,G*W��aA0�e�4�� ~�$�Q��D�����*<'�p\�p�����!K�+����y[{��6���-��I��{�6�\��I_��=��洙�|�q�ʹ�v6�G� j,����t�yЯ;����7ol�}� �\(İYP߇�;��h�/d�)4���uV��3���R#�[f�9%�3~�hl�
�m�0"2�b�lm�>�1$��co�v��5�B<��a�q��e�.��Ls���"�p2��v��/',�Zɔ��0ʵ��V��F_ӝo��u�R�7��+�y�=>5/�K�=�I��0h���q��B��G�S��쟒�l���I�Ţ��!����h�'nc�
���{s�K��sцy��X�,�m>�r�����2r�t��$Y-S�"��]lG-*4����p iߐ�$�QBu����t$Cmv@i����8'Ir�Crkc�%C,�eg?�;$Ҳ��KCQ����h�Lx�u4��#]S��-̲YIn���Ma�8���-k8W��/�BN�J.;M�!�B��u�������c�F�dT�/�Ҵa���;��Mư��)#�#��<tQw\���]�N/_���4o��߁`s��F?a�j���R����n<�ؕ��=����FhԿ���g��i阘�]���0/�\��o!�y��"��sK|ِU0#�:f6�2v�*J�']9����Ю�GYm�˛���md�]`��6�8�@:5R޲�ud�2�ڶ�Еs3���d�kp8������n��9<p�J�IT<p�v���"��~��"�B�����a`���#��eV��m�����*
�<��e�<�^p����H��>}�y�������H����*N�5ol?0��|}w��v8䃏Х��3���� O�q�#y޿HD��c���HA�V�n�|:� ���QF*=:]6��4x��|1ɬ�(��_��ř��㙪_i:J�	~�~����W])���ϥ#��[���ML�1���On���N�m|)�SK�����HU�%L�lRX��)z���6��w��1��0�|</dy8��1N�q���X���:R���3ў��4'b"nL���t�T��c)���-�X /b�c&�%�e�+\ũ������i��%�(�W��y����Vq М�eݧ�=J�S)��M�w��?a�8%���`;��$��힞8V=jx�N��?�ފ[�;��=!��<�IQ���V\@_.�r����p@�/[QwRo�t1^�~L�z.�W
h�\�G��>�Q�~M�0n���pfX��=@�>m�r֬�����:�)�^mg�P�,�#Ä���1N��3
�3����`!������48J��-����*}�=�y�kT��x��!+B�u�9Y�����М+��d��B&Ζʎ�&�A�uV�tB��ҩ����=	�j{Q$�]� Tˍ8��@i0<�d��4OQ����Wo⁜�|�������1��J�Vp�)
\9H3��U����wN
�AӢ �:⃚��%��/L�Ὁϳ-�'��0n��B�9�.��(k��D��� �D)վU�=E��ֽ~��k���=kp�+�e�2�/*� �f�ُgX�X`[B�>bNiWg�`u]����"�Ғk����ǯr䡝���z��"`1�FI�v�@��$�r�Ǭx��y/5~�)�R�X,�|���L~�B�1)W�/3$md*�
���xe���]	J:�f�§�/�(r�3��P��}��^I�����~W��G��so�59��zkS�q�6�cb�R�sټ7N�t�BB�-|��R-���g�u8�7�
�����&�V�-5�� l��t��V�7΂���~���u�'�5���fë����,^�%
7��\�(03�O���*�D��E�������vhm^�����%�ˮ�/b��W����U�
��Q�/?<��Ǹ�5m��LtVc��/"ĸЎ��|�=p�qa`�wLK��didA�a+�K6}�g�Ly���h��@���f�s����lG�� �ך�O�C��|�V��d�֞3�j������з]���_�	>�H�����L��S<l�o���T��m�G#�R�Ҏ��u�1�~��/J���R5��{W���� �7P��F�%�1|?��մU��J�)k$��
]�ƙ^�P���J'N��q�ji�>���>��ȸ���[�oj��8��<�F,=�1+�'b^��/�PX�K�G�+m�۹�d$�P�-�\~��&�����RxJV���n@���i�s~+���hRo��c�Nm%SO�>������Oibt���W�A�|�:�˸W�����ҐIb���\�
t{����+�a�Ϸ�=e�����~�H�,;���Eո�����C��Ix?Mvf��Z��8�#%O	����}�c�p�kf������<��g(�p�e�R��]-¾��!U�|6j�p�U����|fJ!��>��0�⥘���J���o����,�f�x�>�r��b'<���9�R[N3EV��o�z�)@N/0�m
��3R�(�Z��,�8���X7���Ҭ�5���n�a\�2\�d��������c"��)����	KO "n2����1���Q�4�Fi�7��-�%���(ǒ;����|�栮�@�%=KG��Nޏ�0m?��M��F�Zl�U�+�2��,�N4�p���	i�&���}̍5A�B����	d1>��>"O{.���р��j�GO!?Y��B�hw�z��uKױ�Lɗ�r�k�������D2����$bA��@�_&�>V���=+@��w�z`T%�0�0,�E�P���sF�p�h��֥`�V�����4-w,l�FMG����Z�X��rcjl��z��Yp!�9���Y�kϨ����'�?�2�1��>]n�[*NF���;�5�&b�C'2�>�t�?8v���e�Ng�,���ga�R���=!�,��T��N��2�]��X�0�8�4��<�P�2U�2��B"����}l�g��'������`��;o_P�Y]�܈������A�E��*�`�}f	��i�[;E�(@�ɂ" �����L��~��za�i/�9�SD���3���k0Q芋�N��v\��8%����z�,Z(Y5��/˪�Z���|��E���ةN��%�Yd����H��iO�|��� b*a�$�=�d����R+PfNj�[w5�����|~3 >�� ��K�s���!�T�o����a�d�e�`��BK���6��#�`��3���F;����b!/�b�Oœ��i�cq��"��"Xly1ҫ���pF;��Izq� z��'X�������Ӹ!�����K�4Z����w'F�k����Y���*B�sx�W��ӑ���.���	���#��.۰V r���pX��^d���uTJN�t�C�ؖm�8� �'�IK�M1)+,p2��v"���0\ux��.�53��p&˲!{l�(��Q.~��Tv�r�;ҷ-N8�
�΢���� ��8M�C+yt��k3#��cu�}R��K3��
qӟ�&sݮ2ȞZ�d���w� 5�Lh��� �q#^����.q��[	Gβ{WG��}L�%�=�A����;��aN�w� :e�8��]�qog�����K����� ߎG���n�����k�5z�A�PE���մ͙��b��hiĶ ʺc�}��c����쁉B��f�FCQ&�${�S�1�ۏ��\�>��P����]q�`����'hd��
��SĞ�����f�����,�{��p:�@�N�i�e;E����'�ɐ�����Z&��"8����1�o���_r|��J�PV'@�J��F�+:0:?-5�C�b�hC��>�2���2ڰ��Qsnq�ʷ9]6�B�0`sj�_y_�.�$+}�G�����4aH�b��'�gPi�ζ�q�$8�-����*��_��ኲA�cm��t�C+>���ƈ8�E�c�K�9�'��"��9Dnv��D�\i��2�v��<��*�����Åz���;X�{{���_6J;��o����W��P��(+`/8<;A��~@pv����5tP��r=�d��<��^ۼA�+=G��I�0���Gtn��!BS�!!>d�ӗ��PJ�2��(��"��j4Qr�����u���-&
����F�I����U�B&Q��D�bW�5I��4��>|a;@Z�O�I�q;F��U�F�A�"�k�7���a�0���������c�.?+ ��}�'Asҋ��kA�64�R=�]u�;��:�)��mEP[���o�-�c��r���g�	z�������<v����׃TZ�x��>R���L6��JA�?�
D�čM(6�~rˊ�<dΊ�JOL.�y�W�gy�7����S}1ZZ��Z���Ixi4.@�����VhF��� �)hxr6��^]g�l�i���+hI�H���sb�e:�ǁ��Y�����_^8�;1ξ(��+)
�IB�V��Ӵ}��=*��'�UU�#q6�C�i.p��+�����u�6�j���~���Y�nxN�u�.�4�E��3���w���%#�^ϮLs�e�,�����'%���T/e<��T"&_�ոq�CJ1ySr��
���Y�����%5J@��W"��%@�C�bD5�6�SB_s��� �@�Q����M���X���$�FF�p��#�e����Q�C��$�8�h����� J��CuUʞ�5�B1���s���,����9X����Ðy���%�xl�(�k��x��]�;6B����"+F��b�~�lz|�AvcX��{W��,�k�'HJq�A&�D��!U��W�T=6�ld�.з�j�C�":~=E.�_ ���r�Uĝ^��
���
Uߧ(��A�'�sESs
$:Rۑ�]����L�΀���(*�.'-!�J:[�pqo2� �B-��l��v��|�+}�
B ���]͛�-x�&%D2�M��t�c��w�O	�Q�0�ȈZ���
3�8m݂a��Ǚ�^�4�ݞ�ރ.b���!U�W��s����`�\�=�nS�Er��>�i�==�4���{����t�_DņĤ�?L6��img�r���@'�=^�S�tc�㾅7���\���g�����h�!�q|��������Ĥ�)g$I���d��c-o	�V�Y@WZ���^.�IL���?;�=�g��Х�B{�6�呎	*B*z%�i0p���b��s�`��rk��ӝ_&�B�s�gIGi�����u����;g���R�,j(9Gx��$�����~���5%$_C
��H���wn�(i`�e�� ?�C��E�䆛i�@yF�ρ]�O�W&���E�"ɵ����	q�nH�̂��R�7�KK�۾�