��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>����w,.��n�Pm�kN���5(�=-R4�(�y4D�i}���kEʴ�D�Q��ʹO�t���^~M���.�^0��GR�wRG}kB���� ��w3�V���,���i��x/��[�f8	�=q���tM@2Ҷ	��5�P�(����\���Z�%��*z�	�h�aq^v����7����틻�c��bCc�Gm*��r�i���l��aQ3<u��K��]�Ml��Lh�#ԇ1ޔn�N��XUN����>�s!�+f����g��P��把űa(p��iF'(΄W�q�T�t��h��p�N|�qӶ�>-����{��b�kȄO�����Y�X���w�����=��㞡>yU�6ݝ���2�]fm�^��-2tO�`��~B����i[�~�F�T�@�%�����3���=���x�</�
h������*N�����p��oG���P����د���t4˨�:qUc��ʷ͠gv�}B"�X��Cj=Yru|�ɜ�X\�i2:��e^��6�c�µ͋��a?�:?��j���a��Y%$A>N�#����ClY�<S���g�"���Nq��nH�Th����`EK�aJ�YQ��m��T�S5���T
��v�[�6�/b"���QL����l��Cr�L�'��Q͕�w�!'��ǋ�s�Չt]��Q�5Vѹ�BHL����썡x��
�Pa1\C�ĳb�ROR+�ּo���ZS�k���_�w� �>8O݉�Z�l�N)�Ș�̝xH��r+09y�� ��S+�=m��y��m[Sϫ��:%'AS�x�;�Jv0�*VK�?PěW�T{Y5U�h$R����Q��@��hk'��G�Ğ�A��e����/����*J�nVll���!�Cf�u��&ܧUDO9V��{e�)�L+E�#��0��[w������ĭ{�H�
Э�E�9=j{2M?�jV)u)Z�D[����S�F�U@AƾM����ʿ~0�!��Ȕ&7�/6�)h��(�(� ��J��	Ԙ�S2��՛�ڊ�T��b}�M�,/9�[�T�j4=�x�^+�Jp$��<�
��Ӏ�
f=<�6��F5t��~N��59Fx}o�ղO���V�[�"����us�G1��u�8����c�~�˪D-�9?]c����Ȇѹ�8����Zn��V	X��0���
��s��Rӛ�e1-h|���jT4n�KLқ5$X�2B2�$	 �>U�	5h*Ј
�ZGل�C-�X�����2���t�y���i 6�8(Z[�N�Mv,_2��ҙ��p9�~���d�#�/��Q�P��@B�"�
���k������=�3��1-`�(��*��c�fY�Lg.��@Iw�����KO�7-��Un��X��R�(5O��?�����f�����
��2�lcS3��s!=����'��~�ʙ[�����] ��T�R,y�\�_�$���_K���2VҳAld��R��QW
�&�Oc�ze8O�͊)9ҟ�B��_��t�M��83��U�t�Y�*ԫ���h�6������.�2�;*�E�2�nP�� @��7FԬ�1�Sa��F#����Y9;�.��Ӗ��0t[������4(K�g^��| ��s�]��;8���:�w�C�RL2!���a��6��8sı����8��zC��B�A�sq���Y����cK�.���i|@;�nH��p-ET��.+�����V��U��h�M��W�{����P���]���/�Ԋ��nH|9��}��q���Z �� p@�/�W\�>K�*Q��^�<��w}H�eA3�Lp:�����>��م_f�#Yl�Y1�d�Q�d��o�LQ9�q$�!��
�@H��3"� �,���ax�#\mvg0���B��~���ip.x��J�^��f�	7s�g+�-��3'(�*�\a�ڊ_C��[?�V1��4uj�+�MiLYaF�����iM�}�d�Kf!J� �W!k�c�"��H�n�y30�tU���`.M{��(^�T˧ُƵ��[�z��-��IBe����k{��Q�p{���8���!h��uS./�S�.��|^.�Yj<;�Kw|X$#5�r*���n��'�p�C���Aj���1�k�N���zf+)Ad~8��{�Je���Y��BS~�T�J���h�V,���Ց��4%��Xx��QZ=���
�0W,���E��&Gmj6&br[�	-c�H+5��R�@��_l�Hpr����O�7���n/�Ń�~E�X(X?�_TV�9�Q�n��+ �c���0���B���p���i�_~�y|]���~O���W��R<�G�Wb����i"^�����rX�`2�l�e�_0cf�Eoӿ�,*�!I�[4��SܡD�f�Bu{�MF.�#H�`7�l>r�1Cu�Z���Iޥ�
٨�{jtaZ�Ź�>v/׮��T'�"yh�E�
�V�%A�}ѿT��_*RjU���-95
����[�HZ��HT��(L�F�/�+ǵ���k�/�k!EP{6n�Z��bi�ul�i��s��]4�}"���u���5w��{�ͳ��B|�Ͻ�8��jЫ$��O\�8��55��[��\���7"��*�h-�8����p�p��~��kEƃ���W<"�Py������˅d�~�udY��j������^�v`n�2f��[��%+)������,�7O[!����|�G�?��U|�I�g'�=�������fo�x�Ƞ 5�"3/�D|+H�*�X&��I|�I�ӈM��׊Qk!����w��qc���ˤA,,�����I���<{�o�W52�h^N��_Z�m���,_7��ξ�N�}Zh�_������!pXu=q���'Ee|�K���_F�N�B>z�	�Q yq_��Q|�>X�U;MC������H�CtI��B�{'��� ����8�#u��Z�y��
�W֪���O�a$�ٱ�Q8 `�ܲgR'y4��.����.J�����t�r�Q|e?\�F����g�'X�l���ͼ�Bd�(�+��G�=�B�7��S����Y���@�+Cu��s���4(�����)'����������� �c��o�\be�F�V͉ ��U���6LJ*�cF������KTx��s6��49C4���;+�jҵ�YT�%�,uh"�g����p���Q?��Ep����f������yE�U���YzI�*nT�QB�ގ��68Y��io��\>��Z}��5�8˚����%��q�`6�'�삭�ı�tB�57�Q��i�6��|G�ۧK���X�Т����������dep��J�����HVi�@Q�����2X��%���5�D�-UW$�3Ѳ5C�Dd��	(�̀kaKv,�E�l����춨NX������9�t%~"N�9:ކN��.���4�&��7�<������-�S%z�������N����.
��M����0`��z:_M���u�1p���6m��)@tA��s��Ħuc�,f2LMM�N�@��t��"!�b|��٣��oݤ�w�GP�Ad��E��C䛖���gI������L'�s[H���p��ݡ�U�5�~���]�|�T7N��A���~�Q4����vn莍 ��1�J�j��E�zZd�-^C4c���se����I=��>� �~�E�b�T�ˋ�M!x��c�����-(��{�
�|Oc�J#7lF��1�ώ�T�H���B$���{K�fK>���J�v�d�ʨL��è�@��6��7�^"fMY������}��*�[�i!㖔Ne� ������2�<	������'��*��<Y�b���f��R�Ö���N��n��h�H 
���C���q��G(����K�5�I&Dݥ�w���&\\Gw��m9N&�$�9K1�5��8{�/�f����ݯRts4�Ȳw�H���#L�q[�)���Z����q'e�U0$uM�����hoq8�>TyF @�E��������AxG�i����z�_���q+o�7 $�\^ �*�Q
#"*Xqփ�~5.Є�}��W�^nS4{>�Jحl�.����� :^9�(���0���,��E��8��<�病Cۡ�؃�^S���_����=mS�8^mrL� )W�~{��4�kG�A4�	�=Rl#�K�R�