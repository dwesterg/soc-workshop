��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t�ă�T��i�W����%+��;�K	��n�{��y��k x�Sjǥ[=�?G_�Α�b\�m˨��8��:� 87_]�9%��zf��8u:����.�Y�\g��jZ��0�T{~4���3n���#k���0�ߍ"7yO��kdk36>O$f�����e*{\��Y����0jx4���ē\�/;�>��294��Z�5d�����~3w<�^8�d�y��;��D�Ԕ�I�Wh�b�j��`X���� e��,X�[�º��"���lQ����v\�Q7e��1}��'�!5�Nm`u09�8�lC�#3����nm��MQ��g,��J�neI�7��Pr���R�42V�ݶH^pkw'Rƅ�쟾 �TEyӄ����������-�}�p�=d�}�vR��y"�f��%���k��Ckz/��6��%Z)��tgo�Y����A��;+m ��&�	��2Ar@�0>m������:ԛv{a���#�:�hmR����޼��3�7ձZ��cr�A8�^S��ѩGx�nۼJ��:Ϸ;MU��ld��T��_�W2������ߝ�&�:jc?x0Y�ۉ(�[��;�~u�@G�[�@�e��5u���R醐`iv���)�5���ىl6�ɦ}ƅ�X:M��,w��Q��r	��G���?l�P�B$�~��f��T`3�1��Q��ɹ��u9*����j�Z�(jq������ʣR"�D�u��hՀ��6��Ŵ�<��EH���¢�6
�ԧ�g'�A�=a�+N� ,��MJ����!�r��wh_�6�NVN��9��N��õJb�?"��������UM]�>6O
SS�i�_ O���o��>���=�/,m��4�� ��1?Q�_i"G�Na7}���i�MY��Oכn�a4]��J�w*�)���`�\��]c�X3&��0ٯ�8;,��RA�z�t�Y����m�Ou8�����m�@��0��E�7�}� ֭��B"�����i�ɔȑPK�mJf�����Dac&0�k�d��ikԓ�-6��Lk	��Y��5���ő҅���(��gI!I�Tr�t[�</� ��~�		,Pƕ	�-IN�Adׇl8��f8�B��?B�g�KV}:1 �0r���^�09�5��
OQа7�f�t�2���+��WN�*e"xx�y�+��XJe�2����#Z�զ*� ;����04޻��IH�@�ºUx�fE�pyۗc�4z�ϐP?r�0���{�0C���[[Z��Z���̹,��������'�����];0�l:N@.�����p����K�qT+Ⱦ��~�d����|q��|�w�n}fެu�j���b��Vne�S������1����q^��݁.o�a�Qk�W�O+Y�ɱwH�K��n�I��"|�:h�����i����|z�U���
����O��~�k�$P���Sd4|���#��w��T�~P�ڪ� �Jxt�3ށOp/�A����,�g�����5?��8m%]�����_L��lVg�n�3.�À��Bbp'f�.�I�����N1� 0�n7�D�ϳ��i�-� V/%?�b�������U�7�]���>�i�EgN*e�k2�����V����� ��T��9ª�;dw��ֆ�z�Ta<Ø`������9'hR��~�JgjL�����鴍rh�m���{7��'-�a ���\����N���xp��f�$�+�!K2��deǫP��WK��ᬦ�p���)q��?����u���wH������P�����ˣ*7�m���mE�g��vi���*�	1�4\�S��d��&�M�x$'�X��	{�qD.GB�vl�+f�}�B+�L��@�A��N���q�-x���@��C��S�ܦ�����`ߞ~MQ9��V�&N^_�l�OG�m�p���P�e��2��8� ��=���?��U�x�cS��P���CťHǃ︻�*˶� ����Z�t�U�(���l��jm�qL8��歑 /�}`�T%�0�tgM!3G,z{�e�h niU �>�K���m�Rݳ�	������R|��mʷ��;r��^��I؂�W����TS�Y�"mv���g.bEj`�`�n�?�*�9�� �AE"H)zR6�I��U�ԇ`&i���N�܆��v �D�,��E	L�z�	H��s��\��5~��
V�N�B����޽�F�,#������
��J׹����$$�T��lR�+�\�ΧDxR�t%����*ļ�Ẏ��n��B��)��FZL�e���-���M��D��{�ˏ���-�j<�D����������i_P��I.3��N�K��Y�Vg�Å�Z�%ޓ�!K=s�Ѕ�#No�U�r���%��o~j�i�ɔN#�+]��20�u�/�b��[{�;|��X�`¬a ����7�m0\��+���Z�\!ا���sX͋x�[�rHp:�`ϸ_#���|#��7%E��=EHV�ci2�<�dA���R&4)�hN�$�����j2M��p�R�O�2*�X9�>�sw�I\m�Ը��l�	�DT{��;�/_Q�&�/��a��?�,����q%���Ö:�[7����^��v�pک�5M���4�c6U�v`�KC�$L0R��S���ک#���W�.O��I��n���۷��~���B�J�mt�};�А�P���rJ��n�Ğ���>z�p(��
Ј�+���ɽ�l0.s�aڻ82~*`F�$�������*p=�1��L���_�0���{�����b�v���x�I� 9�M��.DC��8_P����;����oG�Ԋ�U�dK
�3*I[>Ǽzj7J��yia��'�aۭ�_��.q�(7��X<|��Xu���B/����#�2��"�m�I���$
�A4_'�'�V7Z/D����Ģ�R�)�ҕci�a�7�^�T8.��F�s�Ҭ�
F��2د�н�j��Vg��sY����"pv���}�����r�(#
z��%�:�:�r_�?^�e�d�4X�~re[yf�fL���A�܉&	Uoe���z+w	?ﰫ�C�1t�>��J3V�e�r�f��Rթ�v���K�u�n�׻�	9*�W�%$IN�$,��+���H�Rq>��Q~��R�2ƚ���×,]���c�US8�'#��"��U�3%�?���xD�:�^ ��l�I'�=������A�^�S����Ӳ֣,��O�9�EnM�ۄ�#Ċ�.#�[m���8.=�Ԉ~�8a����5����V�,�Z�qٻ}�H�r��OgǠKt�$��&�
wH�J�iL�"I�X��B�I�M����jv���VGI��y%Z�0��u�9-Fobo,�հ0�(S��z+�?�\Σ�v�T�("��#����>\�� Pc���P�8���.�5��(hP �?��N�[<��;�� 􋫊�b�%F%��Xs�I�ě�0�r!�1zd�*�N���+�\�`}-�>~i�-�{S�m?���T��\�8�~_��F��;"��?vv>�$&vEdS,E���IR��۰3��
60@`����M[��ĩ릯Z�EP���%���2������?;����S�M@��:����_���krd� 5����4���k
̇�RܬW��ZD83�2Gڬ��u���\M(g��M�	5�Tx�{��\���|�Y����s���!`)�p�:m�Ι��bZTш�fU<�;�����>i�T�ߌ�ҭ̚�uAmNI��cu�W���k��"?�w� P5Y*;C��oO��Ol�Ć�0o�1����H�\E={ 5�¯U�'J�m���q�N
a�������o��ݡ9�:�"����4��d.U����g�j�%����S��L��1�֏۴�1��za�^Z�N�V��^M��x�1�J�O-��	O�p�_ BJ5���k�����wl��dsd\�>
�[�P���(�Z(�X��ёN���^�1nk�;ǳz�e��5�v�'�TF�p;�j7���ʣnX+���S.2�'w��m�EMĞ\�XÕ���\Cq|�cL9���%�>�I�`'C-�ʞ%��j���͒�Fg�O�1s�
��ЪL�M��`�`q)R��������?j+T1:�ӫDd�h�/���ϕY����,�;�h���'��	����2��t�q)�=k=\AT7�*�\��5?���
����)�Ĩax�����گV�ڞ�ͷ��kj��(��O� ��#����8�Zi+L��'�ZIx���p�B�9���C��i�t�ʻ����5�)�}˭��ԧ���c�.�ԧ�����,�* �c���5�e��ä�n{Tۤs���J����<m���n�cSvE8}4q�z��.${QK�N�
2Se�3��R���TJ{?������0�����E+�M/�����kB���a7;��9��7�}���[i~$OzF�x+"5���`��zi�4��G]�H��:&�e~���_:������M���V���au����_'�\��0�J�2�i�܎�2/��j<o/4���tU�v9��ZO���Pķj^��̇N�L(\u�#0��TE� ��&+.�8�ް�����(R�eD�:@UR��28I��rb7,�Kk,AU���=����Bk����d	's�3���?�[Cgߌf�4�ǆK�{xџk���@�RV��8˴�*���`��;�;E%�8>d~�b)4�� E�&�g���[���c�� �H�n��]x��߸a)��Ct@����(@�ZS����jޮ��IԱc�+i���h�$��0�0~���Z��R'^�*���F���E 䧲j��D��mK�;v�S���ftƉ7�7!����UW�0n�,��!8��R_�����g�5�P\�
V��\�$�m&������ZJ%�nӱ2�-�X�B}wC�(�rh��8�O^S
|���}��)N�~���x>��=*��ށ�>7�|=Nn(t�H�<��`�7��-��5S��O�~��id`��L
,f'S��5�y,��Z�m#����v��@-%P����Q��G�઎2��ze@�b&�IՄH��0��g,Η@��������c��4急�?�IS���_��τ`��&�<�	�+�W�M#~[AJ=p?4q)���2]?� 2'�,'�Jcb�N/D�xS����|��s;�\3��s��r�`��8h��ȥ^�&���֗<�ؿ�š��#��o�L�^Y�2*b��U�D�(`f��3:��]�}��(�}��<fm�AQ���	��3Rua���Y�Tj}��nM_ ��.R)C_��)����rRB�٦ԫp~�*9�htI�t֝���!BI�Ev<�����@��%stP8��y�Ů�bDG��������v���%2�Լl��R?�z0	����ܰL;�XN�2����]��yyo��!����ǫ$�p: ���Xs9iZ�L#4a���0J��'�,8�AZ(�4�F\���,���uIS|k��*N�mlT�ˇL��K����3�)k3J+(�B<ɶf���c��`<�m�dϳu�'�ӂ�K�a��≢�>\��	OW�e��K�D���1s�ܢP�&>�&�"�Tp9H�Os�U����ƵA\�-����[����$v����{�y h�nz�E5���=iT�A��֮��e������IGUI3�uʬمq���!<��d��v�i]�Sy�N�I��r#1�� `�}ƆBr�ɿ��U�f���h'�G�τ���t!M���q�NC��,:L"����xzG
�k��+0�9���Q���ك�=2B�~V�n��##����+�0��^�~�3��h�!�.etv2��1�v�}����5������$�߉�	�@�d��n͡]FJ��褟�ea,�>}R[d���{F�������V��%"F�W����zD亏��*j�r˚��u(�p�H�|����_ԋںG����V^'9��s�h?[Q�����e-4�|����U���%�����@+�ѕ����Y�v�ù!�fK�I'~ˆ,CM� ��F'���?��=�%6g���i��,O�3�j+�by7ؓ��`��a�� ����ߍz�nֱW��r���;�{���l=�Dp��ۊ�VIRd�3�ŕ23���Yz��r�C�Y�6�JI�$���f��ڿ�¶��sRv�,z{��+)L�yde����
}*K��]���M�m�Asó�f_��I%�r��!�΍���Ϧ.���!E�P�AgS!"���cf+��ל�-AG	������LQ��n��:`�y�Y~9z���5�F;�	#�Χ/���Ɍ�G=�~�"�����lq63��B�@nc/������z��������=�����7yt*�K�6a]E���i_����o��oPW�Y��s�J�f�^]H�����g�E��NIm��Q�d3�p�Tb?�a����:���6�#�t�p���I���;�]*^R���2X5�$y�.Q���j���TQkG�jm:�1���6��u4%�x�*��Ew7�7�PA�ۿ�Opڇ��A`-����h��x1&�@��R׸v3�"�U�'�%)oh��[�������]�!9 �����u�z��F�_�uG�>��Cf���R�n�	��.5>��p:��(έ�y�'*�l�iզ����!�IϜ�^E�H��6�g=�q�	xW���]��i��3e&x��o�<�u�5=��4���L�����j��
��M��Y�'kM}��]z*��3�.J"`��
,���9k�/�����׉���
��/�m,\۳��z��x-;�m7_Z'Q��p�s�_ Nڛ�y�h�V��@/C���a�����T���+|�L݅	�oS��9�98-��� �FkX��>�J�"2_�}6��
|�;�}��D�Y�X&�|8-��w��M�U4������	�;f�L�u�×	�3���G��l�fj��ݼ:�Q�&���uudp�@����?�5� M4a����e�J�ɗ7�'�O����<�h��tA�O�]Y^ar7w�g�a� ��O�b#<*M��B�&o��"HT��-OE�Ocq�Ev+�:�Vd�vA��-X��_|Ae��GY�\�N�#����`��dc7q��"�|�>ȼ� ��|�N8d���-�w��D�lU�mÕ��m(�4m��B����&�tzhs�m}���L'���Ԙ�!k�(ͫ�����W�|y��J`TTv�i���UX�(B��2�|qu��eJ���ɜ{'̞U�A����T-:Y@h�R��r�W��j��K��	-����S�c~95��&w�.'B�?��s!��o���9����O�~i�pq*��W&||hN9�Bu5
Xz�X
+j�<��kt0�
�*\����W��u�������j*�K�:S���4h�Z�[*���eh���t�8�Y�eۉ{H��_/|p�՞�(���եa�I�i
�+����`h�q
(?�?;%뤚�Ֆ��#��	Tޏ�� �]�L�^�x#$�5���	�8�.�����
�l�%)�c�^@r���4s���/>`u#+�_���_�e7⳺�o��f��|U{��lɳ�E>���L)����Ұ��?i%%�H&9MHGt$\�K`Y7�8N�塥��悡\����V`���v!�S���ѕ<q�'��� pP�e�l=qk��9$�p]D\�;�7�+SO��烧��RԻ�G�sv(P�б(E�����hҾ���y��Z/��3�+�1g���-�l�wM��#C�b����?Ll=��Ǩ��bB3���GTޥ/���'`�$�T��3$�PH�W�7��oON�z� 
�����6��|���1q� �_��i�����'I^�`v���/�9o¿;�D�i�����<J=}5(��u�A�º�4z|ŵ�3cL�|�-R�Qs��ҼB�&�M�w� &7K�Y��Q-���6�u���t8�΀3`G\�}���u}�p*��`��q#e����&{�p����d��"��4�K�>����c>6G�i
��B2��4��d�0�Ʉ�]�?��P՞�~�JU��[�'�B�&���u*š��J5u9��
Z����\�����{/͙%*���᠗ˣG�GV7vIxM1�/J'u�/�R���������Q+�0!4�����nu��]F�����K�d"&�K}������a����F��z�=�v�C��ݖ��jw��Q!!���H&��v�9��>�86�+���%�m ���fzA�R�ʻ��1��� �+_��	�].�&y@��e���·�<��Z%��7���e�U�G��������#��$s�]hu�����kE�L�~�P�ț�~�97B�-�QɨM�����y	�5��M��ȓ\��Ps�Pϐ)����d�m�P��}i i]�u����}x�
�$1ĉ�
D��o�x���4FpԵ[c����A�p��˺��"�p�Cr���:���<3v��ʽW�+����Gϵq�`��"e��&X�$;�-׿��x����h'6�y�߻��C������ݎּ�(�kQ�&m�	�0~e�q9�L������߮�hvW:���j�ai�ʯ�F		�>��Аk�@5f�$�/	��W��v�@�����vt�|~J�5@qmP�x�'�P�Bnpb-I����V9�0�Hs��O��p�:R�Sh�Zi���v3]���$����N��|0�c��u�ӟ��ƭ�U���wf��?���.F�Ց͖k�qs�d�m��*t
�lMI>/�C]��J?>��{���K�!����
������{��T?����$ͻ��RʱŊ7��W��������h�%��QN�����|@�L��.����rD�K�熞O��9������7��+�l��C)G-�
DA_�i&�K������(7�`I0�7�Lt�~�l��M(�K̆��[�>�O�����y ʝim?[����R�Jgc?���"ܵ�v�+mEzTW��p���橽K}��)��� O�Qɘ7 m��Y�q0�ߘ���q�6U�FZ1)�	g$ҮT���-tAD==�nv[��5�$�ќT���)��R70u�g{��Uϝ�P�]ntFau+�8����dH�˟�~Z��[FJA����5��س���*��R�����'\��z,l=$���U0�W@1�⁉k������0��RHs��	EZ�H�.�ڥ�ήn���#���QuG������7^��h���yw���M��;���r��gD)���J��}���U��q9ċ5��u��}�u$7+?�u������ո��:;�)�.yM�US��`�{J�	G����b�%4�J�xY�&U��m�A!��{mi�����,��u5h_Uߛ֮�Ku�H3���5�SB�:�L�"&T o٤��ԦX:�����j�m~�K� \Se�DĬ�+z���,��?�P,m'�vrG�����d��g�����֎�	I��m`��������Jo�!��wt�z�yU������i�ǧ#Ր��,�ǹ�I��@Q�\�ln�_��r��G��	��>غ�,3)�Ω�T�0}����)�I�ph�OV�c��z0�{i;|P��
:K7�]�ƍ_�n
�����u턕m�f�E���n�\�V�gv�I"ĵ2��|��Fbث����[�5`���Y��Dm���:]���Y���4���E��h�]W߼��uO��Q��?��z������=��*Y@�K�������T}��?�jb�4�@6]c��c��s\��$wGãD�r�~E@����;���Ք�ͧ�2�������H6x���o
�7 �^S!օ��{�V<�-�R���1|�ԷWh�G֨��0_V�����tA6'Y���"`J�l�����Y�����-�|��:��YV���s���+<qަ ��SՒ<S&GZgU�8n���Dlk����
�%��.��ײW��,��Ѭ�}w�)i��"��!K�ޔ���:J�y�n�^��T�Y�L�7 3/����%+Y�攼Psau P��*DOE�/-�V�=��/�����pΰ̖��@��K=MW�q�Ϲ��;F�|7�����U?8�I�oBb�t���U���_A�����A�b�;�

���V�:��}b�����KlQv�QMڴ��ڱ��d���x���*�%\/���L�KI1��会��^�ҟc3�^Q�7��?К��As�5#m�2䵢�A?�^�
^�y)�.Z���x�X�ҩsVFQȄ�|��O�s���÷2�15ts��ֱ��S������8�lV0I�
����;S@�Ghs@�2�]ֆ�:H=�î�L�]�R��U�`q�x�0� ����&�!����a�G�3�Gq��2����)N>&�P;(r��yqN&���69���&E;4>���Cw~�^2�}�J�D�#/+�-�4��;��r�$�<k��*S���.��K�L�%�V��0��s��h���5z�Bi�_(=�6ڗl�^�&��RW(J7�˘`[
s߶�)n,(AbG�k`�͒��4�S�Ń��oO��r�\���{"}����>o��X�de�/����]=���}�9��\�df��$<�������vn�~+D�+�X�Ul�ǃ9v�b�a��3�w�OK*�Ar����9)5�9;+��2�q�U���c��ٍ�s2u�����MZ�k@�C-^�۽��?iR�9�J}-���d&*�TK!�C��W��S�6�����ʃ@��q^��M��y���hC�gwt4Z,	�K����S�O.$q�A�jm�?�rȣ3Aע�\ ²�Y>��q|�T�7a�t l�Ff�G�_{P�yq��Y$���d�-0;*���GqD�m%�ʮ���k>��.�@�^P5� �:�S��|�j��ў�q��=r3��0�k���A�ц��ё3#��U�����������ф8�`wu6[�:��;8�'�ʇ�H�)��
���6�|�>�ώ�1n8��W�LC$�P��!90q�\
�A�a��=���>�2��F���Ũ��Y��ᬳ/=��B�|:���q�ѕ�S�:Uwp��붃�hn'��Q�q3~:�.R��� C(��U.�b�(#�	��aALI�U��n:�[ �eY#v�g�;'�j�C����/��Sz��� �B�)4�d!��,��[j�듇����E�|�qY!����n���� ���*�%���o�=Z�bp�8o8Z9�y�G�tſ�4=3)�"����D;�7�Q���:5�G��𔺹/_�K��L!�@xR�~�+h�2g��>Gq?�-ϋ.���a�D��lm-Ż?��� 2��:7�{n�(V�.�/d}`˗����[��=�9h5��v�W�,2��j1<2	5[aO��2WZrQ`U���	����	U؝��2��΋e��
W�ߡh�$M!�H�NB�'�ab�?�"�R��8��X
�C�<v�6O�Z"�O��-.�\�g8Ct�{�/��C��B�·~�e��ջ�M���0A���Bpo��G�l,��W誆�.r����o�DE���I�
��J�=��3#�[��Q���f$�m5��_��d�<֘�X�2!��o�����\��|��1փ;��٠^|������I�[Uj�/Փ��)�A����l��hV|�Ң?�:ڻz/�m���O/�cz����D��a�b�ӕ(��R�h�Gp]F�����a�*d��@����<�|�2��%��Hp�S��UL"�k-V�)ӯ4���{`8���,�֏j�jF�Kn��R�or*���gp~�$bzv�&���em�;, +N*��ٕ"v���L�>��3�c��LK��t�[9@2>g!-<�B�G'��Wez��Z.+,�*R�������8'���%ֲ���A��	�w��4f��]t[��t�0����������/eU4�l�l�Y¦x��A�JJ� OHU��.!�zsu�(�\2_)#���`��s�J.Q~�=�VY�S>9�(����A�����eA��d@�8^}��ww�(�a`�-S�uR�q���8|K{�T���.1��ak�?��)C.ƽ_(��+�Rux��s��k��~��.�G�K�~�R��R������$eCVi8p�M����N53�0։G��-�רp�H��k]2o9cР���y�#�����i�@ƒN�)������2t���=�0s�'�Ss;�b
{��U8N:�HB��L��~'��'&8W%�1�vPu1?AU�^���7G��
�1�����f5iu����Pʑ������;<��t5�v0M&��¡��ֽ�W�H���N���X�7{��#Ux��Z�"䙭����2X1z���W��1��]y����D�n�\u�Tk\�]�:g�3�r%_
ȷ�V%�.R�IG:0P؁耲����*�����!ݹ��t܏m܌�a���7�R�R��{Q̼�D����,���f��!��!�8ѣ�k �w��'yq2\����h��2�f�tD���ԘKHx�47�m`K�fG$.{�j�s^��0h�t���ٴ�ގ��>j�7r�C��i3!g�y_�x�qp֚F&<09!��k��͂C�{�m�Q��gZ�16����|2�p�o ���;�Q:]'�����WF��4EIgI����!��Z��\7�뮯j5d�q�Js<�N.^\��k��cs������b����W@+P�� ����`��������&�\�Z:��Q洃�d/~{��[ELVrpPm�)�������"q�1�wԗg|C��w�����i(� 媾o��VV���ۙ4��� ����Q�2��p�ʀ7&=��f�%z�f�*����1Q1y�����r�/��s��xW�Һ��Q����EJ��[�d;�Q��D�@��!�@� �8��)`�<��Y�C�K]�J/\@c���gf���&ae'Z��<
���GBے��
� �O3�U�D���!��I��OA7�����9�Ʉ�%Jt�:z`�9�D�ɦS�����?.<���WG������TǍX%�|�H=h�}�[���3�Pѻٽ-�3�
x���v�=��{CX�si�M�%xxP���pN�����%�ڸ��Y�;�E�쥪�{Lc�[��aۼ�|xH�+�a�����3���iy�j:�L�/<�xg�hj�܆�<>�&��R��C�(sH1l��$M��'W��c?1D�`Ha��Ʀ"V�56��f~�lxXK4}&��\J����L�uOV3��1)Ū�"���t�8"��G����2q��pq*�g�u��P���BBZ0�oq�+�]���kn�W�lJ����O�0����$F�ɘ���y��փ7�FO�l"����p��$�<����*�h�ƶ��$}l���_Ws������J�c-7�C#�o	Ip����dy��r���D�k|�|:н5\��`*!`��8�#��ɑ�$���LwZ�n�F�����c6^~�P�ܕ�����4�8�4�L�Am�G��� d=�n.�����N6y�.��x,`�46�i6�H�"������$�TyK���;�g�+�C_��NWݒ��Dl���ȳ�Ϙ�c�������5�u�5=���
R�"��ɿ%�Ǧ��҉W�'b%�����f��C�mo�����)5^Y�1��)�4�.�&�q�dqJ9�%G��P[^CB���e1A���ةϲ�jh~]�v����6p���ds���`v�����Ԙ|K$�x���>*�4�*�
��j���(�<`��~�:U�� \�C�p&|V�c8�̧7�#	�:BW~�����z�V��_�řV�IdC�F��e?$���ȳ�>+�QJ��3+��aaj:���J�}��.��i"��������z�L
B�%-��>-?�̞��_����'/v�E�n�8�ÊE����{���2���测Dmx�lU.�Eo��1#;'�,�{:b�@�a����?>o�@=��F�Yo��m
�)�E��<��q���eZ�۬ae� � d�t�~J���AJ���#x��}�p��6�,%��#��dK��1V�do5`��G��綤�B!�]%zZ{.Zo�t�+_����}�XsN�".I�]��"�	��z,� �[��aX��~��X�:y9����/�����s���������lvK|� �����ki"ϝ��3��޶������G!.w�I�����0j���/TA��t[<�P]9�Y�O@V�W� ��L���	�%�w�\.�|=|C�ݮ�=h.���N�qֆ��j@U���?a^�ܦ���
J�*ԒS����Ew�:���u�ۥGi��^�<���D�*�Q[G�=�rD�E��$Z:a�d� (9�:0��k��z2��Fl[|P����� ��};G�c�p��]�y(򏈕���l�#d�j�N��bc!�1^���>g�0������W�� |��FHU��
hYudK�������
Ym|�ȥ2s4�i�e�4X��OC�*��+#W�~�c�[�2d��U���Zd���V�-����Z��{��KwI���ۄ�̅�юT$C|U䧴����zYs'�ɜ���rD(l^A����%�oTf�֝��������<��w���N�{�?M���iX�X���y}a�o�����A`͗���x��P�=�c��� ӀwDʺ�Rl�����\��<��:`x�����H�"Z�ШB)!D�c�fL�Aշm�/�=�T�_,��KMÂ��2���V�v#�z�b8-�K.���Al&�ճ�N$/��9���O�Y����b3	�gv����˗!bj��YH�6�	)�����N���̅�v
1zu;J����<�2�q�)ַ8�$��z-��N�I�pK����s��zk�� �!h�}���ӶҾg�N�����W\��pg���.�l}�͔*(��ӈ����:�`���q88�O`uIi��,Ǳ��yYMY���n+��޹��mBn��9�ٶ�,�+��k�|u$������Q������j��׹��0Z�u�UD����K$?w�ȅw�m-l;٤w�?V3�Z���K�Ô��o|��H��)X*�Th5�Ǳ2��Kύu�����$|���M(N"��^3Mԃ�3�j㪧�j��O�M8{.���k7X|:X"�8�7=�;@�R�\��6:Wj�����B
�)X�v���e{�c{����3�OI��_>B?=F\a���u���q"t �s��G�5��v���a ��:�r�F�Q���l�U�T�D�HK/w��T\��<���F�n�z�2O�������%f�� yUi�	vo�#@ ̝��6��Z��.IM�X�����v���i�H��7�Lr��<G��"�޼��O38���Cr(�C�d�okTx��Պ���*�3���w��`OV���w���V���0Ȋ`G(�$��Z tx�YE��h�K`���j��WȤ|˶��D��^H���Km�����2��	^��.�Շ��������H��bY@��(����y#�����-���5�T�0sg]0e�
��e�6���7ǘE)�Z�7���d�x�?����T�W�C���8�3f�b�y���?�U:c��ԺEd�L 
Ϻ]�d�,�c2D�T�R��iŞ�p��l���d&��D+�s��Y5̾���e��4�-`�-ƾ���	;���Z�<GWZ]���5_��@��v
m1�s�
�A�uϬ�P�	�zXUn��S�Z�H�Uc���Q�!Ɖ���_�Yc	{	��_>C	������#�e*�(����0�l�s�6�Nn��zW�n�d9�^�V~;;xʥ��xF<y�S9�qǫ���S�-�KYƚ.<��X	�G����pt�m�Æz]�M�
�x���
t�iw;�_U.��VG:���%�������\�C��/b�8���|d�D��ľ	6�u@P���x���s�B�\��y@�1��'l�?�oPj�qQ�0�;GF|�
�BP�Ȳ��՝��W\����Ťt�H�޵K�̶~�F�c�9�ig>y���6���l헩�K]Ln�2j?�~C�E�N@�$PP�����]�.c�|֧�NQ�����f��[��B�X�<�#C��=����ՐPی�r��@#!���5��gW@9ǲ/�u2�v�<�К��`�C�� �r��ߌ��4�)��6EK���΅��g�g��A��WJ�N����wbq�Y�1�U�}�ذ�����Ig_�:���3 �~��1a�g��S2Hl1�Y�̥>�@��3�
��i���^���>Ԛ鯌>Di�����,�Œr���0N΄�bߨ;�.�j�q$�7�*Dƈ���Q�Bv��8x\8�kk�z��=��������g��B��!�棾F1��о��.����xi����cO�����\���@�4�Tq��)?w�|55��L�e�*R�׉�K'�f]���+�����b ��>���	��uۄ�Ӕ����zk�w�ִc13òz ]`��qK��-�$���r��ꟾ�����b���Q�
����pP��w��Ŀe�4T_n�4b1�G���T���瓨dS=H%��#l��!}[�%�Z��PÎ�J�qK��復*}CqR�B�Eڅ���p��[p9m��<�\�%˔t�yC(��E�=9ڲ�Op^��|�����( Ǯ���T��T�g�z6bf�N����cWS��Zb ��s�jo�%Z����]�V_��Òo^Ec�ˁ/�0R�����[�����lW�)�k�5Y�(e
H��}<���!�/�>��2������}�Ktm�h�	;�9��A�+���[B�*%���ݢWC���]�vW}���pKg��5�l$#���l�'�u���ӏ���D|Nr� G�xP� �!���P��ӄ��A���ԍ5�촆�^��TU�̇7��=ny�g޴�H�IL�;�����`)w{|t�6T�o҂-&�&8���gR*8�� �}��������0�'������V��1Kt����:�i�`smXԑ����4����Y�%�>�^�yUvϊ�>%�T��Ny�t����hߔ�"�3&&ȳ����yN��:H�*�m�M�ć4�.�P�XԲ�ߨ��t(��qv;���=���G��Eķ �����++v�����/�z��*�����HQ@�P�M�I�Κ��lg��Id(ڋ��LF��X9�6�{r�\�����z����j�r�g�Ul��0\�uk���. ��c�E88f�>P<��!)	נ���3����)��/E×�}��!���p��&h�m��sQ�kl�)��3�1�Ǽv�����⡊��W�������
|��:�����h1�Ϋ�
/䷣��:[K��In��H�$�{e�L0ݬ��u���x�)��g��3����:٩��_.E����B����|sx�^檶'nH���rLք�
�q��j$;𶄺��-+��� b��r���u�:{m�_�	����i�w���}|��G ���V!]�E��_"T�6�K$9[ǉ?������>�b�� ��V#���c�P��Hf4�E�A���U{�8���	M�K£)W2Gk�6y��xM��q_�##=f^%����R/��ZV��j�{t�N� ������g�TpIg=�ӓ��x�+�ÃNԲf��\�� z����ޡ)������(27�W���Fr�>�G�+Y-eg�(l��`���x?H����g��\�v��1�x_$�
��lj��5��\�*�B4xM�YYFR�>~�����l��u�c���':�DK�wU�����b��e�vU{�Г�9�jn��Ő�����3b���	2�[�3�F���^�[b/��ֱ;0�G]#�c^%���������V$g
�q�Pm��P�W�M�3��EzG]��	_�p���!� ���:�~ލo�A~0dɪ�ϋ_9Ĝ�Wbi���]�Hn<�����X*���*R� �T0�)���:�ݖh�}�E�,��6��#+��%GN�r�P%$u�ߌ�қk})>������*Z���:r���&���^���`!�k�f�1�U�_Į{�����X:��68E9�)+��gp�h��V�� ��*�9Yp�<�
C�O�����D�<[�������b�{�B �E`���{]먫F�E҂[:5CP����Mr�H�j�9���j1�����t�5%�; ���SF������D;��7��_��w�x@ݿ��̃T�ʘ>��BR����aJ�m@�<1�N�_y%���uj��{������'���HO������g�|3�����N�O5(����T�e�����A��3��m��!m/G߮�t����
�?
�=�ۖ��l�o�`Q���l�	����X�A�^�5pc8��1���>���+��ϕYL�YoS�����c9�5k���(���9x��$�o��_(�K#4]�����` ��ggF����|��*�9�*��pH�p����4��tYkm�pī�
�:���棵ʡ��:3��1����!J��@z�$(��M��ak��ݷ{��h�*�V��n2��.���jj��������ER���#0='ǎ ��%��$t�ǁ�<#�;�]�ge�m�sqTj���Iw1��T��o&b���;��\ډ���kY�V�(C�����~
���kR�Fy�:&��]� �,&��"�(��{�TLn�<̧B³��4"U�[|���I��9�-|����?�!C�{�hm�Ag�����A�"Heu�o=&WIϾ�p�����aK���2�yO��v"B�����ᱚl#�KȺ�\�}&_V�Қ 3�BJ�g\Ms�0摏��i$9iKi踓���޻u�b�8CN����}�x\�5=I�)���姕"����]����<Է�:�|�o$p�l�8ue?��{R۟���]�5!6�[���lgA|��C�n�z��`�d�ѝ��?6It�8]�zh�-��Dz�������̮�@���6x��&��;���Kx�ݤ �'��U����t ɇ|҈˷eĄR���9�vc�{����ڂ�#�co�?p��gI����:��rL�| x@���o���D�gA�F�|� 󱒰��޽`��O�
E+BfR/BY��!h�P�QpQ�i��Z0Z�/��{b���*d��}�|��s�89i�L����*��!.���m���~���n�HͭnⰌt�v� eΊX�~C:t�4~j���*<R^�("�����<����&�hy.�f��z��WF�.�^ܕ��wI�vP��ۆU�c��rNs��������v�h����rU�����~OHz_Y���֍��&!5'�� cJݢv����h��a2ĥM4Q-�K��P�H�y�����c��QzpZ��&��qT?%8��<K32��}r3gw?��D�N��y�8��N1��7�I���?(�"�MF��'[,�#��2+mޙ�R����
�H�����U��L��(E%>t�(UY}T�*��X�\�ǂ.H�ԽwN��4�7z��xՉ
"�#`�#��KJMR��d釁U�L���!^NϹ>��8]�-\�-�/�([�b@B��?�=�>��Tn7�!Z� q���~b�~9�Bdd)ɳ/����ո�F7�)l�?:P��2�W���^+�(��H�!G�𤵊�t�r����4x�_B1g��9���T)��QY������96�'2y󓌽���4�ԇ�|}�<��3����Ѥ���v�-\c�L��\��_j�+k���)nq��d�՘u�̹�����h�6�#.|b���� �S-�3�K�Gd��k=mv��k�a��~�w�%�` v�r���T25��#�e�.l's��i��!G/��'�ӂA���;���6�������q�R+{J^��Z���/ʭ{x{D0+��h���x� ÛB���*a��;bǬJ{�S��xj���jF�:{u�6�ݳ�䦢e��/�'����m��v��K�	�P|[��C$@�A� Ɲ�R.)ˬ� �̟�̸��qݣ��� ![Щ�j�.D��ό��#�yS	O��(])�]k���BJ�(?3$�P�&"[��_��l����Y�x�n�r����$]�)̼����k�Ә�a/i���w�̔���^���/���RdO9�yKS�<jί�7�5���]t����~7�I]x�}��~8Re�9��+������m�1��eGl���yW��q�KH�coO�О.���\oՑ�O�%B]$�3�4O�c��X6�C[�.��:�Нhn�e&�~��"��Q����%-Y��ꓶ��%ƚ��zh�m6@D݌Ǳ3�� i0u�� u�1�F����%��a�<<�o��g����4h�'*I!����J��.׬��vN��>�!���Gz����x�TQy֜p\B��if��˄���V���#�@�'sC��ƽ�f:�	�0������
�CVq�o���F�fL�oV׶�v��DU9���� ���W�@�c�0�+-���"���7�]�%��q5x�N�S9>����JQYY�jh �h	p&H����پ3�l8*P*X'�_�3}�����)�D�q!*b�s=���
��4��iL�3Z1�s
z^�M �&O|҃|����,W"n7�&�S ��� �G�_6	��#Nn>s� ��5-��^���CX��/^���~g���Y�aX���F�'�Pe�=p��D�~/�cH���Gx��c��/�+��|$��s��7����r��$�����lbk�-?U�Ky�6��_�Dc��x�/�$�#��lZ�.hÿ��
-)g���#��<`Õ'�Am͈б����"1�� �����E#a��Ի�4��F	���ߐ���1�l�)oH����+�$�X]g�TN}��ȸ�^�Nvh�+�@6���E&�p*NG�#�=RQ��q���Q;�/䗎t�'F�v�`-��?����W���I��^��a��ķ�#����n�{x(�k�K@� ��G�+Q�t�7"�j-���FKhIMÓ�oTx��/VUdZ�f�}c���,'��jlE��\�Ov���L�<������d�{"�tl'M&�0�<�]};��?��fw��v+�[�WA�0�^i�����&�/�����j�8���'��������Dy+���OL���>ɞ�r���3[F����"d��Sa����R�[z�΋>��2C@K��� ����$�>���e�Y�+?$V,u�}WYd�4瓇�˙y���R�Y�[$^H^yZ�s��)S�Z�)#!�8����@v�ɒ���k[�����	�f��L^��C�+ ��	�P�M����A�|������z�o�W�V�Q^��܍��SJx�rw���4!2}�@������DM@�z+)6���\�� �L��h�H0�1��y��@0���a�ϻ���j�Z��h	ڄ\0��[a7$׫ҟߏѡbd��Q��@�K���ر
�$���R_ƧB�:��X�]L�'�R9O4�&��p���X�ȴ��7n)���F��w��o����UV��>�o���t��L5�&�B����,�[�*]������z����k��#!c?�A�I����r���L�eXLA�@�ޝ�(��w~����U"$���|Mb�`D����9�h�4fj}7��u^৳+�SP�t2QK��":w�!�o=a��-���i�/����|S��R�|���y9����L۴WT���u�;_����$��\�m�{�Ɖ����§��!�p��~�* ��`ӵusƶ2�SԷ�k���m�b�I�Bɨaá�rxn��#����<�Od�ED�����Њҡ+3EgM���k ��bv]Q��q�cZ���a�#��p�E=������Mθ�S'RNu[5	�R�\k�\ni*�{a�q��R�'�Y��`�{@��D���duBЫah[M�98ۇl��5�B�28=c]��4.1�'���s���<�P�4x�:6�trԑ��`��-��6�sg5A��ޏ��BQc�̙�ښ@^���v�)�4j�ȩ�R;j���������HU�ǳ��wy���|z�+�Iw����>�}�蕹n��v�j8D~�� �8d�q��+�4!���|4Ρ�L�ҠZ�%udu�?c��x�Rx�Ԙ���/�&�37��hW�l�5E62�*��JE+d��sGn�����\Pm�cAP1�Kבڷ��O|� �4^� r��\��/�7Y�z�l E!N^���F�.93;m?�XR�V�*1��8LO��M���Q��g=a��;`�� �{8;��R-��P�xF*�����l�V?��Bz8��)��Z����̠�ܛ�sK�&��`�4CjF��I�z	2´(��'���r�k�=�S����ꩌ��-�Sؓ��Op��h?8���!���3;������SZ�4XA�+S���!��}�.�#7���_�����ǧ�Nȅp<p���-� ]��_2I�bH�Km绚h�F�����INp"."�F�w
����ۓv@y�*���TDE�W��?��?tnn/�'oT���ܨt'i�E�>5;9?�R�+��5J�������_�L���T�ڄ̞�w����c�����.+� �/� ����{5���@�	���x�Ҫ;NFW�oG��p�v5$�󨂷Io'u�a`�9��'�����ި��+�Tr��<�(Yq��hݡ��&)Wm��h(C�!�.>~�3�
�#�.�f��SRx3/��F��ȋ9y��|��~����9����	��m�κ��o'�~o��)��P!�c:�&��P	WlJO��J��i,�d 3���G)�}�_�S��:�z�~| �_�E1�q���=�=[����o�ցC�8n��5�*/�B͒�4e&P�חp由�60r{��vorZ9Q�������ov�6��h�w��B�N�m�pv�=W�FB�m��wݟH�t�J:������^2aTShP��j]s�z��.cHG�T��#�J�'���Yܲ$U���,q��b(��#��ΞM{��o3��J���z�h�b���T��R4��8���eW��� ��IW����^5�x���E��-h|߀��x}e��JACp�֥�6��q?�V��t_�Db�ۆ^Q^nW)��$���q����*���phj�>m�v�1�j� ���Y�᫾P�m�(�%�Ov���Bkcv���+�&*_�(^Wݥ+e���v�M�!x�]pǓ!k��1�?������7���]��1���do�([?�~�|N9�z�CFw%;�#���?K�]h���Z=Q������4T�IT4٧�_�224 �.)x�gԳT�Y�J9l���f�������si-�'���5t�	ҟ��B� �"�.MWKː�~+��oV��EB=g�&ِbi�I���l��W�R��
��n@ٝ��L�i�^#��
lTϔ�	��{��CGyn�k�,����kiF�2��6�0kVp���&�4踹 좯'�&Y����~�m�;�����������ҝ�(K���c��O/2�^���<	��s�	�f#�9���/�n(=C��6J~Q+���[3/�Py��AQ����:q/�-����x�����{K��rO�Al���Y��)Ѷ�hcU��K�a̴S͜���E�&�J3���QNR�� z�tO��������z���Qv3�]�U���b�R�.��ȹ��1/�t����\�@��E��&`Q�Rڻ�:p���n�eԹ��C)99>��^kz�̀� ��.I����'%j~�����������)�pc;'ч���(�	B�|H�`� �� �vU]��[�b�X��π��aih��Jcu���/�v��"�^3t�|������>-s�	�u˜��0���q�ݓ�0��k������@���Q���Q���-��)��%s����W����YB��Wj�(�;,���u~1����\ʿ�8�đ���j�Vn'o���9�=��[��PQTE\�� V��/�>H>� r�uN;D_�}H��\t�h�3u�{o��t�q�"3��U�L��=C��7��^a�5�{�����mzf�H�ޝ�K�v�����sd�.��esHHC+o�F#TT�c�ܱ��N���O<�;��e���ⓝ�-J�w�p�� UB���ޏX�n�Qu�<��{>~�X4��>�.C�,�}�� ���Ĭ���B�|�D���^TG�2>�К�@�w����_C֓
0�Ɍ�����)nE�Ǧ/�� %�� ���OVQ�ԣ#�jme����ڼ��u{����,(��O��_�F0�g���`�)�SM/�R���*r�D�VN~����&���l������1��ǔd�sT�����=9U�[zm/�j�l�Z;��������oA���l�(ۨ�V�����@';5�	vrE�Ut����׃;��/D�2D�d;��-g)�#)alH�����W�U 8" �O��hN�p�Nb2i��R�ǡ�81��rD!�'Vo�g�Ѻ|�3��N�I�RwV*�PB;��[6&�H��7�P�{Ы��S�7�Y
A�@�7���ؘ��\��C�H���2��JL�x$�X��xpQN)3�{�|y���Dw!��Uc�&bd�AP�,P|*�'v���rY$��s�^�M� �_&F��@Y�	�Q�Fi��uoG��-�H|�����O��L��|v�����K�R�wT�74G�KNN��o����G�˹�9,c7��H�$����I�qm���M�	;��+���0����!E��H����&������墰�z�����T�]ƿ��U�Ő���.�"�tCH�<�ciZmd#�|�A(O�keM�ʒu�q����мMʦ�w.f=14io`�$�,�O�*��Irh��P�JJ�^��9Y��+��,�xU%Ο�yq^V�5�B*K"���}�PE}u33dL�ɐ�lsdV�d��i�J�j�ٌy�����I�j�SP&+gHV��<�SI�?.��G�?L�~"r��8z��<��̶D���B�z���;_� o}�O�ᇄ�_�8="�K�J�^	!v9E�)5���,����-��������b��d��q��|��2B;r^b!�u8x�"���g��g�c�1x̲eB�g�����U����ژ�׮$�<:�Z�l�~ͮ���qۙwl��Xt�6��e,*E�S䅒���xy�6�{[�7�)����Lbqh���y{��7*n��� k�x!�ICХ6�^`���_�L���N�#k<�'�N���C��(Yw���Y#��ݼ�1��">����O� �oc|��lT&�{5eҞ]gm�kT��pI�lhWE�7�4K�gǫOyyk  ��"��C|F��e¡Nf6G��ʫ��x�V� zX޹x�b�~����<���C3��}���2*p&�ٮNe�P�MT�>Nbu�"6�4609 _&��>)⤮8Ń����kLϢH[�IZp�H��g�9��U��"�b!���2:'|�M�����jٳx�i,P1j@qb�.�-"�1	�7mcr��Dk.oD��AP ^��<��H�[>�A�c���^yCƨY������\�s���ތ!C i�ن'��}�E5����L���*�܉��2���L��1gugȹ�݇kZJ�[]��NC2�i<!������q'�vy�\LD�I�w�~p�Z!`_���	J�"�	�ڧ���Rvz��\8���Ne�
ȸEY���įy��'�o`�z�L;��,S��'���X���uй{^G�Yo��!D��Ԥu�j^�����֙3�]"��Ļ��gz@��Sjp�DsQI2� x�fޏr���7�{vT �^Z�W���'�>����|�.{{�Y
q�!��D�Y�kb�t��^��W�����Sb�B�"�ˬ�����-��MbZ����b�_֚w��^�l�;� ���-����ܗk�a��BP+Jc�cူ�gS�?9���u�g��ը���~6z�+�[�bl��J��^]�=妞&�����0�h�A��Q73����mF �g^P&3���fHp��1��	A<aӵGmi:��9�/Kn���C�������I�s��n9׻8H�|X�MZ���~V�ؿ�������d8�EMvtɃ"@���0h��'��/��|��Z�|��&���bJ����E��:�o��]stVޤ��)a�b$����zo����ƍ���Q$�ȫd�ۂ��7����潸ۡ/��(XC�O�l��^("L	|$�ŽdKǊ��=0�M��T�����r�!��L��:�d_�Ar?�Rl%}3�i?w���$qdþ��ŒW�VD��=�q���૿o���2+f�ʴ��T�/ ����مlW�/R{�8tĈ�O�7��?�z��ӽ�k��}���^$UO�̕]���8�����_�F@�?��`+/H�6�ԝ�t�F˽p���LE�Ň�*��B��a�,�w�:l~yaG�86���2_r׽x��h��J!_��[����i?skMn��3I�a�o@xFh�\e%ޅaU�� �֡�$��}��;�A���a$	 �T�#Kg�Vk�l�'^�۽���r����S(K����2���xd=:sJ�J�K{��ڈy��� �e��8Y'�f�tfT2X��>�䳲E89��_���'�r�y@�|ñ�uI(�N����� ��F4�& b��B�*�%���d�+���8��&�)ޕg�=�};�J�K���/�'���!j$�=� ��O.|/
؎���j��v b�fC�DT���\�[5��[�'6,��_W��tʄ�A#�h+�Ի�a�1�N�;�l�2%d\I���D��(�kLF���ע�<��qU	��f[�Mڙi�hzJ0�G3�����-J�W�	�q�� _2�å�N4����
/H��"g	W�+>~|)�f��oJl��8�%���}�z�5Hh���Q:�K�qM�Vu�\��U�F}R��&�d�^�a�NJ2��Y��=��"����,a��iq�(�a*�{�3�%�з�|%��F�L*��gK���%ոv_��Ia=@����NXxc�����&�<�ʸH9�c�:j�Ze�#4��
S\,,RD� ���?�2��l��V�'��%�Z�q_��ﶷuO�nT��o�!B#�u2��v8�`��r��?X��SBZ�w�Ҹ3o���3� qV+IO�}FWq΁u�\��B�d��a�<�'�G�x��(���g���Tv�֍�	� �^��@;c}�O��'2���Jj�Ҥ�0OF�,lTV��9�ZL���p�)NfhyY�Uq,�"���GkV�=������u��sKY��C�Z�4�,GV|5N�4F�����ZfF�<Fx+y�Q�
k9nϦ�s�����@}RK���a�Y�1B�3i�]bp\>��"od��o}to�~�w��OvY��D��R��Y�����qwl�aPe�Ir9��/���Cf)���d��nRCj �H'��W..�79�a'?/Xo�-߰/REi�N�4���k��w������C��5��{KV^���<K�^�)ψ۾r9#��-R�^��B]�`�d��tx�(�,����t���W��y.
�m^ ����JL���U�@Т������d����-�L�#﹤"^�+w	5��<��kB���D�?�)'I<�P��^|�qOZ�� R�|�#� �Q�(��@�0�o�:��oh��۵�F�k3>	�(��A��a�8��b��S+z�j�NE����C�l�%�����2�U�J(�4=d��;^}�n��H���]��|��+Rߡz|Yɼq�
��Q�wm���W+A3xrӃ3���9Tr=�RK&0.�P���c���S�|���.4���~b�Y S��9̚�q��(�1���G_
��Tҋ��S�v2�3�G�����u*i��m�<#���$	�/>�������@n���YB��He�ϻ��(b���b���B�.�%���86�5��)oHx6G�x���A���?�
ᘲuKūb�h��h�ke��D�g���H��@"P�0%e��NB"4W�Q�5�L�j�1jy�^Kޟ�m���V	�.$��m ��-�?�?��V���ω�<�2��yO�q��n�� ���:8K���^a5���e�CZ�t�1#Ӣι6{�,h����E��Ӳy�kqCՓ�eE�e���Iuq�����=>#aM.���������*�o#�����(nr6���oSX.I����sfhĳ�%Un��1mT������_���Ns$��(����jKj��Vr@}˖cP�䁗F������g�,�Z�	����7j�����*y��j5����+��;�pQ����t���!�"*d_σ&����xL���b�a�b@E�jG(�aT��vB8���̛И����:>�C�x�+�ѽ �J!D�<���f�-f�~�R$mR���p��.�O�?ǃ��:����������tk�b=��1݉Ȓ��
]�ȟ�β��;]s���f;u���U�a<G����H什�������]��8#( �>Kˍۙ��W<i��_Օ��A��*R�X�&��O:kNo��9^��o94������҇�rF��Y����{���-ӷv�r���l@�����ZEs��	" �Ѷ�)5���G:�Tk�4:�cK����F�Ia��	�������u���7_w�:�0-� �ǖ@�S�|p��x�G��謴�O�T*���X���zq��m
#7~�m�7p����k�K�C������ģ�r	��0�MU�{��U�H��v+	/�%��q7m+sHZ͏ڽ�Z�uB:��!�M�X�m嶶e2��j�(����.\�uI�&����6b�ލZ��	-��&�|�q�8��Z�.@��GꡣR�T��=ɏG�	Z��7�4�	ru`����m�M�.v�Ny�(}\f�{������щʋ4d�feK��0XtB��9�M�-7Ex ÕX?'��y�8���Bw0�2�w����[�����Эb�b��5��`7�-��]� 4�{Ҵ�IQ6^TB[#APÅ,�=΅w���3e�4,,Q����ڒ+.��(�
:=k�+fzu~�����vm3f���������z��k��i��#��l}D�n5��.�lI�Z�c��=R��)jNX�����1�i_�����Q`썤�f�Tgg�Ɏ���@��_/S�G�oS$
�-3ފ�>����!hO����>���X</(XHI:%c��%�~0e��+{�A��(�v[ĉ��hvB#�QjJ����	y���W)���7���	��/함��| g�ؘUkW�c�m���uR1���c��I��`}��̦� ��)������T���*dhq����!�C�Gn9��ӊ���q^����;-
I��'xÏ|�ɭ?~�<�8��uQ�3��{��!�ɟ�����$�Mĩ{�P<DϠ�/��.�a�blA�m�!��BR�f��/A���|+/d,�I�(:�zA6��z�Pi=\M���'��"&t�?mK,_Z$��-�i�Oj�jR]c���)����t'L|b~��P+�z��L a�a�����y=��>"'1���-�8=x�p��3�=�C�C	j0m���-x����hX�r��������F�vq5�=��\�p��<:����b)��p��0*87�2�a��'�TD�ܷy�Z}e��c��]탦Q��و9�F����z��O�{�5wR�H�1�������&	�s�[�����t��u���|��r��<G�@0T�����OI�V�B<y�w�&�a��������B �n�B#D-�W�&K�b*�C3I}v�Ȓf����s�f�5O�O��'Ӡ��Ż��x��u�ү53�N@���߁':���Y�Y�5�a�}��aCzb��:�{	uzJE���`��(��$Vm(IR����� ����&�p���FN+����&��d�2���Vi��������(z���
�ݛO����"���8!���P.S��ƪ��x>]�$R-U�dz����E,I��tnTd�Y�(a�6em� �}$X�PJOŬd����x����RG�~��q+,�A�Tm,��� |̉�s����%��H���U�Xgr;w�``
�C�/�Jļ"��� ؉��Tlu�U�ep���s|��E��.��^�%\�����	��_+T�8��/�O`+����Q�z<���;<s#8H��t��u�h$�v��y�o��*�i�|Y&�&�����?���� :�=#}2�U�V�]f=�bP�J ¨&b���A6���5���e�%�yeWN�u~����Z�8��X8�=p�k�I�Yؼ�O�r�?�T���..�XT[�y��341B���Q��p��q>|[;Z����O�"IT$����I)0��hWL�<;!�ٙ6���E���k������>H�z�����qX�YG���`��uBw�	�d��Vu^�n��Zݾ�����Z�J!\D����ƆD�x�G^����]��[O�^�p&}:vݡ��Xi��-V��!M@�0�q��K��{����ɭ��_�� 9�K	�����@<'Y��j��==��WG�I:����;1X�V�Q������LK�
\z[`���jޢ���j�����<�.�-�tCJ�}��P�Ÿ�72:�
r��
�~�3y$ci��&2��9+1I?]ka��e�03)C5��Kz���%sS�?`�n�ׇ ���`~ط@=��J%�P��Y{Xh�)����-�1 u�E��y����M���ߏ�JCҍ�֭&��ac"��ʍ�9�J\�_�U3S�bݰݷЌ��;�:���yɥ�l��#޵72�V�H��>���!�뵕��P2�C������2k������[��4�WQ�9�#�rͿj�֥�yu���Cn.@6R�.["�u*68g�a+u��5��}�d��^��{���:�76�Z�D�ttߐ��:k��;���ތ����ҏ ��mm��lR�ڭ��
�0Z�����kc�i��d��c��l>��ﴱL�Ӛ�B�lؾx_��$6�
�*�(UU�Q�KӮ�N�������Gd��JU!���r�;V��U�L�����_�$~��{!bv�=���Ӵ����_dU�r�`��n6��/����Z2%,i�a۝%��\� .��X�4mM���t�DO��-$8<��<R͑G�1Ao��l\D%��}��8���'�k]~"��_��1�')�H���(fWI:R�ڄ{�îa�E9?f�,�@#�,f$q߃5�����o���_����o���䥈�%]�>�f�:��9)B*����\-����g8֠�ɀ[ac�L�����E�� ��ӿ(�D�z<?��v¢��o�lG�پ�]����~��)�c��T�.�Tw۞K��7�I��+M2E�5w��|UK`h󥫆wһ�?�jlCrD O�~��!u�U��u�����E����������M���4i�f���`��<`=��zwa�o�'}j��T�<�X�"��s�Z��fq@QQof��|9�[wH'��/=�P2_�}9�&���Tw���2��5�굢k*�6���+���߸�+7��^��<q����D��b���:�-?����t�u��?�W�l�X�#+5�:m����qz�J���o���$Mԏ��6�ܢ�L��b�&�84��{%zp:ٷ�UE�3ge�O�׸�����ѤR֮�����r +���FsH��u���L�˙`p���(Z�rc���]������t�o&�&N��%���U���W�sESU�'%"��F��f�#�i���[��
�.W�߱/��<'�Sj���{՗�%��BJ�����>��3z�^��n�,I,��-�'ׅ+�6�uZK
2��8_�F�q w�z8_,�T�����F���gq��TJYziG���U��X����������dW����_�F ��c[+���y��� Vh6Ղ�wc�P�'�-O��ڄ��^xF��;��dsh[���/4�	t)�x�fGM��tJA��R�9O�n���W)g5@5��� nZa���[�׉P�#N�^B'�?����@�e:3	\7|!�n����v������#��JŞ���w{����Y`����I�l��O` �d�,(�	�<�>�������c󾏾053څ�erS��kB����:��ē/XN|G7$i�U4���~=�~�Fwh*~�wTI��:}�˛�#�p�$��G:cz(�Pf��Ѧ��=I�
���\�>8]���ДV U�W�\I�)����
�\]��	a��L�Q6���w��rm��;]�9V��zhx�6�׊�;J���Ms������G���T`R�%�%;K�A���E��'q�tXX��j��Xd��3!����0���Q�[�6��4�p��ـL�� ��%�58@�� �j�*#ȉ�2�Fc,W�U�Ř�U��Sވ��a��GR��7�@�!6���¡��0\�l���%�5��h���i�)��'�g�{����*O�s4Y��v �W�\o�s�ی��R�"�9M���yz{7${w�J.�x��&��,(� ~"B�lG%;X(�x�U:��.�?-}��-Q��z9�����5���-�	+�'Ko��5g]WV8g
��ehX9;��ڨ�{�b�X���+b�G<'l2�2�S�Q��M�L��c��<\�I�l%��B�37<�8H��#�L����e���|P�c�&�V���]W��'bղ ����X+��d"��v�����#��S�b�=dR��O�e�<)k��C`�3�`������ N��-�3*o����K=��̅%�ޜ-L9ɱ�6�wv�
�ΰ�1!3���^���y)4ăT�c�W�������a�N c�5s`h�-W�y-B��m�a�Ԋ8��8�ڔ� � ��W���TL7�r��7�f#�t-�5�q@��v�=�-91A�$D�>9{�|����o��
P��m��v�{�,�*&7�z�DH^p�}���̇[tLm��0"�f���?���Q�G��/EYCx�� V��a�:J��W���?�J�8�`9/z�9�`��;�Ȫ�"�݅M�"��\?�W�qj
����� #��V�q]�j��������$���\��_Pe8;�\��"]�`���
�|(#WQ�L¥d�X�Ƀ�.b�:��P+Y�Ļ'e{�,9�D,:e�P�P�$�=�=�Qs���Æ�xs��O��A��,�k3��6��>]>x\�vK��x���-� ��Ps�Fq�_���	rC� `�;�.�ϑ�=���ʠ�+��0��5x?VL����������δ3ܻ��E��b-5��)��7����Q
\���1��r3�:���5#[�M~��An��1�n�Z��vJ���R�dq�&�D��,��cks�U�I��ax����;
`�W�ǣ=��]'
c���Rh4�z, 	�M���t�!�1l�Z�%�S��qb�4�+�X[S��[V����U�Ed)4e�Z|�sb�V�u�����EbA����ۺW&lJ�b{�H�g�7�l�h�ڲz���}��5e=EẈ0�>^�u�lP�v�9*5�oc.&`�-�'���ڃp�Sƪ$UZ2/�.�2Q��a	���!�lM	TC@�ۡ�^,	��<
��揗!Ě�rc�	�����UG�}�_���� ���leJЇ���F�gx��>T����U�Z�}a��Mៅ�,vv�.'�zB뙃r�bոx��|�Nll�t�2LV�\���j���&�1X��� Q�������-f+%bȃQ���,��������޸�t�8�=����1����P<}�!�ؙ
�t폡*��f�ڲn6'L�4������U�F�]�M�����P��lI)�L9_��TW�����jE�Ă�r�d� � 0��� �~�!�gCl�̈́�<Ta�4��'ľ�hA1� ���+��#>�G���{���P<����) ʑ�����d�f�iw[�E��q���F�>Nʽ]����e����P���z��~u�V$������y��N	����)�������+�VL���VU6)�<���Y��YC��t����4W	�%E?���[� �q!Qa���jF�����i����T����$����@
���ut���x��������-��joR*���CK__��o����v�	�5Ǌ15:?��G|ɞ펰�T�AGe�e��(�x`��|.e�x�+�i���? t��t�V����VFP��W�0�m$2�ָ Pq���}�:��c�+�!�]�9U�L�!�� er���;�aذ���L�G�{����m�ij�Z����4��o��js^�+F�8se����Ã��d�ǹ��j��ޭ>��K�յA���d&p(d���{�p�S ��,�^���jM���Z�ZPGp��..��?���5I����4~]C�i�/8�%��q�"�e����S��
�ݙ q��4�)�B~�\���SsE�a8��X 6Unv�1�SR�A%���qn�t�
k�nQl��cy.�QV���n��s�8i�"�͍�A 5�'�и�[�8��