��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�ͮ���,c���d3� # �z��d�O��vVWp� ��|F0�Ѻy�����ǌ2�#+tIfA�P��(&�ӝ��pԟD�4�j�a�S<4R�#�v���UB���x�&�C���f����D���X}Ȫ��0�I�g;Zq����À��p���fD4(స�Y��2)�����+2u�@���q[��� ��ӿ��5�&~��x-f�	�G�EM��9O�nqҼ�htlo�c���dwV�ov`hr�]yDz�mi_>�~ WX�e0�Z�;<����r�U�:Ǐ_�웗��D7Ǫ`�s�QP�|!fg�Dc r��4��2��3
��7qގ&������;�-iWJ=���q(dE�?vwnv�i�}��^+0=��|��]���f�r�Pu �����8g ߳%�ô����� T��U� Z��Xb�6s�
��A�X�$��N�1Y S�'/��>�Q�}���$akN$]��y�ԇ$E\d��B@Gv&	��������b�݈erӍ�b�F�9����,F\e+7i�!D�G(P�,M*�q��$��Y����. ��IU�����F�s�c�� ����#AG��e�~��6�^m������aw������e(�8�E3_�d�Դ�VP��	N��y��Z��X�+�
���Ԩ&��,�2F=��F��?��.�7�Lr JB���̰�\<��ٟ��v�>��0a/eF��jC��#�+Hn����v��`S԰�����A��������M�`*B����KK�#��)V�z8����sʳ9�rE:��*"�
���7l �z����h�#-�yiu_}��f���c�z�Q/5Ĭ��W��'B�$��������9�NK����_ʪ�[�>˻��oY���� ul��J����dY��@Ԕ�x��4Q��%��c���e4�0���kv�=�������f��Rf})�ɼjMӶ���¦�$c�XZ}�K�%�9�T��$=�S��$Ѝ����๙5�T�DH4wV��������`���ªd����t�frtF}O�A�sK��+���P�`�.�0ٵG��w�8��D�v&E�ma���((��L���у��B��)n<V���b�#�ܕ�\����?�$����g�$L�Y8<ݫ���[����^��U�e�hgC��������9��G� �C�T�#�ؑ��O�O� i7���r���V�iڤ��_��b9����u�}�Wo q���8	�����m^B!d{4�T�����?�Y�1��:���& 	��?;�0R=��W��l#�$p&�pՉG��g�VU�+�j*�o�'������ЈX>�	>�~��;�ණN�3	���kR��>��'쯑�愭mY��q+8�.��W1w+R^�^a]���j���H|J�9���0��*h�P��ӕ�FJ4�!9�1Ґ)���]_N�6��IP8�D�����l��7r�:&9��N�2��6d��@e�(��aȬ(�����=�r�N?����_�	U`�*Y��;9t H���jU�����VK��K����y�)�ǚ�,ӱS�=yz���{W)
(b����E�h�$��$��	B��9��HΨ�ڷ�J5z6�H�����ߑ���eɿը����cۻ�����b�g��Ӎ�w�}��j��=,p�L��̻%%؉^|	�1�K�0$�B��@V��=�O%���I"� ;-����ś���h�k�U�Fn�M�t�[)鼓j�o��ҭ>*�����3N�Zt�����xiaل9�Q�q(=�!�W'`U�{�+�:ۛh10O��l1�!�ugC�N~"9ĺt������6n�=cDeV��	�j�w�,�Y�X���*χme�e�v��%awX�S���=���7��Q|���񪏑!嬪���,h{̼�}�_�Bkfb5�j�j��BG9t���V-�ǵK#ί��@��o��!������u�	�nH]}���V��&y���h>C˪_JH��%�Š�c�Tr�et
cԓ��r!O���q��mK�GA�b������c���HJ5�y��>��3�	(��:�T�Yz�"D�o �{������|����	-!�zi�I�3	�g1=j�C�/��Gw��k��Q��ߗ ôNMK�,��:��8�#�Y �Շ��c1��j2��E����dXR��F?M{ �w��Z�����m��|�� �+Eu|���՗=�3�a~��A �d����zڜ������Mc�6n6�X#q�-p�Wa�ɝ�	Z�Y�_��0��?��s�5�X�I�)�;�|W{V�O\��AB�W�M���m����Z�➺�DPs�qPt��3>�'|���_\��o�+|���Ӕ8�i��{o���0� �^�8‛�9%�+˴�t�˫��>��X���OM�0kK�͒�649N�Z�_����|R������ ap��M��R&�q3�5�c0H\�d�R�Ħ��[���fMv�xѷ��^�~ȡ�lY��!����w�FrQ���|32�7 �)W�n�?^'8�\n�����1�� �B�3��2��.�O���[~V�/�ݭ�}rz ��|�������pm�QK��]�I�[��v8(Z�.�AV�)��#��a��ƥ���Mv
v��L��)�����''���W�|`��䂍���yG����5wY������"#)*�fl�8���[�����<m���B��c�W�{?溲�N`�s ���m`�7�t�i�
�1n�����B$��� �
i���inԱn�����)=!�swƭ�S���E��h"̂S��sN��R&��/���Oq|�ψX�U[pXS�pkl����7,%��A߅�r PK����+��&����B/s��S�}�ƪ^+)��{�)B7P�xy�
��/n�3�$,��q��d̖A��ĝW��x����^K����j��Hw:�^[�M�ԊOw��KBA�?�>3�m>N�0;�VVٺ��]���h�AѷJ3�;*���Z���e �?ǐ�6I��)�+$�<>��/~�ZݷQE�y��8S�S��}�N��V�-�/��L�X�atR��ݛ���3ɂ[�:{�:lgJks�r[��J�k�l�	��U�i�	�B8� �Nk?���!�`�	��>O�����tƜ�����a'�o6bM��5 �ǁ��b=VF�/��?zW.��^�d�����e�.]};�w��6 �>;FH�Cw�l�u8aT���B��<�|��fV�|�p�CԺFg�BN��="�)'� 
!�t�w���+4��y;�CJ��^ ��$K&R�����ҙ�R�������{����˲��8Wf�:�+�Mpu;����xS	�)���\�}����]9�ƾtE	�IB#��aH:��9W~CrY���r�=�+㿭��U6�1z�0���vǜ��Bk0�m�·�~�g�X��$=-�o��!m@�m��� ǁ.�o`o+v�u���D��G���W��'�KB���
�Q���$�ITo���3|���-
�g$��]V��u	�F2B#�f�ݠvo"���m:j�njy7������|��$5!����g��ٻ-;�k��*�ׁk����S�b�V�p)��jP���R��8���B��KZ�9J���V�`b�N�I���M�<�Cd���j���X��ß;gz�R��p�� m7Ql�
�}=��@�i�d�W��ߦ�?:�W�o����-ۅ'o�K;,�R[��F�����<��S��r����$؎���/y���q�d�sqm��m1#\��w?�V�O��'-ĝ˖���5���7޼�X�(�����^��_�~$����@��n�]8�ՉIo�e�k;��aT��MN�綡� ��4�IP�3�˻ �;t�`��n=�9�V������+A&�4�9΃@J��N����w����X_���(�
xq�i#�VՆ��Z&GOO�i&���&4&��;:�����r,�b9���.ޖ�R%�F.����1���q�N���hP�r7^�����p|�9~���{���<~��R�*{ۇ��6�ԧ@T�׎k����|�Ђ��}g{���������VΏ�"�F�b���	��@�i��W�M�ʽk+��i)j/#6�3����� :��x��uKhglW��g �G�6�Cή�&O�՗#v�8�����"֡�֞�_�U�̩ ��VG�@�C�������L�����(�!��s����v�i�Ln!�n/��Q@���9��Lg	��B�`4�1}�T7�H������>�RhG��K������C9�4;�u��acv�.�n�'�|��5��?Q�.͍�]GP� ��~-U'�Y%=Ϸ�Uȣ���8��(1�Kn����GE���M�휩���&m����K�yk�RK�q`��]��Vr#�ӊ%�+�H��������,d�+;�d}�s�@TxlVK:�e=j�!OE�}{���r��B|�@Z��߯���MϞ���1.8��(y1�k�G�#|����V�AZzgI��7+j�J���v]�j�,F*/A��c(�h���yw�s�Dd��5��	; �N~^���E�)v��#<�y��~�V��7��Bv��"9�߁'���E�@,us^�r;��N$6��~d��g���W�����ZG�~���0�uW7�d���L}'�e�9`]�BK��$��Ҽ���<�.4�d?���߹W��V���]L:�������@�.���`,![N��b_|�c��l�߽!�[�q�H����.>� p�lc��k�h1Ef��f������.��õ�2���R��2hc���z4yQ$ſCV�yhT�[����g4��W�w<E�.%�e_�p�,���i<q80`wA7��'�����i�c@5�����P
 7M�����΁r�+Vk�=���G�����������P����1����`�{2��,݃aԳ��vsp�O�A�g�Y�b�1�Zc�l��^-����:3�I~����h�'z�͖y��%P��^EJ�Pf@����%wk��_�X�B�����!L��(矣��0�kd��Z��l�&O�7�:T�+��Xκ���x�*��G�4ݪaN B�e��;�d��Ԕ��� !��a��BՃ�7yj�Q���y[���	��;j�=�-ٌ�)��繺�9�e#�x�c�ǝ�����hv�9�v�54غ�9�}��#+�U��
�o�g���u��&Y蒓����?� mS|6�c\\īl��>GN�Z>�t.z���I酞���u� ���RV������kߘ���1c%~�Y�L�1@vhE(4��!9���.���ؒ1ݟP���y��ۘW=\�N��9�tB%�-��d.�ț��#^�2V�(ڽ�w�0�*p��.@�d���4���k�"&�T��7�!M[y���m�K���CYkp%��s���ʔVl����@���������@�P9��
��0���@�/�Bf���7"R�~/��<r�+�V �mp��n������c���`�?����VE�F��L3Ր���8t���9�M��RZ�b1m+�(��)l �>O��;���87H~>�@�a%x�h����f`�K0����kc^�l�']��)K��GG���F�'z�Yx����5�X����x�'W\��j��>Z(z��Ǚ�p�oP�lN�����B��$ņjk�e�˚jZqĠ�ޗ��+�V�)�Ac��1����B���,�������[��U##�}�Z¯{A�ۿ,�v��f'u���Buk��Q��n�thO���F�{y�RqdQFN�֞���[ǿ'Z�S������$-8��Mo!�Q�0"3�L{�P�����f��"Q�	^��*\L ��������z�W�7���=���QV
��y�eG�.Ƒ�6�f�W���q�+k?�a4h�*}�Yx�+2:§� �B5�ņ���A�u�1xm�����j%A��Ev`E$���T��L�x)l' ��s�`��@f��xF�^uJ�Ft�t�ƛC�}�C���I�S�f�R�1(���@�t3�q��)�U�l|�ąky&_�][��$͢��SR.��\��mUh��r��M2�@R�x�\[a�Đ]�+&j��d���$!�V��`�î�bX24hP��m
��ECB���E|��o����:��/�:��[d}��S�A@���;X�{��8<��V039�J�o֣`�ŝ�'S�}���4@E�¡`�[j���FqO9��@�Ǔ�\*5h���JG��c��i���z�A�ǯ��F^�)M��74p
��nD�f"��n�m�G/7a�	U|��߅�3���[*�}��2/���.*�[w����������M7�(�"���P~��BCx�XD�BbT4�Ī��
�oA�v����(���bN
��Z�q70T5�
_g$B�Z���&�D
S���~�~�S�jd�{S��/�����f0]�����nm|�K�
Z����,|x�C����	�E���Pi���ł����~]�*Rǉ(� �@���ЎS��}��� �N��Y���T6d#t�z0�r��v�֘�sQ�«[�%j��B,MK8$��jlH%���S�إI� �5e�s� ;m<'Չu�/=�p�Z�� ��W��u���𸀝��'��x~)=$|?�+���ݜWl��E�	��]�tb�)��ŝ�#��[�\6%��qC\���u����\
N-�zG)f�G��=�`��Ӟ6lN�l���Qr?�P�j��*��SJ�o�L�س����7��}o�&�[W��ݢE)�׭�.����\X1��'���q
܂�j�ӊ���W� =:jz�!s �`n�NA4:No_^�`߁}��3����S��޷"��C?ܙp�U��HrC�N���b������q��e&q�f{uU�jH������5���7�H�iNO�~��L��F]#F�+��������A��Ntk	��q����8�����!<5�\R)����@�ے��`���FK��$b`�D���;�5A���Z4��|]��'�A0Jzi��a%r}#wMXq�z��8�M� �Ã��%�(ٯ�C�%�L�u��*&�-"!4���VO�H����2��cRL��v9��R�a�8��q�1s/��=o�/{��j�du�/&������������v4��G�?���r�����^/�P��/<����|�-����9bW���������=i{���G��#���+�:��0�`աToiؽ���,�FA;�X$��$g����0T�:v������<a��;�zOp�WV���6ڗ~ع�nv�|�H^�^@Z���M���l6�񏕲���B~��x�n���	���*�c�NQ��@f8wj��
�:��ȴZHc����1EJ!��s-�N���ԍ�]�����%(�"N�/cQ�VL���;�4���vtX-|l�
�@����&p�0E>r���� #��s4�[K���6zL�V3�۔El�����{����<�����2M|>\WS�Ǆ�z*.��n�z$�D>�|�Hͥ~�M��^q�Us()��^�՞�Hn|�w_O�������[t���S�Րd2:�G!�s�ύ��|_l>e���Ƈ�I���ɓ� �=�������_�c���O�Bh�B��J�՘6W$ObX���j*�1R��f�"���5�u�T�GB�pǑU>U8��� {��cHK�o�ea������w	��֫�$9��K��יI��I���o��g��r�hŴ��*���T��TP���4
��
�;H�����!W���	�e��T4���1CC���e^��&�#en�%�b���/��H@��4�m���8�r�8z�=q�/��u:Vk�U�`��G���\m+���#�(ϐ �C��24�e�&�n�ʇ�.h�dF����H����m�#!Knx�xf�Ο>���(d��]8�q��e�&��������BY�JX�W}yȨruo���h���d)TP����0��A��:��^	҅q^mVy�B�e� [�ROX�\�Tm��򟹓�P�Zd���EFQ�"y�r��8f��[��k	�++��(ۂ1X�}�{�p�s��WY;�l�L��Q�g�ƚ"m9�jq<ĕL� ��_ӯb.J��I�5Y�A��#��VZj���rxw���!��̹��	W�fOS����u�Y�BoQ�d6*��_%�'�ބ�m#�o��� ��2!�v9��q�j|�\$<$��͉��B502��B��4v��v�ނ,�N���yWݷD��40���;���[^�Z�[D���|��H�Kh�=��w�L�գN��g��4�i�*N���Tb��쟖�X���9dW�e�`絭��98�W�5I�n ���T����J铜�$'s4��p����6��\9UD�'�x��cW���B����ж(RaR#�rT`�6����殔���8�EK��D�?�Z,�`u�p[ �|�i^��:ZNo�]�x����z~\�$�,��5hFZ���ml2�8�R?��F9�er8�J�k��n�]ۼa�8�Z}�.۝�[.�3&��B��2Ƙ)g�^$e �ݵ��z�ɵ��Ĕ�Y��d�5��)��kQ	�u8LH��T�U�d����'�/y��}1��6Dk(� 76/��e���-#��;J�$��ѵ�};�c$��A���?�ԉ������� NFU�6���QҠ�R���F,x�Ǡ�t[z�˩�d�f�x��;;�O�禓?T�ۃE!�LL� A}�?Wh���+�D ��^��Iַ���k����<hp��Rk-8��9��g@��^�,\��gD���䎤�_e��2���B�AJ^T���־����qj���vRy�K�fHqGu�S$F��ڢO�<��^�� M[IQQ�{_��y_\>�o�gّ�1�Ao��O��p���Y�R���敬|J%�oҵ�'e
2Ԇ��NM߆�K����kpwBiy�']9���c?Q��P�]��������܏:�i�1��K�	%���fz�b�q:Y�Kks{�B@�m��V��pxӱЍ��0!�se=C���e�F9+Ί8o����.���	�I%��p�51��@M@"S^�����YL��O-�����8�Dއ�=v_��VH�`�^C���6 �4�ɘu=�=n+q�JÐ��o�@�C`�O�y2N-,��Dp�����B������"��"J�o�Mc��Y���Um��3?'Xj��}+&��ƴA��,����p���$���P�/`p�#ޞ�y}�{�.���QI�3���9)�h���H(5�d���g��4QKL�Ds��C�����ю\���6y|w��y����W�����g�����NI�߸5Ν׆ *��D�`�#R��ש�ĉ�U���H1h��0�Wp��� ?t���M��ۛ�ف��¥��	��J0@k�'J���5t�řw8_C+�	�-��#?�[�j���CM�Z��(�r��m1��0oyЅ��cj^X���,k��4�n���n�K��9��ڮU�þȧj�DRɏx���(�*����wϠ�sߊ�A�Ƌ��]�Ε�'���h7��/&���|�YV:5v��Z��2°}�_A}�8�ô�~3 ��4����ݳ�
:� b�tܿ�BOA�����[���NV�纒>XG����W��1^�k�n�� 0�տ��12��TQm����XCQ�>�w֗X���~��˃R��ؖ�
��KX������A�B�"+A�mJXVX?t,Y���ۇ�@����l�_cu�ϯΡ2���w诇Z��n+�U�(�D�H�D����'u����Q�{�C~x\���W%7�]'�:I}d>��(�F3�fr�ǃ�R��D����-«u(���՞�=�.�M�%���r7 �r���u��>�h��n�D�)���tKě���^]�4�WJ'�`7���FڗrM�7�-�q��a���� ���?к���H� Z#���;����C]Q�ʞh<�J�=�E��M�I��p�]rt��r��m_}"��a� �yDJ�!Z}Ϊ�d��0�\[i\�C�/"P�7�7��uJ7V�+*@�&˫�ަn{ן�YU�� �~��r�tD��H�!�]��g�a��?]�u;�"9���5�����jܩ���7޹��l"~V�m�F(�咗��>��D�)c�:�
��Ы3@�(�5D6��r����-�ћ�g%0ܥ�$	
� ������!��w���q�mϧ�4
�7��`�P;�ҵ`���:�)^%����Pko���~�0�^?���n�K�K��O�� ��Iq0�mw�|�J��-s����c��,�t���J@*:#q�XK������ �6 |f̈́�0,��T�5���Y,��t����aD�Z���W׸��̫
/k9hV��?ѝY�܃}�!��I�kjb����7ݖ��⋈�N��bT8Pc�a����A3큟J�OHe1�n�kc؞fd�"��{����?��%�&ZS�=:*/[�)E�Us�5\�]/�a����(	r`�FX��xx}��gsG��E�~i� ���a*+U��Y0pDܲ��p�c+Co"g��Q�θ��"�'u�ύ��O"�s(h��O-
J��(����k�F%��>,@� �ù��xA�y������.;��hk�D;��������ɪN�|�����ѵ� C�ndRX�h�6�υB�Ii�/�c�{��M���I��_;,Wl��a�t��Av��#}�=�6���#.����F��� 4�q7��fps6[nw��	N�cF�Tb̷���2`��9y:�'��i�ZGX]�W�?�P}v!��aՍ.����vk�w���W@D%�Ր3<~nBL�"h5j�g�#���kP5�*�@pT�	��b*����_�6@��S=���3� �P����W��*G4�>Z$�|�8<f���̆;��a�VBT1��w�-������|!���-\ݰ�s㘼�_�%��![�Q打��%��n8st������`�����菮p�o�x_�.ݜ���f���:�׊�}0��#f�����uyk�I�W=#!>c����^����x�jp<��������K�x��+'P�}ښd����D�.V@)�4���q�1)MtJd�.z�KD��[G��V������T˷"��y��u� �2�Ga�K\�(�`�n�(;F܉I�aPf�m�K��"ז1�ge���ul�ʈy�1ݎ �3r����1Q��uF�S��� ��a�	R�
�g���L&�����u����'[�4<�"34c/�	d	��0�o?�{��U83���Z5!B]���'C8�����g���o`g���E����\nzN�bS�ZKR�������$Z�\3��σ��W)%���@5!�x��"V�\�r�|��L���;�n�8p�i^��<#B?��8
֋�?67ئ�L��{;�qպ�h�G�K��V�N����]]�{)�̈́_/��ċ�Y���5f�8�av�����3h
@@Kc$ԛ���1b3�������cੂZ��>���y��j��9�e�0��~��x�V����XeG�y��l	�NE:Dj\�?3�;�2�|�R�l�?��]*�X.<�J�{Ђ3"H �l?�Ur��K`�l�E���Ne}v T�4"#$���c\�G�t���"����6t.(7�f9�A~	}�!�p�K��}��4�G�1(�M8bc���}R���'�*G�p)�Ӡ|	�K2��8IU���9c)�QU�A�PV��ōW�>� �n�b�-�k���p��=�	6lm,�{�pq����X�	J�1C7��69�4��=H��J�X��Y;F�U0�^�� �g����aqy��̱��!�1���ef�P�D��gkW��Zk%s���AM��
G���Oa���^8|�� �nDN��!������t8�/a9�((gEI0v�s�T1͇���>��{��$?���A�t�b�������ߠ�)f2WAv�ԛrͮ� P�T���V�����:�ɞ][*WG1kw������U�#�A��f�Q�>T6���q�e�ɧk/ek��۰�)���{	��Y�X;>�
``�u�a��vX�Oڊ�x�1�'� �G貸�;%���S���@�"h+��ʬy4$��(��m��8��غ���0A5�ů��ɥP�!���BC�_Kc���\ �Z���A~n�LbZ/
w���7;Ώ���T��Dx��+��%f���v�Q�i��'�X���<����%��|�܋��u�\|�i�KM�U�τ��GvxDbp��?-�����bɔ�_Ѡ}r+������Dk��kV���)������X��c3�;�T���D��j��$UD�+����� Z���P�1��4�U 9ږ*�Ks�k��q�z����=|*di��o�Z2�4;g5P���CDO/��v	��Ӫ���/.�39Vn�n��?,�*�T����K�� ����>����U2؁x�/a	��uo��|.̃$"E� �Ɓ� �x�"A���a�<�SnSH֒Y��\��M�j�dI���HCy��6~� �E��:���:L�6<1sN�λ<�*�`���4���k�,��b|�k��r8�ok�oL/�c��I�Ǿ�_7��|��g�`m% D|��� �?՝�5�`}�(���:�)A#�GK(���^���	2[�tI�q��9�t�i�n)�(k�%n��$4fb�sL��������uL�Ҍ&�5¼ 6��z�Y�y}�$�9FA	b�L�ߧ{ulQ��S�^n�/�����GS��M��,u⻳���!��&���ch�-%�3֭��6?K�i+ {aѕ�s'����K�,.&�`�=ѽ�VoOC}�4�٪k��R}����Bq��#H�/ ��xK���,����K��{�&���`UK����!�4+���*hN��̓�?��k����<�Gl�#*���Seo����Yu��9���#_;'�{ӰR+^*��4cGMa�yt��;n�fa��a׌U����%�����tE�����WW�j^�_S��&��[�a=~��c/��ӗ�����[�N{�eQ�$k���2���Z��"��ǿ��L���u,-���a�ͥH4w5ʮ�K�[�)���1*�knJ���=��O�7#�d�]�Yq��\�����P���Dd	����
�\�Bc��;\���Vc�7j�d�7�Kξ��L�����Y�DJ;����V:�c"��Af'AD!D����1#��.�=1�S�"��<�z㫴66�O{��d��DG��:H>{��6�,�OY�d�@+I^�}��*�wV�f���M���T�|S=��f��nqۥcv6�ؚ�I셤)�=O)�D�U�L��m�B��U�:	��a
���z�֧�i����-�H�+��AF)�ьW!1�V�n�D�{Z;Ur�ehg�-�z�)��| � �������A	5�4<
HZd�^
��� ���5�W��͐ůa/�c�q]���3�c����;Ɨ�������С�a��y3��U�f��R�(}��3W�m�~g�����7�u!*��M�n��*�~����2�t�+��'8���}�LKs
�Z�!11yPb59I�n��ذVL�搡�7�2����:����E������/<��"�!Q����|;?���, 
t��J�@�:?�����V�ʹ�r�A���.j"��h������Om��`!U��� ws�,jNtL���	I��y�ă��� �u���r�3�(>m��̊���0[���Y+q����r�Ĭ'7Y	��h~����yq(,����#\��t�Z��g����_�G���p�^��|%���i�@A�\Z���z����.�
�|��0+v�xu��h*tD��]z&��r��.�]#ޖ�!ޘ� �iuP�m���2��*&���k�d5c7W��8��.���!������U�~�'����I�,HU�?���ӃVK�B�;��U�� *�iH��prf���#���2��	�]�`c1�%��*����jA�S�Poy#$��k��%��ܓ樋�b������H�N�����W�.c�#Dz�&}�O����j�n�m1��S��\�i4�*�w���B��-��$��9XUa�
n��M��A�����E*���c���CA���'{�~�b[�ӥ�)ob��LC��
�5*��m�w��+�U��mǚ�o��J[iD�������Cֻ\<&y �	�3U�C��>��a'�֮f��%�[�_�.03k!��	��oЇ��w��<�׫�^�m��@�����C���H[��A���ܺ��)���{l�j���%�t��?� E�m=�%uj?�U����]a@;�[�s��34�T^.Z`���F��8Y6� +1�,.�(`�˖F*��nk��欚]�#J��:���h���4m]�VP 9݅g]�@�E��kƳ���⒓\���E�0�-���_n>�s�����������R�$T�c%)�,ʝ���|�x��M��Н'8��Q�V"�lX ˸|a<���m�v����L�m�>��#����}Պ�7`��$ű����׍b�uβ����>��Q�Ը#�q�~�fΣ���������L'��'��#���x�	2��/j�����'�f���׮��*�j�:�����lbB�lO�-��W�nW2V��r���������h���X�953Ww6�%G7�c�4d'�U�P^�튈~{���@�aE��9�CRj�"vH �?,`O�՗<�x�z�������e{H4!N���]��oQS���ƴ�YCa7.���uR�A cD~3p��h#�򰆺r�Xݭ�u�5��sH �n�ʷ{�4�1e�������;�� �u�q{����ŗ����3�ӿ%�<�Bkh%����-�3�#3����(��b���该�Pl|����I}5�!@��wn\(���x.S��%Z�����bTlcIG=����>E޶^Е�`����:��Z��v7&6�tJ�2�� �4�z:k�:P�Gc(�ƴM�#�x '=k�U<��o��4$�<Ү�C���i�f�f���N�2�V#n��I��[>�-�5�R����N���s���4e/����X��l�� �Uʍi����0F� +����Љ0����R��:��Dxc/Ҵ �+��P��4�8,���7^d��4�z$���C*�
�*-��-�Jm���*�1�Q5���D���gW�[�L�����ol&e��ߤ�]6 �0�\eU�/�o��<6,�JD�Xۑ+����S�fM0H��	������N�	��Vn{�#W��#<>7�d��L�T����
QX��%���I�|n&"���he�Tǎ��0�&}0�3�붓,�DM/���4 w����0����B����\�`�虀�f@�1�>p�-q���+N%r��5��9��:ҀV"$gBnoA����EUГ�\�M�|!��r��j�P�����u��8�9F�i3g�3ToY��z��vWt8g����8�Gs�� C���כ�=k!W���Y�K����(z�ʈF�i��'7��3T����(��XJ���/�?����'�"e�k�tQ�����	sk���,�h�%d�)Чm��?�;K�F��n6��)�H2S��L\��|��YTʭ���ڹUa7 J;���e`�+�E�`�<ސ>� 7g��3Dm��-S[p������*��������p��0j��"	@�~�82&��	�9jWv��ËXZ Yv�Y8*i�c%l8�>���Nh�S,�A,�+{>��~v�9)��6/�H�eŸ�$��*�h�)���T�Y�òCq%�?t�t���g�s��!��7���%�R�����7����w����Sl��vt��abF=b������&�g/�;��/(C}�i�>i=��S�*�D䑮�b�����Qm�
��7tnVu4���z�S���E'����$ڦ��ڰ5w��}�d��}͚��޲��D��� �ݓ�������e���ᒙ)�Zο��0Q��xe*��݋n"�����.2��MQjv�ch���.���=��#��>�y��=#�ZO�"A^��۴f�����[����@�rS��6��V�"ț���%�\<�� �	�|�SƓ�@�4���J�;��E�ǂ��2��g ��r�,Ǿf�%1b���^@��P.F��@ͳ���#�9����B"���z�@|!⇔�2*��� �Կdd2�φ	�]���Pxo*�;�w�H���i�A���%5q�_����i���tf�`Y�8j5-�q�4�������ɓ�PC��<�dDN�A3�W�;��~�R:tG?P��FD�n.��C�[�ڨ c��L��FY	��m!MėN�<E
�nԲ��x/l]����{���Q\G-�q!p^��'�'����!Q��l�7���՞HX�W��RL���N�3l1��=}&��*s��v��N��W��9��~a��sOi.uo�LDe���jΏJ���D)�$�_5VrF�	 MH��?�$�A�����P�cf�}�U�b�q�N㮊,�.��@�I�<��P&�P%�+
#����d���:��4�����E����Ϥ_��
X�4e�0�������.�x��/7�M^��Bvwcq�_u,y��=~�L,�<�!>i�+���-R�Zà��ʈ��M����)�^v��_��cQcYj�<Y�կ�3y�̝���wX�����r��b�f�T݅�uY�N�7�[¯f������G�[����3�������윪�+f#�w9M�=P����l�P�E����<�qF�v\uds��v��0��cRy���c�)�wy��|c����'=�F[��4@d�����,H��6ɹ��8[f��!�I �/�O� 7ŝk��>� �C�Q�"f�R�I�#r�0�H�%���3BicR_7���ل��VL�fyT�:bQ^ؠ�-4��ϋ+�7]��1���<r����+Q���o����S��N�����Z�N\HY�a/��,@ג ��_b��vZ��ߋ�Jm��yQ�O@svI�m���j���;	;��:<ȔU*I��ozHqsش�)�<�P*�̹+f�ۦ�^ţ%O���m�R�m�^���۱��(�ݗd��7��P �H�}C#;�۽d� �=(ah����J���C��n<���Q��_C����I?��ą���/qƨ�i0�c���Zq!H�x���K:�Fw���wau9N�׹Xf�u��{�r�&�~+��y87���|UT�!Ƚ�(_�TNMm�_�g��U�q�4�wK��PFp�B�0�cD��c���|��v�d!Z�Y�A��ʁR&����tۖ��x�^p�Cu���W��oX�'Ff�!P�6}Р��w�){�����a�k�F���a�V���0�� 2h�,>�� @#�uUQ�*�(A��x��5n��X6v<bXu�����!����h"�vDf���Q�4@����K��'��~����Q����='����D�n��XtY?���Q�����FU[ݽ�������
�phA�³&��[�;Ps"�z��P��.�i�	;��5�V-�(��g�)뛁���#Y
�>��R����3{�p[
�%X�F��^��G8�9���·���&�.���"��R!��G���a"�ݦ^ i���c^�O8h���uIM���o��0����6TW��v��J�K�L�u�=k(�IE���{�$/�R��>q��o�H��9�zt���S�p�!�;5��	��T>fq��/�}���I�e�0�^����6![F.X^��	�0�7s]zǈ�dl1=΁V��􂶭�ne
s3�86n���O�����0���`G��[��ٜF�k^\ Y�/�(����i�Z�*�bv$�}��rnP����`دk�~�>�]f�#����$�#9���'R�ۚ�93YϦ����_+m��Ε�j�R��\�ƭ�|��B
�x�Q2�\�K�C]��#����h��MZ�.9#*l롽z^�L��`��x���i��O�d�����ڔ�&���js�":�e"mZ�w�����|�W�F�h�b.�bE; 	Z��_U�#����׈��C**�a��x�E�����zs�"�\c���fW�*�.1���b�0�{~q�����V�����a�@��
�WF^ƃg����o�ڌ��W-�E�V��a�`WsV5ïLB���J�\�����d��:Z&!Ć���`	~��Ȓ���U�F>?��2�������W�y�.�U��
�pt���@�^7]=�P9�� *⇠Y�&��Hhp�ƤY��3>1��6��y��wJr�L2�|6F׉�1瓣]`3����8�XL��U�FT.@M��h��]XN��S+�-�Ҟ�a�,ˣ�#@L��$,�����XXL�ݏ�k�pà�FG�3%���oY�+�_�y���g��q�F3�"�	�.��������\����B(D�4{�_�~:c��ߎmѨPWqz��8�9�Q�}�C��X��ǒ�(��i��2��`�1  �ς�5P��F_��.����R�?�x?�S!�'�9kE?��P��x0�3<��E��l%��V�^7�ߊ̘������9;6��� Bx��+��܍�QR�$ˬn������\�b	ʙ:�?hB�uYk�?Q�1)x����}����D\(c�ύ3��@SkZ�(-��A@1z���R�V�,�� s�a�m(��X2P�f��1X\�4����o�IE/�$2y/�\�=�p4Qˢ\�c~�?
m�Z�F����g(G�!���^�`���'ϸQ��b��^R���Dj%�T�ji�� ���E��(�b�@j�%��q,m�hi8��ޮp}��2U�0��eE#��������9�D���_�G3�Lw������w�.'G��HR�S��_����>�?r�->:�.9�A@ k+GI�q��,��D��/�+ ��`�)�q�p�Z]Y�5V�7�m4�6&�%�x�#Ȫ<���h�ejQ�3K���t^��J��%4,,���ۜ���N�˔���/�l B�Cj�K�6Q+���l/�S�\T�ܨ�;�[ �[�ڱ�]^.��^��7[�-&! �Dڋ͘=s',p�x�Ŝ��?Vk��}��~B�0gry�疨I;J�*ʽ����A?y��>�M��F�5]���>��N����-(�RRy�Bl���I�(�{K�h��ִ��O���?�ڙ��,ԂsU�a�{�����9s��۴����mĒ���
��(}˴KWr�d$��a���k‮��%�����&��MRed�d�(�R~ƒ&>�d\����ȰE��DY��һe�7��\P����$�ʷ���(_Es'/ܥ����v���X�G��9k�Áz�K�C���:˧t���Zd��,����Ė-��ɛ)\���u_)�j4[���OZ�%���bс��ҩ"Y �|5��H�|��<0�Xx���"�|M\��S���%+ *����j餙*?����[�A"�r#�9S3�,7*�X���FdVG�Itp<���^d=Θ���n		dT��އ��UqG���C�����X��hl�m�2�[�R&���D5�<�ϴVAx9��'�v.ܛA��^�E����s���S{�>@��_�K�.۟(�Y���:�|�r�/�:?f�
�����.����TE�f?��Uߑ�o�3���!A��ﭛO���n��q;�WS�6!K����Sf}o{��	�:Ėr���Nf8c){�����˄<��(�k�gn�X5��
m��)~�i�]?�Bz���ga��}h��"\@�S�+���;�H��+.J��vNr��m�Ԛ]lk�o���)YY��η>@jY����w�kw�۶f�3.Rj����/�?�!��4�g��fHT�/tl�N�-��w7eľ�L�P��x�c#��(�h�_~,h�ރ"=f#�>D�gu�ϧm#����iTۃ���`��Ѻ��g�ŭ�T��	aCb�TGC��+��O7M���A�Y��+-՞�=:�@�lct�ӷ
d�T�!��R/?�a}��9|�S�&�c��\Ǝ���mDlN	��s&��em����LCx	��azU���mȵ|A4F �>W�p���!&�r�������|U��"T������t�3F�Dd�xN8���M�Z�c鯝��s@�'=Y��3�E"���=王~0R�����5 3�} ��Ae���ư�8VcQ�b��`�l����&ٟ� #o	`���é=@z� �i����-�ގ�'μs23~�c�����1���H.1g�ޕ����������i�-�
�3�B��C�Bc�����2��<��{�W#�PÌ=ZV�t��I�5�Wo��;��&��.�Z��V��h��3;�t�p��Z�Z0��&�6_R/@sǜd�w<Z�[�Q��k"�J��!���iq�"���r�!�|*I2]�?w�|V������yG/q5�u݋<��"z���I�72@. �^H��P�cA��/��n��D��Vj���@�|�K3�hO�T5S�N�a�í}�c@�[ԕMI��O��|T5f���_�	�P��|{Ϋw��VvV ���"���T���ZGx�7�����Gvy�s߶���[;��B�[y��徃��f��YJ4����y��ut�h�d���5u��^�5P�19�S�
�C��R�_���9D.��ڔk��!�"���%ʖ��gq`�lߤ�&��w��zXPl��+����Sx0��_(Ӏg��B��'��K0��F��S}>��=�F&�\�/�g<����QP�!�� ��h�&=fU~��{0�+,����k��B���Ļc\��y�06��%�O���<c�ψ�X�\�z@M�j<�+ o��n.����^~y�`t�l�_&oJ�*���<�*L��I(��S��#���E-˛�*�`���� ;u�m4:o�K&�!�e�Ui�j�}���*S.��Y笮����: M��
�>{}0�܌�o4j�M���dB����Oz�V��n�
�\Z�5h8��y�Ĺ���i�������)"�tx|	(��9F8���r�w��>I־�C�3��ȱMp��)8�*�a��h68<	��>��e���4F�x��E֙���I�g�
Y$��$7Y�����1��M��������ܦ�;;��
d�AW�Z�ucX��������Sˏ�2��&�Ev�Q`i]�B��7�@ҷq����N�գ$$����)�����q�koy��z�����KT�S�^|�cK󉌎�YF	pl��C���+�MG?�Y��_�{��+>�����!���[�����O#>�
~CMW�҂�z�/:5�|���T�t#)��>\�;)�8X*5����*s ���%[�~`V�R�,W��D����V�`�B�N^ބ��2��:�B1W&Vb���7�t��7z�-2q4n%A���Y���g�l�߶��3�Y�2d��6��DB~ٻ�E��(�	-�D�q�h���.�%���!i��d���U���_e�0��ʾ_��#���0�;�a�����Q�8r��⹏��.^�e}W0�>M,��<ҵ,�"��G��z}Q�6yg�L̚�� h����-��5t��n��T都ւ��-�T�Q���C�Vb�X�O-�oGX���a(��XS�%����-p�Y�Q�̧(���J�S�#�/����?�o��B�wOe �g {���hN��L�qX�Ү���%�Qv��o��B�#�>��6�vT�"����v�]�d��gL�^�{g�ܽ�%�e�$�� +hƿH"�[�a����RHx����y��S�5 5Z(ʋA��H��Jv�[6�8SS����4�5�j����v�oK���M��ρ(X��n�1��aȮsg��W*�ZD�H,R�(���re�����![E��ׅ���*�/�85�H�)�:pp���
a�sOڟ@)��y�s�Yc��sehn��4To���f�j/Y٦��?).L���@���K����>�n�<��1i�)!��}lO�oy�,(�qP��pavH���T(���
��"~���w�zH�oZ��P�׍)-��It�����Fh��{��N�4X鬐Tm_��%|Gq�Y}	L�z�#|��'B1ށ��k�����78�Zz��ֶ8���P;B0��:t�b�.�@�PmK�?@��_1��+!�*@\UY�3�"��eD���|��oKO��R�zRH�S���?�Nm�������o�a�m����`Ff��s�؜	e�O�tZT�){m�C�} {��
�ZB�${�b�i�$�4�@�x���K1^���"�Bf�s�\�D�2w�C��(��ϼ�+oZZ!�J���t��p�������G��!�y����+�f���� ~�4tXj�x�!��>�����|u��C�n���ϙ�����#%�i�B�j�p�oԣ6H����vLy��R���^p���g �1�"�|���i�$��>���&	Ye����`��cJl�u�d$�_N�5��f�˿m�bޠ�Hj�o�i�*�9��(* �f��+Ш7~`6���J�����Qʴ�#�灵�X"Y肬#'ûz�P��!x�x�b��+�ns���k�N^��K�7o$�T��q�����?u��f;�)��0�(��A�<Z4Hv�}����+;�L,#2+t��Ƭ��1��z�P�Q���<�O��oY�=�����1.
O}/95�j�:���w�B{�n�Ղ������\7|���@'|�"��!a�q�r�>w9��j����K��[x(�"�����?��za�ٞ��=2�� $���k�!r3���c����,�݉��Ka\ll�p�<\�G�p,�sì�.�Zhu&i�[���V��E��,/I6�=���;�tӪV�F\3���SZ���r��+G� %���3��(�v�T](@��D@����A�Kٰ/߯G7��x���Ja'���V|�9mV'�5�߭�;�"έw��m��#cю #�J,9�d���7�G#����I�2�^��ރ��}$��-�T	�Mo���6�٘8������|�i�:�b���`E���-����o?tyf���<��B����K�^�mG%�x3��$T�p��] x�l p6��sy��5�':�FTc�Y��3�#T������ )��0R`��xAT�)�沌)Qư'�{t|����m�;�$l��mz
���S�d�>�c`�yUd�BH�𠈱��?�d�t[��{�f�r	�G4���s�u�]��k���r]�4���mb��<�Q�r&����
�	A�-���k�1����H����фq@�<����Q��!:k��w[9_�m}4�� gq�G�>[��=�
0*��k�fgJ��,��i��͎�=ڠ	#"X݁]���bQ��$^��^ �V+K���$�ҿ�}����0s-��vo-�������;pLx�v��BIȌ3�0�z�5L���H��^��k��6���Zٰ��!p�J��r�j��|#
M{��'�u�R�2���aHg��1�����h�o	g�]2��Zc�)i��Ŭ���]�`�xv�k�����ۖ�?I3
�Ls�����k�@�΀�M!�A��p�\NU'�[�ųK\k=�����H����/JJ��^�*7/S�}ߦ
_�OK:yi�<�K�s�$ ڬHO�c�l�h�u�������ӭ=���t��.�.���'LMS֗�*�ě���!�g�P0x�� B:q@��Pˀ�c�6�_���]ڼ�z��S'�xok|�}�4e�;�
7���hH��O�0%b�Ӛ�L��U[�Y�e�ܞxԭ��A���N���*�.���cD�-�A��Hrr�D�(��V2"�d����YA)蒩�wlh�Cv��/y�Ħ�v	y�����nД�Q�ڡѢ�jre��|^���\��l�{��OёQ��̵�9�l�Ae����d���r���������`Z�:�u<�-n�|Z��]����d��T�z�l��kOP���7��HI#NGW�T_��L`����K�AF39�g������Y~�R�~#�g���_O`<('S1��Lk��.��g}tSiZ��F�,y���,~e �5g{�՗��Y��ߵO�C�Kc��iD_3��ח'4��$��Y?29�ė���3���)������ݛ��
׎�rlӑo�Sܗȳ�G����o�I �]=�>���j�}�ƹP������'d��.4��})Z���N���P�ׅ���U�f�'��7���e�ڠ���XB�S8t_t0�π��!�y�)���yE�نTy�E�2��ĢQY���O6���iF�]�Y�"�"�/�T:�e�5�P^Qb$�<��	YT�I2/�lDGE����5QYU��6Q%&��?M{r��t�f���������_�0�$g�e����wܟ�@���!��4q�p����%��h�`!|�g��:U��������IO�6!��X�:i&ݐM6}%�*�IL�u���*���:� A!l-X6.�@z�u{��ϡo4殮ն��?�����Ǩ��f�E�������iل�-�)K�d�^r(�e��g/3�G]��U��H�k֟�a��C��h�S
�ĵ�ղ)�M�NA�-[���b���;����83/��G�E�f՜X��p���~���A"[w(ؽ��Zb�B7�-��Q��9�
08J♑�u�-�]���dg[�pWP�<�md�#�|���S�.IBlv�����ʔI4Ԕg�N7h�2�3��qt�g��a�j����,���K�'���m��!�Jv2˵_�|~�8���9��j�|��� {Z�+�8���}�cظ���uY!C��!C�P���� g�S�+}���om���uϭl"� �U{ ��tz����$��l��r���uj��`o��s\����=z|=u'��L��{��� ��B7�I���gB��A4 ��BA}!1��6g�Az0���F7<��`����3^;�K\B	�bl�bn��p��t�>����e>1ȉ�:\�����#�y�1��_C���I$��ĵ���؜�뷙Q ����-U�9j���O7�	�Ryv���5� t�k�����ς?�r�"�
�ì{)$�r2|�rw�z��V��`E�<���~�| �7Ch �37˃��4��w
'���Fw�۬��|�#*�gt�P��#��Dr##BUU�j\��F�7���	�_O���X��b������AZX�����wؖL1�ۺB��-O��Sr+�ڀL<Լ���\u�ݣ*R��*�Hn1�顁�a���§�$�@�Wl
_r�<MMBv���	U��_�*e�wxķ�,�"4�_��)�N�3q��ok�����f�8� SLc��\��'C�o���7��g�k-���,�Q"B��	�����D�^_�S��!����NN�����h�[]h�]��vD�N�c�Ażr��"�4} @��џ�l�����&�g}r�B���-�� H�Ƭ�F@W�DH5�܉��"[Y�V.�b��M���K�s3��⑧��E��L]{�'�{];�a�pb�h�s(xԏR��6h�a����^���$��U1y��+��J|�Vߛ5��m��ҁ���8�=	��$
6�+t�F�*�^����=�Q����w�?���ϭ�;��v�qY�!����^9�U~U��5,�Z	��dFش�M���1w�Ծ�Gb	(t���d�ah��8b��G�"� �����ߧg�R�?M�x��g��vHк���!Q<��lou���NO�66 �~�}���N�0�Kݯ*}�6ng�Qm��aO�tv/�>�� �u�$(Y [��h.���U�� ۽�j�;�p���P:���XW	�^h�;�L����]N�������S��iP,���9ׄ3� қ�.���䋾��7���͑�R���@gE�}�:r���(�.��A�[���
"��(Ō����N:C3"����ɷ���%;_�kvJ��=��(��܏����=���t z�¯Ƿ������H�'j�Sk��~^���u�}h����~fj�g�Vf�p���WgC�����H�tLn��u��%�4�^O{�c��^���<�o�e���r;�z쭟N��Q�ρo��C��EA��i����=�m�_�� &�6�Ó ц{cH�l�>�4�m��,��8� P�%��nGoU�Nv�XR��%���M(N�x���9� _��>���)ԛ��5�@!�ߙ��=AwH��2���y>nxA�A�M�P}�a�8�+N$��\�`+��U��
�&���Ωs��Vͺ{��e�E�K��K;��3U��%c��/�����ٟ{��I����>s=������V|��"��^�Q�O��[��a�#�)>·
�ۨ/
y����t����#-�����^�PV��a��7�D��MQn�"K�P n�پ��%q���gS����� |ׅ̑������D�4)MG�7i0ć"�0Y� ���]�*�g,��Ӡc���"���:��Fʧt`{v#q�ce��r!�' g���r�ˊ�06<�S0;�J�O�ڪ�fT�M���� �	�9j���R�{$Mo����o)�m@�K�!=��U7ˉ�R�*�)��d5�o����W��
�D`p�dC���{��0%ɛ�x,��$����S�p�y�|�����)E��0����b����s��x� +���-��>����ߦ����]�TB���1��=�4!��<�V

�$�هOi��"���.����鴎hfY܌>R�����`��2#��9�����,� ��Z�\�VfC�br4��x��<	������J���V�c��g����*�
�Z�ubi����1O��6B�W

ǃ*���ۆ�Y4I�����*�O�vP�VQ�6?�ނ�:=��_tG���A�=F,
��S�=*�2�VB�����i���nR�ĕ6i�p�L˕{^e	�IkFVo4LP���q����p8h�B��WaiD�N�8�>����=.�(���P�f �A<JQ��o��̶��5�BN�п}���hw�tw���`m�0j�AI���{Ia|N�v2�"�S,u�K u�D�������|	^V�[ʜ��a-�"��ai/���������}�s��?�������#Q�O"�V.�sy�`\u܍&�[
�6��nm]��_N$�z�oY�H���mǂ|m^v�wo��IT���p�4d��gt���`\2H@�j���Ĭ��!��T	3�bT1��%C��<Pz�� �Q��+���"P�n����.�d��0�T�_N_�g�����%��8��9N#����DV k��ԓ��~�����d�|j����W�c�ԇy��ia���� �k��C=���C�.�%X�[e�aH�'i{tzDF��/�Si��KU=R�����z&��Qj�,���v�k�uH��u��KF1d��Z��N���7��.Z�h9dvJ\�_��O�l)������&\���ο�ʐ�u�PGMݔ#�ߕj����f�y�3�Q�.u9tv�SC!�_8�ތe�HG�������ڨ���kJ�����C�²"�G܆�*�oGo�M�@�A�rO�sluz�C��tƮ��d�D{�aqΆ?�j3}=0V�	���#�kQ�z��\��S.њ�W��֤o@��Çg�QpLr}��G���j)�t�E�� ��zi-������)�=R�v`hl(�jy�1�	-�����㸕�|&Zh��֑N�2]{�y����H�Kv����D��Y�������OH��g�Id���s���s�n��)��x-�f���U��r�o�+E�'�R6=��*��6P�PE�"�"ۧpw�i��6被A�S<F=��wfZ˂��u������^)sl�n��	���:���*���©��Nh�㍏�����i<�o�i$�3Ζ���Y��1m�T�\�D�nɂY59:��.�D�����@��|G�ᵺ*�@��Þ�Uq�Dв����$|��	\����0懩V@!��ZSX���b0��o8]Ir#Q�)/>U��eW	%�����M��~��<��B���n�%��sرO����;��k��Ղ��ۺWN8}1�����:�����y�l9��?�h�
�����N���!�|YL�"1գ��H��� ���&�{W	OC�tH�*�68#�yDfvae��Nw|fzP��D���-�s���R�:��tt�9�ё�̹�,�|�
ccʼ�S���V��頚a΀�0
�{���
���к�)u�y�he�ɂE��Wp`zG�1˼��#g�v����_,���sfW��xh������:r�k�g�3���A��B)�G��x)Na*Mr�Ko��������.�p��G��]�vl��=]�"�.�
��ƪ�؃�_���]�;�ɥ��(D�ԥst���4��P��: ��EP���C&A���~�8c��|�
G���N��)�ӑ$k茯F�#�C���}�l�!���s|U|bej}�R��(-�R�d!�|��M��,R:S:D�Y�(!;A���k>����-�����?��?�l1�T�r�&X�9H�ǁ��Ӿ���z�g�[$����7�浦b̎J=���V1\a���IV�.�fy
�3��B�.t2^
��8�- ̬n�QO�/���$v�5 �Z�ke>��aP����m�ݰ;z�>$H@����`ZM�\W����D<���_�H*��D�ht�<�UL�6�Kgf�q��gD|1�&� �����k�����wΚ��8 )q���e>�3d\꼅�~x�������v�?̡�X1c\�~k�D�1�fc��y�*���օon�Y@�7��TO<ZNH��C%8]O�{��V+A6do_Fx S�"s���ũ<
�+ǌ��o:n�����}E6�����˽���U �z��L�^�ԵY1|4�a��7)��M��F��� ���3��4�ݲ�ۯ���q�}����!���4�n	ƹ��Y�dBo�p��k��o�6'H@��x�	F+gS�דPe�(W��	�,����A��s�8��F���j��TCSD��ˠ�כ\+S�>�����8Ǆ&�w#��5��@M�6�蚞��ѵJ����C�=�5(7����S�F�aV_3���[���S4vX�Ӆ p<-�e�i[D�n���<kS#��A��񥇈�A3�(T7
B��	Yh��+B�XT2����镓��/�,�����j#R��YdE��UM�\�5;CYH��+�J1 ������|KA�������&W�i
ı�|�׺O#�M����)��e	�Ӊ��a�9=�`�b�i���Eţ	'l��ts����Q��WTJ��)ޚ��pP��N�2����w����0t���I�*U��l�OM��X�7sF��mlʋ��J F�A��82F%��)���A���(B~1�v�y���}��|����e�mx���~����,�2p4''G��YK��̎Q���|�X����>_+���=W*����͠��D�\9��C�M4�<kw�{?����_��>l�������c@�L�Q�������5u7����&c��jdCΡ�(lD~�U5v-Ts+�C�rY�T��%��~M���n^]�1��n�E��f]�:KΙ�a-gL�Z��
�&�{��F��xc����"��I���>���&��Aa��;f	��4� ���k�CZ��/�=��!�GU0��M��֎p��6���)���@���\tUjP�Mgq�e�{�CE�"�39�L
���Ex��U�����7�A��7�� g�"*4z��qK]I4���`BĬ�Y�ȼ����ć�պ7��ō�[u��z"�.L�I	cb*KyĜ��6.�a0�c�|�j�H*��$�/�C��gG&���W��ja����;�W���������^MdY��JD��^��.�8��4E�e�zG9�H�{�5Cg����My����J�2����n3:d��o��[����Յ��ӣ�Ҙ��X���i
3�<
���󜿋`�haL�����k7��B��E/�(͓k/q�~�f���\�Yň4ŅM��7�r'_Fj�!���eP��<x�]<�+r���#�I�`�o�X�F�ΖSa�����ք�ԑ��r}�s��*�{��t&��r�x�l������c�[@�nIr��s#+)�w�/�_Q'1�v�usa4��<�_I$���缍���W���묐S���`��`���i	�05{��4�e��j����Q���GV��dbSqK�&�J��r�ے��!'�G����^+����������T��$���єL�����n�8��o:��d."�˛|��˔&C�)T��Z�U���-���)�P9�����Q�폎��D��D%
�U����Fzje?9>)/��qF��â@L�}e���O\O!���<�:�n�5�E�h����AU@�G�̟��bb;��sP��C]w|�"���͇s��<0#U]�E#l��Q�5V�� 3�wg}��=q:Ǚ��յ�������[�&�J3���!�HOtb�H�/��v3����(n׍Ki�i�֑�,߿N�p��'�~��)V��(����rM	�	��F���1l	+N��Re�N=�(Z�|�:�M��	�^�a�X�y�dcSw2�Y�� 4��4�c�$$�%��?��L��ٟ���Xj?��l�(U���(���9S_��T�^W�ή��CV-yk�ʥ���<���b�I��(��o�G��j���E��r�%��t��0��6)��<�Z���-��\�e��|��5��O�!��I��������d#x����+���!"�7�@�pBWy�&&0�<�M�gV�gJ�@(������|�Ղ��O�+.�:��}|2?��\���5���)w�A�רK�7�H�Q�y�S�]�5�8��	L�1E_����b\����g�zs��]���tf�I�����f��ZH�{-�<f.��X`F��B���Q�_����O*f��6y�Sd�G���Ou�w�ƽ?;ɶ�����#?AU3,��܃v��|��,*d&%{"�� ��RtfB�"����r	 $\İ�)�m* ��׋�aWuF��p-��2P͆[��Jm���ԟn��m�=/J=|<mm�Ԃ}��;:Q��+���W�R��Fi�>�KU�\�'�a{����u���H�)��d ������|����aFdgM����!��{c�0��	g��ըEu[����LY�#��߽��L�"��Ԑi�?��ݓ"� ��A��l
�Ѕ�v��Tb��@�X����T���2�I/9��F�t�G��Fo䙗�`�m��.�_������Yr�t�gp4<od�z�$jn0���O��ZP�J[Q0�=j�vF,D��}DS�i%29�W���;>ݝG�N!.��t"�o�*�@(nȷ�\�����î?]�!;��[]U�3=#����S��w�Pĭ�,����_5��әQc��6xJQ�-j���S���Rl~��9"�(�7�ɛTZ>#��{F>[�7�GC�� ���ZK�z�֢!��>#%}R�i�sj� ��K�az�D��&]�� H���w�4J�����)5�V�ӳDU����������~<dz\=�ߌƶI�W#Pv�*����@�F��K�`�򹂗���W0�Z`�]�P<t _*V_�ȅn��w!E����؜�rG�����Y�V}��q3��-v����Ꙩe�*۳�2K��p��<��3o�@���I����VFJÃ�eڑq�lf�i0z�}��;	�=ê��[���"���z���R��x5�A����ẐF
@��U���)�df38s(0���� (3���O���<nwbێ�`��ɯ��v�� z�|��%S�t�nO/���7iA���1�OɊOj�A�� 5zq��ed��٪�`�
�Qq�H.��=�/�OÓi�op���v�c���%9�c���G�"���^�Q�Pk�B�o��[�����R��#^���:?I��X]�t�1)�z${�"4&�4�h�3���l�q#f�l��LT��u�_�	�r�,�����-Ke��#�$|�ړ�,9�]�C����!ػ6"j�fB������BqA�Ns�/:�ˁc�d��;�|��Q�D�����ڈ垘�Fn�`����s1�,+�	�?zCla�k�������\��w5|��0uG�8H�h��	SNׁ4����G�}���ث��Lts��&{� �|i���'3���貏㑒0q���?1����2���/HNu`uc3�]��!5Þ�o3q��泰��s���:�9[���sYl*�q��/L&��� f��F�H�y�*k�c�w-��W1�k�ҿ��e���J��+��c���i�̓��cO\9fg���e�揮IO�$t^�H̺ h	yp�c9��D}�P��� ��i����}a�����AS�DE0�9��l��B?8��D;��3a��,	C�M����Q2�����j�0�g�7�H��n��L(,I^�b�c~8��N�����7���R)����,��w.'>y㺲XS\$���=�����`;��z�s`>��}Կا)a��ܕ�dEa����;E÷ޏ�WR�l�MG��X�j�E} ���������2���J��3��s��W���V$}�`�x*�MHx���'�u�҇B0���9��K^0��a��]'�r�rm��<Y|!����@�/��U�9F 9�Fך����n�[@`�
��V�n��~_�5f�g���ag@�a�agG�X��w7K2(���3{Iz����v�:Ԉ�S��ï52�(囧E%\x��e�I|����]S�H�p�4~C�)6�S*�B7y��>�sd՟� hM�ވ�.+f(��\n���l��t=����Mp�ՙ;Ÿ�]$񠯇�j�hR��N�p9�����E��ם_
���E^���ήc�~�Wu�`�GU�H.HY����a
��'��#��D`U4����=o^%�3��պ��ؔT7��"dm��wa�M�g��K� ��x[⾠%�̀��o��\Q�I	��wWƒ���v�L[�ʧx��v.P�g���܆dw ��
�J��|0���]���7(��>6iv<^�f
w�����W��4��ڔn3�����Fz�W�ɝ7p�NTG��5����̗a�]\�.���H�/�xۮ���2��>?vw�r�R���QQ3K�4�����&fS7��4�����0׌}�Y|��/-bސ}eR�d�"��m�0_�[M*o< �]�k�vjPy+�
ܨ�H<f��f 8X|���*4 ����
R<[��u)O�Qv�i�Wӣ�RO�����c�󜶨�v���O�/~�]���1�е�����T˖�P/j,���y��v�c���wTG
Q?�I��t�܍�&�u���Yy��{��)��+�#�H���G�n�J�nP��[��k=+�_k��%�2ХN	�
M���m�bX7x���t�u,�c386z��NP�vr���'PNY��:9
��ɼ&�
ģ�R�e��`u��ͯn�(�n��WgF(ت����F4�C,;��4����Bd���j���Dd,ŃI�V���b��������}3��c�#�GZ݉�e|'^K�$"1�Ǔ[AT;5��ɬHfH�tm!��[!���*�GZ��B�o�[p��cQ��wѰ�;O��<lr��� c�J2rDQd��.9YΤ�`ӻZ0BG�ӆ��w�},+r���ߖ������M(؊ő���9"��9���sl��Cj��4�QB�q!���=;l[�(M;:��@d"�%~��;�"�(d�w����2�+	����%t�Mx�8��F��0�Rgw�D`���Ȼ٤� k�5�#�x�QQ�J�kh��MzJ��c�v��.�k���$�Ҵ6V�_��)���=ٷ�.����d[�����:e%�@ñ�cP�D���
8��N���ԍ&"�#+#�A��K*��ε������u�y�?μ��͸Iʗ�zg�Ж�C� 0��[�br�n.�NfI�=��		�6N}�89ċ��m��)�z��
!��az%$����[mK�s<}�._��=�M8!k�ݸ_ݨfH���t	8���,�$]Ĝ"|�T]�C{D(I#|q� ��gz����e��ţ��̀�zJ`�vG�YxԺ!Y�"Xb+�d)���1�C����h�-�y�nE*?Xü;�S׭�{�i��f6ð�+w8��ac � �V����q|���40�s~� �;BB#Vc=S܆$PmL�;R=�E����x�"�R\�����6����y�N��.Q��A�v}�47nn�/�#���	�;}�c����gGi|��s��Ekqx��������X��q���a�^�:��Ҙwqm^rx̜���� �9��$;�,�n��x3h�~��np)f9�k ����-�xP=�N1�x���5�n����K�s33��&������_�J9ʣ��Z�䭦�����T���"tz��fl���̵�YSԴ�)��;J�p�	��[nx����8����o�'>8���;����D�p`�fTuܒ4�=5T� �R���,z��./yk�E��Q�i�W:���X,{��)x��d����,�x�����/��� ѱ �g�Sp^�#R��i�%��h���qr2�<�EWW	3�A����K��_���G��� ��XDs��1���$8���R���@)x"���+�C���bL����mW�?�=�yy�PU&��P�Z�\� ���♢	A$�������������c��g���x�Y;�%g��N���'����w~�lp���(��/A���C���A_�.��A�0�9���8��Ը,+�NH�+	�$�?���%N�a���C�مݐ\T0$h�:�sC'�w��H^���ƪKw�y%�\K�J���,�U���rz�$X	q�5&5[��ۗ�,-�g͙yy�6��F��>��d���.V����X�b�t��&�0qm7��}P�������{������Y �H��X�H�����q+�R�Bp�)XM
>�������eDUi�˦�1�P5���̡����o��V�Qݢ�	r���R���P���N�B}�	����Q^PA�r�=��N�x�Pڒ=c �� p��,�-9��[r�?�N�OۺO�gK&U�#l��6tpB8H��6�E\^(ڢB
�B47��,��>-���Q��}*%��><B��|�d�9��Yǭ�_��;}^�������4���a¬`elw!���l�ڽ�)愓tT�������쉣�����7_�7�c/� �ˬY66���pl��l��YG:ES�H�偪����\�sB��f]���/��Y�U�`xx5�lyS�S�W�΀=�s�Z@�w�)��a!��L ���EG�	Ā��`���o�uD�f�1[����\�n ~�o����B4��	�ѼG�҃��-���}e�=�~����_���N P�H�)���
��w:�y���胋Fձ#�L�@̷�?!w 
�V9`~m�e�3tj�>�&m��--�_����mNf c�O�����I�@��?����B?�5Z!�R��s��=;I'GN)�F��V>����v�"�^���]�AZ��IO
�y�B��m�6X�'���,4�U\|ɮqy-�Dq\��������� d�=.��!txn��$��&>����#|}P�G�=3���+���x<G�fUa
`��e�t��~QQ�~�5Xm=F��s	s������m ��LC�Q������<�BKg=pm���UaPB-��m?�LV*H��-�� ��Ch� :�����ƞTC�u��Ŝ/���W���YK����^S� >{8n����d]y2:Fp p�w�`��{4$�)D
�T�q�3#܇�"4��h�����'���G�;�<�1���b5�hx��RK�k˼^���I��v�u��<(Dݷ�|P�v@�j��Z�'���G�&�z$�l�����EB=t"[Z�2���+��G�١��Ъ�8�<0k}��H�+Sw�*�=�e� ���v���k����>s�U�숇�<�u/E��f�u�F�,%�:nA̡�3*�PՅ�4��:�u/���tS�X{\�Ֆ������~W$l�㌷��-N�/�@�q�8�z����Ȟz���m��'��c����|��k,��z�j��#6��p�$�pJ�%O�d�kty;�X8O��7|�L�g������O��a��L�D����URll�&-�'�?�C  .IKp:%e�1V�
'>�j,�6=���ΚM5�V�}2 '��qGT
ʰ�]rb68��CҾ?�γZe��
6��j����b$�D��-�F���I��/�����@��C��y^	�~K�c'Z�7�7F��7���5������A�K
���vt ��������X��ʋ!���.�����Ƒ~�j� �9G������߽Q�6j�`��]ַ�.��L@�z�݇����rזF��J$�E7��O*m�fgb��*�����M���"�Є�kHK�Y�~{ui]1y�m�Tn
�3�Xw-X;ő/��`-�uro3�S%6"p�j=��ƭ���n�Tb�hU�Y�)Ǝ(j�7<���pۇʖ˿��oX?=����=�?n��V��
y��ϲxw��R��1�λz{�W`�-3u3�iV�Jr�����n^�=	sLx�-�q׈兩��-Bݖ���un�k�s8z��d��6��q�G�;�Լ�]�����<5& ;^l�;���_z�*V�1�k1/7�2��z/���a�g�	G0gw��=�or�u���ӹ��55<�Ne3	��Y�ܖw�����E�F�����řލ`m6�v?7F:��&��s��Y�Sܮ��P�����uo��w\��S�Վ���-d��h�X�\�o���R]�A�q��һ?��/�����xO��+ ��g
��9 E�'��[�ںI �"qX��-"�m��L�����a%>� �����6$���Z��O
�<���>Bt��]�ü����?kt�g'İ��ܗ�F��+��y�a��	h:���t�j�n5���ɷ�E����v�� m��X>��3����I�� w%� �L����(F!�
{�
�؉@C�������ji�`3�b~wG:|�N1"ޖ����.��5W4-FgyVfzv���.dg;�?`SJ�nF���� �N�̌�e�2j�X9�k�卞�:�FۊU���8w�8 ��"�J���T�����ց�������QQ��8 �&V�s���܁oD�
	פ�)���Q���ܖ�gP��_-��Q\�,wꋀ_O��W���	�G����qN�z�sͮiN��B��Ia���W�|��Уt����Zթ����3��T�b��\6��wT��7�	�I�(�&�|SEa9�ظ!}����G�;L��~�ԙ�u��0���^�MS����ƆK
���lGo�����{g�E*�;V�� �֢$�g-G���Rtf�\ѣ9�gDC��Ɨm��eAt� �~Ѥk�"z�eW�$j4(��A�p�/�%��}9��xx�{!��O̫�\Az�6D(r�ӳ=�C�'u`'���\��~K�(	� A?D��UGJ�ĳ=�S��7�)B����OvHA����q�>�<v?(0�	ɻt���vQ���D(?��ad�Q�ܜ/;/%����3��\Y��TH������ ��J0; sw��|S��N5�r~G�~�np����QD���i��kM���.�����#\�?�i��� �vY)My6_��6��M�Ҧ���{�tW��`�%�^E5�貀�xH��;$p�vZ�<������*��������~='oFR��u��.Rɟ�L��HB�b=���Al㐄}%�a/(�պ��\�	{��f���ChV�^Gd����ދ��#���{Ѡ�=�B]�#p�	�.���GӇ�`_"�U��F~�'�ҧ!��R`�:� �l��L�0bH�t2(�|�Q���>�`���D8@�)C��̐��>��w����S��)�%i�j7���B�#�+h(M-�b	I��@����+^�8pX�)���ߊ�
���Jw��Ф�Wđ�<Y����EAO�	J�CuJ�	��,�V~7��}�/�a�����=�ͼ��B��\:���	�/�D��B�����7[1�4u����'�l��O%��x;K�[�C,1p���Z!��0Y����؞����R� )� fos$&��Y��O��(�{�r������~���(�hyDFEh� )�Z"�i������y00�g9w��`=�{=qY�Ф4�ۡ5u���*�:���''hx767K��S]Iѐ
��xJt�B=fLF�1$L{�fn����x�L��Q�L������b�3��a4K�ȪrS�>���$�k�W��Qt�� �K���C����&�q�����2}�e�k�3�5)�!�/�k[-X��@}�̾��(��e|`���k\'17�����|�Pw�3�^W�L��L��#a�R�]o�]d�A�EQp;�~ciǞ{݁1*�n�3���s�"|��q���q�Ɒ��50��O�ˌM��g��_��c��DQ�7|��.J�@�����!������7�A� �z56��9�y��GՔ��tu�w���M�e�A�w�p�Cn��@��������a}���3<T�Z4o~���\��������èh>T6�=F��{C'C�X�����l�b�e��y�<O�����c��&�2rC}�1�aR��[�t�0�� �$�C�]�xM�5���T��_��ز~����eCЈЄ8���o����9�`\&�M����02w�.��%ߜ���T�mſ����	+��{��>2+O5\�hפ�� �)�8Ut�n�?W�f�r���Tv���cPj��{�k:57��p�2��`m7��h��t�.�L�(GW�Ɉ~&/�@x*��B��7�� hٟ0Z�q��I}Mu�ra�a  7���%k��͸�wl��%���~��gN`�tص�N|�B�~�x.xN4�a8s��c��X��.f����OOH�92t��A���_BFf>���\���i��O;Ps\����x5gF����*O�I��x�7�f��
���jl\Q���A$+M��Ki�#�bogcb����e"��|u�(K���Cx��^>n����+X�P����~(>���� c�i6��:.�f?���K�r����	�惬��l�]�������5��T��r�<ïel�5G��ښj���qUVp.����e�e�1'Y��o	l����Jv�.��ˇg�JD���$��|GHp��u����7��03?� ��]�+M?AV�6YU(�坡{	Ɔ��s3���f���lOE�y�<�v%Ң��5 I��q�s������	@l���g2�?�������F���;0Qլ03��B\�ſ+��#j�A*�'w�:�;i�h�'��o���>ZO��4��ml|s=�A�9�&�>X�-ۈ�7�� �����/�� ��ѵ���?�V�nϼ;��7ʽ'&�%��z�Y��U��}�%U)��n:��t2GFlrqy玪fE�+6;��跑ς�Y�W8-��0n���LS��������]�7�����#q��UU�$���b�����X�(��=��6N���&��ݵQP�Ol[���w����f��l�3;���|T��AS�D�n_?�+W&�mhU2o��^�>%
�V�VI�s�Hz���r2d��UPx_`��׾�F���Nu0A�a��|c�x$[��R��PJ�Ŧ�+��	!�_/J+�"��+J�rq���;�4o%)2Q
�{tkE:@���|�7nPՓd}ټ�le��Y{Ϝ�p�"�漈�E11�Mf@{$������+�A̖���$�|�C�����T��_����,���Od",�&���1�t�h-�'�{0�'�X\�n���2b���N7��=Xm�PX�P�gh�>�0�B����	��͉P�fB����V��㋀!�=��`��1�G���}�UT#Չ9vM�@L�a�>��p#�(P���Xl���(/CY�SŽ��XR�x��D)�ҡ�g\��W/���?lI�9��{BUNh.�߃Ә ��dP.�I|�`����Y׶�����"ĥ������wKPu6���S�x���6�8�q�-�'uyNV���c��W�nm؁b�ťŨ&�(�{]���i9NjoM��6,x�ڻ���9���f͋�����9n��<��&]���>}�&y���}n��@���ת��QoƜ4���l��5��nQ�#��J8�޺���y��;$m=�P�
�/�Ɔ]\Qׄ�+���F�1kDW�=�����8T�Q|_l.d�]�bLad.R�͔ɢǬ�]�sWb"	�,�53�US�uI��tZD|iQ��x�/�~��Rh��,}2�,>J~�ұu�E���D5�u�%���@�������1��� *������7JT}X=�����i�Jǂ�Pb� ]O����l���H�yL9>��8����l�7�K�=LC�9jx��oTl�����.z��"UVЉ�ƥ��o��N`��y�e�_�K_�1x�N[��R��6@�?��Vb���s���Y��V�ui��L�[QG\7F,g��jؼ�6�ڷI��C�Oq�B���U{�)0b�7ԅ ���V@gK����$֥�N5)�_l�$[��HX4\�A0(ߘ����m�o05Ω@WN8b.t��4�����L�&?�ز�%��o?KQ�<��A2V^L�R#�޺��T�2�,�97�P3��V�l܎I9�$��Q�DE�UZ�Lʾq;RUW':�v�EVd1T���hhU����zUIAqh���GI��^	�ӥSYsj[�I'�o��A�A���5z鄠�Ty؇�������W)�y�ӊ &A�k�V���#~B�~��J׶s�^��Τ�3����1�U���2�`���zZl"yGAK���<��)}���b��&5Ǎ������m�j��xߝ��(��W�g@W��^ҷK3��`Wﻤ*A��D�S�LE�3u��eI�!dm��v}"i� &�T1��GF��IR�VQ�Ĥ,����}���<k��.
,���l��['��d����*���	�=�Q��?k� 5�J������m}ΪDS@�P�P1�����]d�e�Cs�t��%�B�X0�=��r�Q�ď꩞����@"~y�)nYB�d$u������K�=�*���I$� �CI�20�a�;iR�+s]ݡ�/�ѷM��O��CS��0,#%*���U���KAF<�����m������#�qi�#��4���q/fޮ�I2�m
5����`�	�Ľ�GI1ʧFR�dP��&�F�6����6W��r�ƚuP�7�/��? f�Hʊ���^bw3����}$�^�|S^apv�FMh�h�I������[;��BoA�{��6���E�������u!@9�_P��q�@�^���9���~�Z����hg��C=<��ʥ��2p�eJ�3W��UD��Ė��F8l�M���3�����*򲺧V"wt���W	g�S�����Π�K��0p��̖㒖���n������O�ތZ}~[�j��h�g� B;��5dD���S��񿡧���_и*� )f������8b�9&#ߺ�B	��;�}K>J�M	���DO_(.�՝��P��`�� s��V��ܥ��nś�B���W�$2]:���/Pԯ�s6��ǅ�F����K�?��p0=ӾPy.%�~�֡�A4q~<;yo��,!���9���CؔF�}����`N&o�N2�e�L����������!�����MQL)�����#���B͝�r��R�?���\�L(��&^z�#Ǟ�Rۦ�~�Sa�k+���0}�3����ܗ�O��v�%�of�Q�0�~�벬[s
���]z�Ԇ���$�$�Q�����x�.Zg�Ųc��v�mys�I�

��f�Sn�y~M=P��!�=�����Ƚ�S�ݑǵ��f�?����c�Gy}i�����}n�<n�%��O�(NCs��߭D�Q�2H��=��(��qD���ִ��%޶r v��i��q������~[�@�fnj�W�b��IFM|hx뎭���D�*蘐#�H�]#�H8��[�D\��l�J��DZA� �q�Wu��`����.�8��牂�M�w>EV,��1	#6e�_�s��d���+���ߢ9�c՝H����`I�{�,�Þ�i�<� :�B��;*�:��ۃK8lB�B�7K��1.)���4e��Cb�h�Nn�1"3�;'�L�)��t�u<�b9*OvM�]|UAiE"el>zf��΃>Ά�G��M�w�뒾(f�X�=���}  ̜�j���Z��t�L�3���4K�<�_��e�[��o��|��9��ʸ�F�ox��KK��Ey����h�Ae9�u7��|@��猙��5Ɛ4��{ ����c�i�5DQ�w�e�e�mP����T���Og���z| 83^7�>ӗ�wǋ�����0��	�*q�Qn��j�Vڞ���̀Ѯ5{���_}���	��[K�e�Y�b���׍Mh�Sm��yb��7T������"bޔ�0Z31Ocb��9�]�(�-�J�ޛ�oM��W��*f4�=)3U\Z���qn�JՑN1E��<�WV�H����B��C����V��q�2$�J�4�n�-d$;�lj�ƈ�'$�>�Zy��ɒ��-��p�g�����Fd�� o5���L%U�N5K�I/`SN�//Wy!���$}}?`II'�������s�6ǈ�[�i������~O���� *�e��X�Q�[76�$����e�^���h\J��$�V�Ѝ-ay/�f+	u��*�& ��¸�͆�%�Ъ�fz��e̙?縼w������G0���wmo�gԒ�x�6
59�t���f���;Q�����Bp��0�\�K��3&����D0pbel�dF] �^5����{eά���1�곃��kf]�ån�-��,$V����LD� ����*L�m�ԇi�҈*��I;����a��B��7�"��N/�7�Ty	h���}��16���9�!��>ʋ��o��'�zn<���h�R��c�*�Q�B��̢��'^�s�tY�!U���\ؘ��DOR(�n���9>�֊x}�^�W�W�0�rjԧ�o,����}B��>�`�f"P�7�k�P�*��l�Sv��܄�GI��e�U��g<b=��J�����(�J�pf <�Ye��A��G�V�x�-f����9�,0�,�Yb(GыW+Xخ2�{�+�6�X+w�}�E.��S>��J��ڲ���^g�s߶�TV���R����>�BԹ���2o��fR�B6��\ʁ���qM:Si|�������ᩆ��d�;���H�E���M�_���R}i�.�tjx�6�n5��E3��Q�=#��F%�F��T�1��������l���A���{z];��k�J����%��ҹ���p9��w��Q%�f� Sʔ�xhr�#��}.8II�D���<�|mĵ�#K����RX#*��Y�8&�Ů;�(�����.a�J�V��c�I�"u@t}e����3����B�B����/1֌�?I�}� �E�R�������[L]�8��e��R���L�I�
�M�b�`�7�p7{9��H��A}�ٟ#A7�y��55tE_���%G���M�|������8�b���O�� 
�g`��Ii�yp��iÝ��q�4"��A�?u��f�!% ��q�&Y�7���������<T�%3ƺe�p���"šΘ�pق�׫F���W��]��yc&�^1�E-�u���gJ��9��JW��̸p�
n�K�ZzAb�d�'���2��+h��De�t���l���qw1S�J�¶�nH�qŇ�#�f�F�XY���Ly�������j��N�o���XPy��FN�G��ƈ��,J��4so&K��|+�R��5��7g���\Qm�%�,]Oc��@�C�$�݆������i©�8f������y�����n���Е�}@2'i�n����9FȚ��\ �*ݓʱyy���{��ٕ<���X'����V�i=��o�|>َ��h�=vV�N� Ps=V|J������.}��yn��f��.�v�3��jJ���Aro����ļ����v.�pĴ��[�\ y�;y���֔�@�c.鈠ݺ��IS�[>���.��^3��k#�w>f���h�䈲�?v`�ᜥir?��wBs`��*L��"��ùk*؍H�́m^>]=M4�?ݦ�'���C�������0==ۣ%�/�o׷�u� ���b�K,��ųN&7���ea`�׋Ěr�m���X�fq8�NOO�T%��[��W.`V�=r/�v��:
g����I� �s���w���|w.�	������܂�#������j��uH��{������H�ۧߦ�����4�O�ե�����ǀ�Q@3F�>�VL�^"c�;�D&b�(1L
)��帗���}��`���U�}ԉtC�C^]p(8^�mZG~:�����{�1�y�n��F9w�Qy;=eB�M*�8+��%g}x�6�N�8�i9*qBRC�)h��W)��K8��(��5��s����cFǩ[�d�I�Hz���i��ߏ�+ل�]+W�e�3�ڀ0��2*��~���U�	��?Ay%L6�Sib"�c����� ZR�qhhxTZ � �mǊZ+�H.cU�h�$��}�)��48'BgU���)ʢ��y�V|�z�>��>��|sqNr��l�ײ�њJ�;��$��(=%��'�H��;�v�M��6hp�o���N���RU���#�G7k:Ն��S{'gAAd�V:@�X1n��Q��zI��ra�E�e_dJ�(zA�������asN|.{�ii�@X���;���A�KO�jS�.���������ɢ��A_9_��Fr��N���T4�s�U��j!oX5c�U���ʻ�ճ�%����>���d���(��*��:}�&�z��}u�1�>Sr�K���>�0:w|��N�Z֪s�9S�B�12�%�n��j�Iѱ�+��y�tMWa�D]�x�Ln�C�5t�I<�J:;Ԁ4��ޅa�g>�)o�LI��c��oXn|��oP|q:yy=�7�o�@��=�����w�@@;����sz*+Y'���9�[�����L�ym>���=Lr�+�����Sb>�2�8�s���N��z���[�?d�b�\�D+���j���;x	��E;Mx��VJ�~�x�n��v��V�CX�������ca��L�ސv�Y{��e>(�J�|n�o<����[\F�����-[�2�B-PW~@~ȟ��<��]D �KI,�ظ���p��O������a��O)��o�m��M'���� uM���އ�Iz�ߵ���Lڵ����(�X�5Q�*
(ɝ�em z�7Y,��>��Dw�2�<����nIR��u����:2��/  �<�l�E�Ѧ��~y>8Գ�ZR�,�6��ƂA�g��}uSϠ�W��H�Oe����"O��r$1�J�,�1�/��&!�th-
M\��%%�F�º	V���O��Ң��6ҟ:���E��+�.�ë�N�d�vA��G���6�?hp��/�FI*w�3H���	�mީ
�Hs@�oSғ�w��b�s����؏�+&��+�Ӭq�]MQ�6}� P9-�J��/�;!��n/��i��	q�JTE�܋�E_Inxg��c��]�0� ���	D ��&�x���ILJ���N��P,c��7x���K��R�4*Ӌ�ޢru�_9�ׁ/0����w��lQ�'�# �I	��]W��1�Vo�S����:㟜�#yx�"�e����XQ� t�Y9��c4�x餘�F=��/ΫG�Y�бǲt������\��C�s=�r��g��~�by�^*�H1�LB��D�Y�!0ν8&a�?�>�x�.c���Z��¥�Aɂ CK�V��+)UZG�v� �ɔ�l��O��sî{sb+��Jl���?a�L�m�
3�Zo��
*~?������6?�`��,��?��]�[x$���.�{�j�����!���`}��2������^�GofXy.'%'p�>M̈�j�3�/]j�$����Ǝ�֎�%��b�8�6�;��J��1���F�l@�& B<r�و$��t5GyEÇj��:p旽_un�	����\�z[/E:5S�+�n9]ƪ*ϥ�axæX#�ٔޡ6q��T�lR��!n�ťZPjl�N�F9IDs��.���P�(Vث�aJ�⏁c�<��N�3ﹹ����7nW�7�-"`td��<��u�$������]
�;j�FW��Q?(/�y5c��x���O����-�T�z`k�p�ROEr`�%Ot�yV��ob�N�%�+>�(mc��AV�D�jM�@(�n�GV��h�:�x���k۽��K��?�U�&��5�^}�8��4��ɧ|��KF�>眺� i*��8�Vp��d$Y V3�9l���êjLޞ68S k����nj�n�%�K\|i_��/^���x'vv�x|.�IU����Bc�����r�+�I��X�Dr�\͵�=ks�}�@?���:�0����<G�����y�cn3t-� N����|P��|�ﻓ�����h}�F��]�.hF}��	��j��齜z�N���-�a�����֝l4>�W~#V7nY�Pٗ�x[��BCgq�5��[���
{@M�%�u������%ř� �"Eg9�Ȥ�
��3�C���jL�������@�*+���`l5g�U��� V��>'���`d�ekP4�3�z�g�=8��K�����9��*�="=�u2v݄*1�0�����!�������G�̓+�cקS�`������W�Q%�в�rDq��&�N~�E��M��il�����0���Z-WM�c'��g�L#a�Ч�{f�� ����b+������bi=�Ձe�!�M�|6׵��p3��S�q�Em8��ݎ��K�"�S�M]�Ep���C�NyB ��IkӦ�����5�m"4V�6q�����J�/�]�g��H�P��D�ɡ�Zw�z-�YA�>
��f'j!Q(u�	�3�����zB��l��]��l�n���ܘD�[����lL0SQ���6���I ��B�M|��m��8��	�-8 �x�;���a�zU�#�|�ym	8z@��$��?�z|���8�Kc��녗�Ժ��^�~V�¤uA;�f�㛸�醌��WG5��F~�j�Nʫ���۴x���S����*q�;2?�9������ ]A�i�I�Fݥ�Pn3���0�=��[O�ۙ}�%V��V`B2n�v�8~���Q6�uDž�cq��L�d�A<� Qs��X	C���ĉ^$~E�<$>�2���Vૈ�)�qm�%�q�P�u���۱;7����VIm<��~n8ҥ����j�2�ǋ"-���R����h���C��?o뤏��#�����I�)�u��ݼ*�$/Fn�l����K��?�.@1=3��%�ߝiw���0?v=�Z�a�S��S�R��M+�s1��	�gi���x�pX#x%��M��j�u7?.��b���|S��Uq�L$��-N��Ը����#�	C��)Or+�k��(w��`�
X��=���;�o��=7�9ŏ?+����;�GY�}/�f�y'z��cy[Cl-ݞc�s�dn3�r�Sd@��5�c%��y���!D��FpfY�f������N�k��
�S���%ի=S���3�����2�W�����	,����d�1�8_�P|h4'���r�b�%����4����`��Yw�Ę�@	�TR����O�y��=	��k�"h'���Y�bGI�}��v
�	Ȉ�knvkZ����M���TG�G��3_�<)6��=�hd�gzC6���r���G�K|�mM� ���o�����3t�r�|by�;��-�(bb�O��k.�w��s�����5����Ӥ�#��5�5r�������Rk�䔔�!�AG�*yų��ġѶ�|J8 <�Vi�VYhrK���N���pI�Z�)�@v�sV=�[����M��s�ޕ�������8�k	I��k���p�x])�6��8�$��qwmB�2D�dC�u��F`�<EVuZK^.b���	�;���VWf�P�����-Ԡ�%-�~~� F ����!�bF�2����#|����ݠ����]�/$���L�&���\_ڡ���C!*C	|DR�u�15�F���6�I��d2m	H���m{ ~��~�ևbR%o7{��>)1��v�� �Br{�E��&��EK係�S�ddu� $0�\acW�A� ��e	�l��<��F��6;�QupJA���7��LÉ�FŜ��z�*�p-x/�)��ӒCWx�Ư���v�8G|��̜�?���� >e�t{p|Ug�Gz=�>�����@zh�2}mD����$S�l��x��g5�����j�P而��>ؙ�`1Mm �~�����FL	^��5e�����{���;0�Y
9����Ͼ��~Pu+���_�(��uر{H�v<�{�u�Ѣ�S����|�P`4)���1��>�=���=�|F÷ a���~���qy�����;a1*�u���t���M;��$��BMI�j��mlN�K�hF�[I ��λ%��(������A�A�hu��Ū���JlE],L=̽&<�M�4��#C�J��'�8��j�rF#���<vF��t���?�=��2�&�xR��C��xD��
�A�E:�;���"�C�Ua1���B���H������\�#Uq�#Sp� �I ��W��;L��r_ b���k����5:�0D>W�YH:�شGP��j~�]�t�w�#�@;�`�Vlǵ<Ԝ��Z����Dl�p_���HRǪ��)��=��o��u'9���ߞՉ�}�|B/ �tʑ|!Л�ׂ�H���cvW���vٶ��S��$�� ���ëb	�������)Xa�O�4A��ac���Q��x���.*��Y�����`V��a^�N`���Ȗ�{����QD#B��m7P.np�0���[�Iq�6�Yz̛�d�M��'�~ST	5��F6�/�z�(0���vgs��g	�ִ��eD ���:~N�o�`�t���#�xv��:7��O��跖�Rz�+�Q�F ����%SHN���'��I�~����T��~>M(��x����jV��|�I����,�1�郁鿶�_f4t�K��Ǯ�/��7��)XL�;5��Sx���l�/ΐ�x���m�=�qM���NPa٨4��s����r��
�p��#Z�2��;|�9E������i�^�~�:+��?J�~�����$`\´���]E\��oB
����dX�����ч���F8�;���r̆�Kw��NS�x<'�|~]�"��� F�h����:�r�+��~�ˡ��l5���r;�Q�٠������r.N�ǐ�3@�X`�5�=���Þ��qX�0�6�:y?i��yb9��>i�&CU73XǺ9�ɴ"
�{�̊�S�v�`���ebs�bM�(��%S���=�m��yI.4��^׆^�2$����!{'��Br�o���^�����$ɸ�	Ld3O����ߝa�yG��H�3sX���u������P8�B�f״��x�c����F���3��}p��O���Y%dQe;���b����'�̙��S�l[���i8����|�Z��4���� �C:	�W�� ����f%'����v^X})d���e���������_��$����-�Mޙ4�nB��B����.(%e��gl�4nC����>}���k	S���&��?V��%��e�r�#��FJm��s���]���>�Yc�b�O|!�C�$�#�~���V�	o�pUG;��PX�RmC�pFUI���|?v͜����uY�]C���c5p��ڴ�7ϵ�	v�t�F��3Y-���Ch�2N d�������SӖ��@Gr�rd)�>@j��V���_\�z'��!� W�1�Ud����*��M
)E�J��8��~�@�1<��q=�A��1�h�(��eI��Bt�E�Ȃʶ�n��$~u�@J��@x���ⵥ#C��Sdt)�
�L"/;Y�1��oX���J]��x�k-H���������J#�]g��:ؒc`x(���ڐa�E�v?.$?������ G������y���[$�0��dp����|s,0�<)�^��cۂE��`8���z��'r�`s��F5�S�N�x
״�CL��"����Aم� ����=��+/ʼ�������Jga���,�$��GYF�����|TD�C� �-�B�ϗ'�;�$�G���194+a�i2Ǘl��:_v�1���>`.��#O�&�fL��(�\���c��a)W��ٷ}yh����nP��Ml�^�eWx��w!?��1^;�Rn���jW���3}��C�ic�H��E��e���ep�}�z���ʚ�"S<}j|F^�����z�!�M���[��.%@C�;���;&��ǎ,%�ۤ�x�ٳ;� ���Fl�O�4��l�u�Z�5���H���p�8�T0ȡ-�N��aM���lk"OU��c6�`�{�`
"w\Bu����x#}����0��)��?�����R/�?Ih�y�i��Ne��}y$��[!�{2a:�)Ɓ�rN������zm�
i�-�Tu2$�n�5��+�� �����x�W!<�� :[<y�
�A2�E��s2�-H�-�g\x.�%A�=ʝ��K��� eNe����W%�Bs�.�h7��p� x�~-nV:�H.�h��Z���ǒ=e6*>��#��HY&4��MSׅ�!�Ffn�Ws5��e��|2��Z@�s���g�mjh���}��%�b�Zt�M�k�7��BA���7N��6s�>��KL�k"_Z=����l�dch�po��q�\p�diq���Qw+���6]�pM�͔�D�
�?�OWٻ���t6��v�hF 7y��pQ���t߻䇀���6iO=�X�`�r��"?��mx��n:ę����l$ �K|?�4��6 >FͲ���$7���I�jF��� �Q�z�>��J�ICpt��lI̱;��r]���ml����@Q�)�5�FQ�"K�[�=)��{��.����=볗P�Yn7<k��}�C��,���Y�#B'�B�Xo�$�=�[����To��!�,Vq_�/��ϒ�M��ub �̽��il�4���Ve�킣dA~mūژQְ�!�eX��>�/fIG���E�3xl�g�'=���>Bҿɞ8yT߾
�?�&����2.E=O��10�OH͍R2�KoT%q�$���e��C�� ���p���趏��>�b��f�7Xڕ�5q�{ y�p�V����c��j |/r���X&`��~q#<��'v;�Z�n����w2H��7"�$ۤ����y��/"%'5r8���YA��H�7���n^6�_��l<R��J��t��t��y�K�^��ΩiX@4�z�$e��+Z�+g�I�w��ݚNJ�,�"r��f��ǿfb#�t��t�ƀ�Y�Kt�.g6j�ڵ�$KxdU�
��[K�G��/��W�I�o�&+���5�=���FU��,�^� u��~�R���a��I5���"K�/�&���a.2(wA�Z�ٜ#�=7��Mk* �[b0�I�]<�䟫V(��Q�^U���A����3�=Č�U�JS팝��K���FM �&��7ve��[|��0�%���Y#�I�69L2����q���ϊm��G�d�7B�}�\��ŕ���T�N�k/�xkeV���H��Q���`�Bc�ŖD��8x�Wl��b�6.z���($4G�r���K�ǚ\��KK%aYυ�(5��X}z$@�;���UP��%�uY.8��0���5���*�h49T���PЧ[�E6cV�hd��ڵ�[6��#�HBR��`���Ø���<T�N9`*�N���\rU�	^�Q�Dx^���1a�������=�i�R���T�U3m�#�<J�����v�f�/_�_�J'S���b��R��.�&��:�8��#@ ':��C+NV{�W���=lw�v�!�X �oIX���\`���O�U<��Kh�[¦st��7��'�����U���d�pg��mQ`CDp -�ˡ2Gaz�T�R{�r��/��KRPuܩ�)8�K�?[�A�	[�ߘyg\C`6�Y����|�����1��E6)�hf�/�d�f�3�?��r��]DJ����']՗%���.[s�b8���l���W_��6�-Ac�q���a�jhL��������\0��n���pT�F<�~�5Sd���\9�7W�¿ax��4ÑC2$�)��5����2zuξ��!`ᘍ$�rD�^Gc��B}�����x�kI�%s�F�l���K�'H*�e���/��]~�ă�o\þӮ�;G�`�y��;P�Ѣ�L���+���ȃ�+��-��OF�=�Ō��[.�o�ǽ�����H�`v�s&�9`-y�w�sۀ���51m���������PG�+4!�����j�7FU��X�Y؎єm�Aq���	ToF,�r�L

Lc4���ē���LA��I%eh�6	�F4�v�&���ٯj��;l#���knrO���wO�;cz��e�-u��>'���Oh��#n"T�� �)'@�ڦ�� �k�l��W��~Y��=ez����,��W"�?��sa�>��0#�%�t���s/�Rab���b��p#�A_NUs�+�9U�dE;lNA��p���۳�D�Z�/|�M���BZ�`g�䙙]Uɐ��w������@ ^<P���p0���?�����
����WCkZj�)�Ŝ<,�������Q?N���D��(�~�|�4���[P�RH���
Ѫ�s�1�͒�m��w+��$H��/��m�~t��@���|a0�����`8�-`�$����8=6ͼ��S�GH����@0�^��p��RE, /T��g%�� ��:�4u�m<�M� M�y`����$v���ε�������^X苌�E��LR+��l��ox��HT7c3�9�Px1��Gp��d�TA���wq���H.l(��J=f{p"����:�Z�b4;Ƹ�.�X��R�W�,�)�"6��^ %on4R?��!_��`I[lH� ��!�?�ρ0�E|N�����KDD��mϭ$O/S����!�^��x�X�s�#b[����k<S<�k 8C�o�u�)��n`��I@u���n�4C��9�H�����ϫ�s8���@]�-$�2�PR�S�G�ʆ�m��V_�ME�"(WY9�Q�.5�@���#����md#�P�hQ�ig:�~,v�;7���jk��$�-j�86i����{@�#$7���MQ`w�<�IR��+��,m��nNg�J6�\p�;���z��jF�^��{Y�0� g�3���7@E��s��^��Ν\�>'��n�g^�H]��dڅ����3.�eWI��5�[I�=�Uк���_�T.�wz�����P����*U:�,����cn��j2������(eH���C�Y�Wmk�o"���G�ȃ��z_NaU�w��.b��N��8��"�W��Dky�|�{�V/��fQ�-̼�|.�Ġ�R���cI#T&������������5M掠=��7�$���ܑ��7e�<��Ā��F3��%2̤������Ԍ�@0i���	z-��ފ;^^����Bհ��E^.آ�@�b	@�׮���������I���]��@���E>��G��g���|��1�N<��;���^p�l���'����~`�nZѿbz)��4�~R����Ԃ�U�9�����O�D��j�����:�RM"�}r�dӑ�ӷR�ɠM���O bPvI�ʨ�Cqȱ�gu`�DzA:\��^��]�χM�_��Z3����eKO!\�3�f2������'��~�6],0'�h\�ӷ����i[�_�eh�������)�%�V{��϶�1L�Kơ E�>K!G�V]4�Q�(~�M�����)r`�\�w�꬇XA����9<�0�� p��	6�T�c�Ps3U�o?^A)��A퉸�I^A(�Ųp'Lq��w
�ƞ_zXl-�+pvJs�r��3�Q�n.��ơN�	e�(�ea�7�9}t����>�}x��8Ļ?=������<�Fcn���8�3!�6�"�C����L�b:�a_-�� ���Nv�P;���p��=ڭ�(sz���$����A���t+�Z�qVb�7��N	��=�1���oG�4�_�^1�����Iel��		(gS.$LU��z�y�s�q!�M{_	���b��5��j^@�:�~�i��1���u���u����2�`��d��n��P8e/Y뭦�׊9������Z��Sz@B�kZ46�'
BF
I�n!��/�f��̢M+M�3�G��߲>L�g/w#�� ��ԇ���ڄ�	��ǒ��<�c�����񶉢6o�S�e�<� ����eJz��!��.�ܿ�!B����ՙ�uC}����Bc��xM��l�aX�& ���=��S���EK�'g�MX�e�yn��}O��+��% ��5K�Q�d�꒙�l���<W�3u��Q����2i�jo��G���M�/~E`�]R{�>ۈw��%��!t�	�A߰��R���?��vh����!.���-U�]�H�d��5��B�m9���&�ݟ���.�
ܶ"�&����Wn�٪�w�����(R.��3�b腴PD}BB�I]�"7�C{�����0�PK�����A�X�>�f�F=�&��I�Tjã,#$J������-F!��Fb$1k�ōtț�ر�k�+Cv~'�t��Z9��t�yB#}�� /�L��Myg�B�ʁ.�Ò�V�����si��-����l<����J�7O�i�Q#o�7'��"3r&����^��o���ޮ(*�`4��$K�7���=в'/�C:Q��זd�T�Č��:N1��	��&=��?s,�"�����4ǉ��w{p���4ȩuiBw�W%���O���P8O-W�I������0֢�/��	g��Z����D2�yl�s�s�@ G���6�
�*�-��u�a���n��[�LD�zj����N>�Y�̥e?�`��[������_�o Cv�[`qt�ё5 ��㒡�Y�i�\D?%K\��ƶK�_�GʩN]>���)��_��D>'�e�`rK�I��xR�-�=m�^�pق�Ʒa~�FV%�f����U)�N�Mm"���inj8�G,�QK#�O�<�., �kv�u5�@��,�٥Қf�=�����/����G5�Y�����/'m���	����78Dn���۸�]����mƍ�^�Z��h�v���=~c'�ŕ�/���A��M�ԟ7�Q}'���O��P������)�/��EhV������SWac7��X��d��NM �o���a��j@O�I���	�k�<��hv�8�]�`!L�(bv��h�
L��GK_1�X����YAJ��3z�����0E���c/9i�L����A���HnvbOLq���ܐn'�1Q\I��g�T�Hv��։�wr��iI�17l�m����~��!I�V-U�L�k]~/>�xtG�S�#��e�_|��kѣ'��Y���Dq�pzz�-�ia���j���n���1c�1_��)]��	�#���� �<��$���;F���.?�ogy�sd�I-�x���V`�p��h13���R�R�҇���`y�����ݕ�����r���Oa\��P׵�p4��i���S��&��X�� ���x)[�� �-��Bl�QZ��O�W�7��� <9V�%���o��1	�;��'߫��R�E�q�7�?�w��&�nz���p�������Ӕ֛hS֭u���b�+1�q�P��K���9��X�V��p/���~V"&
4y���*?w�A,�s*QS�������(x��ʧ�Ʀ���}�/�Nve0
���V�����u�m�[�xw��?[���Ӿ�֢���!��S�,w3UĐ�2�ق80�PY	*�`�v�����6�u���R�+�����J�d|���u������ĬB�E�oS��\�6v4нŰ�|X�t]"U5�(T.�﷓3��0��HE#�g5�	K�O�<��W��с��Y[Ԡ��I7-d���	�7���u]�yy�6Q�5G����Y�.Ϡ�5eT|��h+RI�����t�9�[��[^��߳�bM��WuF���a���O����s-��K�=�o��í�9��Y�Ł� o^�NZ�%��pNrƚ���I�T��Q��q�2��T���#�u�r�{8�4b"�o�E������~4��6�2넜s��ť'���0�yU�f��أ�*"?�)d5}ԏ����V��׬�ą� a9%k��2[�G�b�(Ԛð��\��Hc�6�4CyZՉ�O�@�g�g�#������x�5c�ݿ��ܜ�Q�I�݁#�3@������N`P���a��m����y4ta��I��5�<۲堄��b���
��XYI)�4�֤�R"
zދ45w9<(�UG_�;p�|���^��e3X��8�ANĩ5{�iF[�N�ܬ?�`�np����ܛ����,�i:q�^L�亂�,JۻPI�ե�_5����;z*���?<��PE{Y[ZZ���>Ҋ����T%y����lA��tT������t`b�@��48���מ�ɳ�c&�N4j�t+Do\���8�ΔBuX��m����=Ո2 �����p)�ϟeH|z=����?����כ��6��t´�oh���[���]�վ㤏��O��6o&�?e�$mu=Z��t>Sg�U��)?�<j��hH6�Xso���v�_�(N��e�^jޖ,�DV�h�@u��ZҮ�m"-a1����.����|V��, ��9�i��"�OCYdJ���<1����,�(;/�8۫��~	���.~�T�|b�=;'4�<�ߡY��￳�W� (�Z�?ܾ�d��6�� �/���m���j���R[�I�m���A�������t���s�I�r��9ӥu�6������U�NM%�Y8o����D��i:�LС(��yy~��$�̋4�PR����Z����E���` 7���Na���pL_T�@NVx���3�hz��úЇ���I����[�jΊ9��8S��-Z�-#��z�3�އ���Bq�Z��3������S�Po{��LJY
[���^�9���fG�C*�z��v�G:�������d����LG�	�Ս�,��fK��SϮ�t����u�yBF�c7/���Y7�T����a���:gh��FŬk^�.����t��!Z-:�{�^���/�([#=,�-8���x5|YlMt�wdz��A2,�T5�ω$L�rq���`%��r��k��}���&8Zr�@�a׃��$�Ւ��3�o�(ݚC{ت��Ɉ���uQ�����"[��R �#�k�gDp����SA��X���v�e�U�-5�R����x��Y��4�q#7C[���L:N�u�V?Gm�D����c�#����H�W^�T�Q�bfa���eT�N��tZ�P��4v8��fO��3}�~�ٰ\	)���F_���v1����͂ҟ݊m`�zYL�G5$YNh$���w����K��ƣ�}Z!��~����?�i����Ѕ��I��/*�k<4`��s	:f�?�6w(���^�Y] ��x�Dq�DI:���;�́I��7+U��oH����R�B�޾����OGJ�J<�m��7~DO˂��E��V�fCo4��(�Jʟ�-/0S��G�
Q�40�=�R�k����Vsp{ ޖD�Qh�Zwӷ�� �t�P�1Z����vX>m#>� �FGYv�Hn�'�$�����yX
O���^dy^ \��Y�����?�N'��
 ;u��$0� �3)I�`�h	T�a��9~�˪dk���`yMyq����%%�`O�s��eZśD�܏i���!�ɳ����X�A�} ��i�zʸ:ߖ��s�����B��&f�o�b�V�<-;b��}{��R�n��)�aS�z-=�n`P�T����;�B�����9Ot����8O�=}q�ר
6q��>�x鍼a����PF��e�b�bI>�NG����u���{�%�֝<��lM���ʄv7�L��1�<�0tU��,�1Rf�Iqͭ`xډz��o:�З���9����?�i��p2�M�l����	���܀$�u^;�7+��S�<�¹r�����٧.�v�f������	�px�;��NDk��`��'n��?ESe��ncf-yN�qbG����U:-�V���B�|n�=O�/  �M��dܨ/�t��B�����ۆB�?��)��VȶC#�;�i���o�-��"�&��fR�/f�p{�]�f��?T�oNF� �L-Єt6��)BD��
�Ab!�|��E ��[Tr�ot\�Mԋ��(�c��[�v=�*Y����[�̀�"'�o���.@5'!�9�)|��}�1"o��w`�z�a�vت��@A��M�i���:���"W$��A�H���`�U��-F	{D0K�T�cZ���T��!�.�Z�>�To����n
x�{۹a��<F��]$�L&%��
�/�Fi�Or�ւe�=��"��后�,��KF�:��~T9u��:N�Jn�%e�S��~P��^����}	O���6����G��9�����ࢬg��%Zj_M;����+�Rh���������Y��ISz#y���s|�HŶR���@����TFGi&P���nNAv��7�c�S2 �����'�c�����q��#$�niW��>����([�K)%���C�&��:e3�2}�E�2�uN�^yR-@Zh�\�u�������_`൪�A)Et�T�hk��K/H8N�W&���K��*UE@`�H����>�P��{`��[f���EDa#>��<��+3�H����*�s���ZWs�S��9$>�>��#~�v�T�+��D�w�V5�%��f�H!@�#�]�MB)Z�Ȅ-�i��\*��z�(d-:c��/��{$���wK
ޖU5I����A���C���-Lg��]X�ؾz��
�}	^<0�O��ވ3�V,)��ؙ�`(�Ƌ���w����+gq
��W�j�������\����t����'�g����!�"|��@��8�j@?�I���������E��\�M�J���p>#�����)����tK�|#b����n�����\��UY."fM���\�j4�	�'.�Z����;s��.�, �@��i�I<�[9�#� �u�)�׽��iR��߶'6���1��/�J_��oA�o2��y(+���J@��X�����*������X��8W�f�8��cF�V�����H8kL~�[�$3�u�t���G��T���)�_� �[ɮ]�}��w4��WiI{��$g��k�����B%/,�;�2/�$&	�e�A�B�P��K���q�Z��P�繹9� Ԩ�
���9k���KĐ�CS�����p!�
7����u�M��*7cZ��Uh��9J~Na��-�W�H����8��bU|(�_�(�m��3"���]�%v�Yqp��R�q������MeR&VW/����iD�d�ս�+������T�\���b�1�Ȗ���R�Q��y]������^�M��98�$���R���[N��\udW�Кt�����.2̚78��Y}ܩhZ=/�[I}B�+�V�jۛ_�t1\y�+���Iu��_��[Y����5M�Z���G�(��t���ɜ���� 
����1
����������vصT�������5�r�� ��/��W��(<8[P�#䫚���~柮r�����h��?���8nۧge�vڸ�l���)�f�/V�l�k�"m�-媎6� M/\��:$!E�so.�c�+�̼I�ǽ��#hQN�v1kx\P���T~��.<���������F�Bpv>wl��G>�9�D��*����	y��E�+�?=�s�
/|ʎ�L
n�r}��6<�zO|���	�� E� � q0Aok].zI�%r��L?�p��u#L���t����$t�!����?�Y���{{ 0Y���8/��!�C�$��Ǖ���թ�C��0�'�J�������cJ@�-# 7�1G�n�6�_��`�/�>�Z<�c�Wv`����)��ȍp@�*���č�Uҧ>����ߤ�*y?�A�4^5o&N����z�����G��aEX�E��=6[����0C�8fT��䓊=]1T��(�8[���î�*�� �@Ǚ��!+���Y��X���4�+�޻F�k?;�Cqn���Ĺ^�]�Xjb5Y���d�Lw��e?���'{��������#�x+L�{-�m�,��ԩxR"��2�L����H�<�y�13�o�M��E���P����6�ч�T�.B���9��\����{"Ĩ�$��S�#�
�U����͔��:n���P���^3��4��3Y��p������r�̧7�͡ylº�|�/q���]�2�bG���&�Y�.��z%��~E�
�6a3����y;�x��k?M�0�F�x�Z�E�:���Z�z����{�@I����
C�d�b2�OS\�.�y���%0��[�u�V4�stj��mM��k�KX���|��.pzq�#7��עn���*���K�%�F(h1C�r@)�
H�k�-��}<�Z���T{�4!��a*q{/���"&;J/��
��k��`[�L]l����g\S�3�A�b:�b�/�׶}w
�0��^ds��Ї���4T�I �/�s|�x�n����߀���k�I����ԭ�2������!�Py�|�v�N##�n�1ז�k �&N,����(�Ԙa��
�ZT�����zf����Β���vl�شd�MaJ>�+F��ƅ����	7��
�	}�sY�]�� 0��b�Nv@*����~��F�w��O�$'P���ݹ.<$1�Cpz��@�	߁D�4 �B��]��P��&�����Ⱦ�m@Y�y�ޒ�0Yav��%����j=�89���,X��*�UC2��,a��r��wM(�q�皦��	ej���{j�%�0�+�h�Q��L��{�M��O��6�����z��kh&�s7��8g(���Y&���,!��6��U��8���R~���<4�k���D0!�����v��bĘ���M~|��矛��C���!r���ۗW�"&<���ѕ����+ ޻߯wz��_�H�A䶭K�<�C���L4Nǻ܏䄟��*�a� u�_
�ǶÑ�$�6��|��!�Д�߉͉Ӆ��E�]! 쯾��w��u��}\��a�R�@2����2�M�����o�;��r�H��q,&���=�π�m���9Za/��|Õ<"�� e!�Qz<��$qOۼ�W�B�9h3R�iC�jL_��+sj6]���8��A/��� ��0 �K�Z�2+ZX��m�;�8��%�rޘKXw��7�N�	^:�da��ta4B&A��%ə��	0��=}'{�û{n��[ә��>�- jq�پ6�i�,>G��(�/@:X���1~cq.�P;������]�}\���+*=�8��G�W�Č�����!oAc86��Ɖی���s 
@���뽦m���`p�\������%r��FI���D�Z�-6��q�u�qD��
mID#-e���]e�l��u�N����Ȅ<� ���'�f��c��Q�i������*�B GZ��M�򙯤���4��B��d� ��6�o��גr3��T�J���/�8�v0P�V���V��Du�\d�ߗΩ)[vV��Z�u�`�ʡg�:4P�c��C��Z��S ��$���3,�C��:���uঋ��/6Ӱ�a8�zZ=ڙ�Ĉ�97�f|�dk,KR��4�]>,d�A�ID.��f�,1�)���j_�;/&�5#v��FM��z*J=�<Eع7h������qt�01،j6�ε"M�x�P��^x�Z���yWiZ�����]�6�� ��ȪF��h���ڎ��-��aM�Z�߯1��:	�|�������"������������bs�(�ih~(Tvs/47�s��|�` Z#.�� ��~�Q��q�%�J�@��ųj�����0��W?r��a6���^���3�r+�/��ft����Djƹǰ�_����`�򉼵�a'8�Μ'�� ��\�Ę�N<�pV"�!�*WxL�����P�)�����9�-��ˊmफ़^�hj�܄g�D)�NK�"�n�dr��gZ�Uoڰ�"|W��/��_wjA}��^�r��Q�W����?8
.@�!;ۣ�S�'k1�ݖ�{�k�>�����!w�3V�2F�8s}�:����G~�7��:Y4�~��`;}́k���i8�2v��x���&k�=��y�:-`갾9��ԇ�"��I�f��Z�f��"�jа�^FL-�0- 9~�*�/�5j*>őEA'c��~�]͌G��?S�@�zA������C�B��B�n�[+	ed%=�s}�#�T/�l�U�Hk���U��s�Y�pN`�%oEyje��)��)zG'��΃�*p0��^�*���X1�я ��^�L����6�ȗ~�Z��l �ȩ�a�-�M��1���%?��W��!�� Kէ�8FI�N
c�����pe϶@$=��� z5A�=�ee�7H�xC]��	m��#�<��u�3}cT���c��rTuT[0۟ȹ�#B��-�G�`u�Ĵ������Q�ӏz�����mm����3��P���UV��^w�*��0���=��;4!ȧ�kB��{���k�./�("�;p�߲ԣ;���5������$(��6�*����GH"�f����,�	��`�`�0k4�tYOs�ɓ�<e������O����e����2�W�(���+��d[I�З���PU+YJW	�y��������Kq��]>�A��C�%L0.p�t{�|9�@�*����ًg2��� n�Ho���� �Ť�"8�6j�H)D����/8|�(o�kSe�aG��fLn���
RI�8�9`y‖�|�:ò�Ҿ���R�A� ��W��X��d�fH�AL�r�P�z��H��Z�ϩ���|QMe�������ft�}&����%�ؖ�~�����C"�-���v�}��9�Uq�'5{������H��sc�\t�њG_��Yy5����E��t>~�(��8t�?X�{L���IJ����r�Q��~LYx}�';�J�i����4{S�u�o�$ĵ4G/Qy�%�)t����L����Vm`��4�k�27C�ƹ������]�-�*���i����#�a�S�{�:ړ"�t��N���������  6\�����
<�,�f��8Z�e!kSC��a�@�������8�<<�g���^����3&'�J"n���(���]��+���%�F���˙���)�a�U��"f)�E瞬	m�)(���3���
՗o���z����P�\<���3��<�����T��l4�9&%�\_s�j���yv�㾲�ڟ�*J��O��gעj3د�[J%HO�rhg7��B)uD�%;��e�!��@9^u<pt�(�y���4$������9AtE�3�5�eȭH��Н% 8[����s�f��,�r]�����@��>9�T=Jf��b��^��h�F��!�0v�c@:s�z�}�A��y�gv��ku�!�+'0|G��nɀH��420��.i�M�Lhp���r�FBP����E��T{|�7�`qa�����vD��a7���5A���i?��8L�Q��̓��$u�eM}e�ׅ��s#HC1<P�_r,��3�%/!�-�NK�Jv��[֝�x,��Zw_ݏ�۫�������@ȸEЧ!�ݚ���`,�+CǾ�b��P>^@>ng
���)HD�X��8��-z�]r$����^�X�5Q���
Ǘ�3��Ou�kM3�-_I0ߢ�6`�kw��m=�)��aU�Wm�������.̱ʻ)3`Lp,a�Te����6a�:� �4sO̭뎰��Hj|?u^�R+&����cp)1ɝ����!Z�"̸?��yQ١����a�jM<^�P+TKh��C��~��e��U]ZCǠ L��DG���QI�C<l�M �v�s(�+�E�O�ڳ��L����_�THo���S�SG���w�Go{5%��������6}�'�^)���{�4s�ó�2|��ܮHT��іs�aު!�ܾ�5QE��p�K���oq�GS�!dc���?���\Mj��2I���iaz�uN��Z�]�����~���%4���3i��8�]B�D�a�������7�w^�x�.*��!��SD*���;�+�C����@_���	%6+��wg�z��;J�(PXPS}d 2"����Y�Wy�@�N��6�R�AUҟ � ��]��`-vy�P�z����"!�*��2�e�\JW{U��2�|��7�t�9w�Oѳ,
��e�/l�Չ��a���VU:/�ߑ^N;N�w�,Pg��%+�_2�3�B4���w��K�O���n׍�}υ�2a'.���>������f�Z�E�!?�����됣�z MIlN��6YV��H�nzh��t�uh;NP�#}����o�L������ \9)���O5%�y��Y8S��r� {t���EҾ�Z�"�i.�8"r'=r��s� ��C�M.F Δ�@��}��\��	�G���+0�,GH�Z�cZ�E��"� �ں�4|�z���\l�㋛���y����ZoHS�Y`��Y�۩h$�Z���PX(/��Z�{�g9���g�q��f��}OY� їt��^�]C�
�dE�Lw�I�՘�<�!L�_���e���V������~Ò���h,�B@��r����B��J�c������s#����S�d���Ʈ����R38�xh���I[;� GR����d�)%yr�����x��u`�wmn�Fy�-�U��D��G����2�(�s︶�fX����X�L�Ǡ�l��л���8�4���~[�����2���s���k����cy֟m���L�d�����%$j�T�|{���Y8��8$��8�����q"����f�tOct�%V-��L;����yO�n���!������L�����U�s��ɀ7:�_+��zͤ� ��w��D�{��uLǼ��g�Q4fi/6�k�:?i/;�]�,���q�u�K1w�����9��yXM	ܨ�����t�|p����$����d(�������IAh�~��k<T`�w_,���V�ZV���W��� @^u-ٞ�
�f�w��NP:�}�%�C�O���cN�H�o̡�[	����It��R=��H"�z�C�<8SΆRN)�I�h�9	�3���S�����=�+Q�q8\U�C)KqkǞ-���L�Z�u�lK��%�F�@�	)���nQ���_��+�TV�p����%��l���s�N�$�{�>7o�j}?RҢ�*)��1 .)o-������%I��}V�	���q;�u�׌�}�|ʐ�+
���b1SS)�&�M�y����ރ�.�	tJh�Ԙ�Zq�;{���L ��F��@��HKݻ�c�03���#�n����9+_W[��W��U�'A�$&�P_�V#��f�ΐG}{��+�F5��E�@���ֱʇ~�Ua*Dq��UB�1LF�M52G�q����@��\b2`�!J�6������gv�E\P'��r��1iP�c�w��֬zIR���U�e��a,VR(7x?%�t~����*���y��<4�xpM=�j#�$�j�|SY=�f�&}���k����!.���	V��G�h)>IS��l��:�6�vԃ+�1.N�64��36~Ex��G=H���zL�j��`�Y
����,�E�������S6��㼛��B�|�ڱ��q��~B2(á3t ���F�5�,K��=8P�1��M�bd��79��̽�]�2�&N���OqU-�4�[O�p)��R/��+i�����i=���}�E�IVx��d`����l��"��+
^�C��@M�g{�vo�竪�%��Rb�u�ss�8��d��7��*�еd�J�q���_�I��\�n#�g�b)�G��A_I�Z0S��D�:�d�nmz�G{D�I�0 ��sd;=��M�臩T�g��Qݻk1��x�P}S,��B���n#Q�p��ƒ�8�ȈA��"&o�Ņ}"��i�!���K܇:i��ߍ<��PQSf�[-��r:j�:m�O�P4uB�h�En����XS�"�'�w�0�&�4
��7^��i�z�?Np���ko<O �Pb���cL8��Rg�y��kb��O�<��֦�CV�Q��%�q�0R�`�m�hZ�1f��5�u�$g��5�CЙ�.��9{l�|�mab���u����Ͳ����1�0�I���Л��< �T|x��>X�B�t��$)椚����5�:S���*!d��/����@jN�Һ�*i�$�k�����_��O��*;X��=�>��F�]fG�~Μk@c�Ma���q���?�@^ēy�G{�n5xfAf�s �7T�#��AQp�)@m��^�ށi����3g8��`�Jt|�(�TQE��}6rQӟӝ�d� B���'�Ĺ\��s�jz�ѝ?�9l�5\�S�I��{�{7��1��{����_Rp�>���#�`�L�</Ȑ ��>�h�h�"�e����2��fYN�骾G�k�f&%?C�ْ��=޲+�}�����O]/�ؗ�e^�,n���^���	�{��T-����P�Lj��Ï.������V��6�/7�f�I��=@w��:Ҭ
^!�}/��G)�� �i��und�g�?+k��A@@"[����~8u���%"q�0�C��ćF�?�"���͚����,X����i6�`� p�?k��u��d	�O�?�����ʯ�<�DBd�G�})��m7�!G=�U
pMB����Z<0��k'm����Y������++� a<��Y�ʅQu������'nY�ia��c��S�7�Xn��H�S���.��^�<��Ύ6�t��b%�o1���-*�_|)���-�� �A��"�&��k0��{�4��yi�u�t�+��
&e,�2�-�!S�v`��;��#�?;��M5N����Y�'�͠汗2sI�+���<�����RGA����)̛�R����l�}~FΞ���AM<�X�0�5���/���;8���Џ9�#!��-�ئ^�
�
{|8B�~<`M���p��i�f(e���,�+��ˌ��\�����d��J�_�;��֘C��v��t�nJ�4�-Q r�����0XJ\k�g2��gL&O
'F��Ip?��C�\��SH����ɪ�<�%͸���7A�I٧\"�Kjs0���d;��%�(�/�p�E3`��c�
�~i�E�g�T�HX�8�+s�i�m��nrC����	>��I�Q�$���DZ.x�|M��b��0ig{#�,8N�y�Vn�V��/��M�ȥv핑0r���������8u=$0��\�Rs%����.#����ʣ`��8n)0��Ϡ$�Y���rM�դݿ���H�88��ۭ������2��d{����ɸ�Y�&w�ڬ�� ^��fz����m��٨�r^����2��Ԫ��#0@��c�O*t�:f�����qOgz.N}m�8�Q��v��<�(����r�}�G:KY�݀ը�;���a��q�������R�
��`kk��a`�iI�gn\0���B[���N|��G�Y�d�*\�*-n�	�2�:$�y0S�?�c�Ѓ�k~�����u�\:D���^'=p���^�xЮ�X2�A�)�>7�M�j���M��eI7��]Rֹ���i/�&����e��d�Ct�k�g�u絧wuD�y r�pmC7U��*���{��`�K�T$���$�5I��aɴ[<ß�QTK�V��]))ɯv�E��0� ���PF\j:5G��D�UWs'�!��{�3*��5�p�g��눓l�@d�E�>}6�9�NZ�|���&xt�F���7ne�@�Ƒ��LƟ1���Gճ��xb��K�$~��.e������ ��(��92I!l�33l�]��y=+�=J&������rR�tY�C�;�!Ft�Kj�.`%f��|�����k�V�v�mF�1[�Ul�����6�����&"X����G���Yt?����:��dh:�Z�,�������Mѹ���أ�:��A�;�)�M���3vT?-�l�0ӹ�I<rz_�5q�%�����ۖD��߭�t"e�a�����|�_c�)�2��5�IxΦ+��Q�h�Q��U���`���J0�$#"˱E�o��dcT(0��(��Mr3�#fQb��AQ��jI���e����|����}�	�ɇwq*���80
`V%��[��k#��F�h)���Z��<C����O�r�a��dӺ����*��"L��ى�K#R�5��av�1 `��;F������y���Y�/�v^������4�|���}���7$4��+z�Z�6A+W��p�&d<�V���μ��9�tEs��ڈ���7T!�����B.~������mN� �.λ��_�r}��$����m>���0� �٨zc�W��"�+��k��t��,�u�D�Ln����Rv�EK�f+ܫ�
�2�^8�餜#$��'�B�H�L3r�� �_�SJĪ��DOe���@70Y����jd�$=����֢;h�l�G}���2��Z������zm���}��RĠ[ �Zy�cO�d �k�y6r�����ٯ����-X���Y6�[�(��'a�ʲ�G������BOgb(��(��j���	.��I��u��A�^��J3�b�Ȕx�0�q���th�`���ڨ�'�E5��(��5�B �Ť|�d]�5���2�u� �����-!G�$��]�%0@���3F�}���4�Y�\+qq>�~�#�"����j����/~v�.߾���<�v��;���e$�D�j����=����J�-޹��Y'�᯲��R��)+��[�#B�Z� ��\9A���y�C�ؒ��H�8.n^���s&=DѪ��7��c82+��@��~�u�I�\��|;
�}L��``���0�diX�A1��,ZN���8�4�h�VE�/���z�i8��d5�!猆l@qPK
.��]��P1�F4G<��V�,s���β�I�,�at�K�]�i���8�;P���b+�^����f�&�6Xc0$g�W�YA���V�C�����Vs��V��H"Zž"M���mt��Цp���	/1O ep�3���%�U�'Ns�N_C�VJ3��UC��yK1��g����㩽L�#�(�3��L~u�����ʻ#��w�U�ˁH�e,�{��Fה�`�z��7Jm�M�*O�\W�a��Hl�3%���k�jS���.���c_�4�,�C]�(�IMP�Tʢ���_�n-�ZP�G_?R�_\,�I�d���@.W_4�o�mi����D���Z�.�+�$�!w-:$c�8[A��v6�-~���CMp��U�\�ب2���Ѓ���/�]&(��k>:��A�}v͖��h�J�X/$�
���(��ɣ\�tb]�(��i�*�醇nuh-v�Nn�L;���Zȋ�Sw�OoS�^�s�xV�H��D/�%D|/���o_	 ���f��Ë�o~E'�;F��z㗪L�$w>��F��`k��I5wA,�\!M�4���aD�����L^�js�EJ�J�"4�h��cO����d'LWr��	�m�.��E^V��ր3\Z�IE�ݭ6�hs�?����Q���Ն���6J���f=���6�A���W� ���`3o� 	L�s�=�5���t���>����yi��ݘ�W]��4��U�6ݾ{7�XA����9L����=<-���v�Q�lX��21�\߈�O(�%[:`��<8p���5k�&l�����0���|�JT0"����b<�T;�~��7�X|��v��(Q���\+�6�9.oac���o�֡��p9���TXS�=�~Ai�G\w}~�+�z�+��D�}Z�2pX��Im2�]�?@�~A�]�tۻ��(�iX�w��x��"�����C� ��/i:C^l���X!��o�k�ϸ�M��c!M�i9s0!�SH2�H���t��xKD \ɖ������Eaj5E(���j�L�'�zx���X��V?�xp~Dh����޺�;w�kƴ�c����3(Q����j�T���WBY@O��+�»Lc!����"7�6�oC8���F����+�E�DV�c��O�)��/z�\p�sƓ��I
���܍@t���$�o]�<�*��IhJ�Z	N��~�"���X�7%��#�ȳ'�SN�5�A#6�U�rʆ���)�7�Y�Zg���f��̶�;����(DY�����t�&O(yk�?�y�E$Y����C	�RAlD�V�މ}�2	`�r��
2�Z�b�1p$a�`��"���Q�6����YZ:+4�?���t�ݐ����^�Ɖ�o�^��߽j=!�ʱ�y���z2�iUX���K����y��9�r��Ր�2}�r�~aܼ�\�tPIn�t����JӅ��7`��Z*��o��ȫ8�P��g�#,}��%��mI�{���HɆ?�MH�b�hQI�*�u)�⪱�_����K3BV�r�fF{��$!�[G�~hDq��G�#�2_3Lʃ;5͹�ᦫ�aъm���^R�G���|9^��,�#�F��R�"o�H�+�����f.=t"N��E_A� �Hxt��yϿ��B����f�[7��Ւ;&S��`+�"-|:6��K�uۮ��M3���
��Y0��4yOU��?K�@�GG����BA$�>���D'�G���84N�����x�A��s
t��Nu���BLH.�=Q6�.�P�f��*�ڌ�]Ίt�ſ�O��9��&%Yq��W����Y�OYM��?�����#3ހSg�͓�֯��ьff�&���0�{!��H���P
R*����12�{c���Y�)��՞AI9�)EN=ٶ%.c,$I�r��hf���p�|��@��Ku�OaYus|4��*Qu�Vt�����g���K����	�_�;�Fq���.�F��܅��`q���Ն�GkO�=���~v�vV��^�Vŀ��?u,��1��w�����L��	Ѣ��y�+���>�My�T���Fqe(�@��"䥳^O����ɴF#���[�.��|��檾y�כ?Z�Tp�3@������{��5Oo#�è���N�l�z��c���3ZRb��U*����\!G�үa#��j:�^�k�>����_a5����uq���Mf쫂��+<�o�@���ä��1����!���|Jc���n��x�Ì�3��\��v+��<��K-Yx*��~��ڔi7��C�͆���2����j��\��\eڲ]��'�w���i�az��fg�Jw0ub�_>�H�?�}<u.7 �);c�<(֮zڰK��9�8��`S'��i�̥V�J �G��#[��d�="e�0�2w�nղ��8l�F�=d�����<���wz��w��!����k�Ѻ����OZI�Ǿ��7C�i���G,�S��MYj�$�6އYi�Zq��n�>L��!hE:�F/ 5C�_���q�
�jĺ��͡T,վ~N�3z|��z0ьvT���7�Q<��B$)�_ur����Z��$T��gu3L�J]�O9=��& �%���#�!���e(t`�J��rL}/D��I�;2���,�@iu]7�9+$d�_<�'ړ�����DV�?ۢq�d�4�����}��C�..����\��K���\�r�(����5�|o{{Q-=����`�����6Op5�B���ʗ�����`��v�@*n�x��ւ�*)�k6���l��+�	��s���&���2��K��_��-�8tB*�u#�.$k�����qG(`a�0��RGX��)���*�L�2WE�A>L�r 3�1����S�y�!��.M�g�S|K9Ԗ�?��{�1�X�є>�-�"C�GkdCu0�`_��T�nvK�I��#,J�K��ɉp������j�vy�6�<(�INU*�R�vbƺ)��!�T1���ʃ��:s��*߄s��~�W_�{y�}��V��ϋ0��$���]N��?}z&�0U|��,��z$DۄWߵ�ȶY�*٤)+��L��+��b�	�=�#G\aNx��r/'�����Z�&��Wn��e���h��f����d�?��P�"F�B��T� B�F���.�-��[���� ���V�v����$�2����Z��0�r݂��-��q����#7H?l>�Q0�b�)Z�$��y#Mx�X`ذ�HC����+�5�0�,��_�24e�0�'-
I�[v�Blx�������]/W�E���#'y����l��G,8U�n2�D�[W�+��-=��\�]��C��ϻ2J�mt��+�s%+����C7;$�״��G�X%��X\t�"x(��B���3�<{���6�����t֟AI�}F�Qe���D���$*��.��IO�/���礧�,�`��<td������ˏ��v_s>��Ut��W�4}�j�rꪋ������N7_���;ޘ���skQ�$ルRm,� 8��h&��-�����R;�+B��քlN��m��[��D��I�/�p?��?q8�1�X��ln/z�	i��ie��h̝c"]����t���.mi�5�n�.o���iH@=Ɨ})�3,a�9�@(������aV\���B��G�KL��^��n�3DM��S�7���O_  �A���ғzB#� ��-��"MK�+4�@��ȗO��P hE%�f'�_l����X�'B�&G��Q�/��E*�B�3!e{x��'��E�� W'�� 1�5Q��mᬀ*6�y�~�fk8,���������s��rl�����{��=s'��7�|�\0�2ڒ�g�[$i�y��%z��4���t�#����#^A�Yx�)nѫ�j0H��j�?��[��C����P���	���O��>�	�}��Q�R_�5w�![���8Le��20���4��9��CX�'�P�*@����������Z*N:���2*S9Z�%������܌��#�70��B6.՛
�,�\�gDWO~�c��s.^;��G4)_����^����S<��EH��f�����]TU�a���'�g�#w��;���j���B\a���AP��-_�46 ��G;�6�5�U�c�h���yq>ʾ	��+��]ѻ�P���g��H�Pw��%��.��&m��x���q���ER�o,��7������fm K79`���	d�V�B��uvE!r=����n�ֵ���ig�r�	d5�����9i��~zr��_<0�L�Ԓ�-z�����Pc^��HCW�%�=0�}9���o7'�6�@m�k��2�jR�R��F��d ��o���."S�\�y,�=�#�9l��ܩw|���&���ʨ����n����A��Sⷼ����\��V`�(��N*w���smHE(�Ғ�S��^��](���gp�������,�~��==]�jIмf���?$ȱ��tbE�-�ύ5]W�<FC�����ŧ�CE�G]O����Ts2E$������sS��Ǘ`9޹7w�ɤS�Q�,>��SIi�Yz�2�03};��}�Z��	���V����]��[s׈`��(>�P�����v0�o�5���Tky��9��孠���c!5D�sN&g�=�	��!g�iF	��&��Y���6���\f����	x�ī$ff�����~�q����tan	��U�9�b�k-����;~�P�}ٕ����U����F���,!��$ ^(��5�]�tD|���80��%�@h�A3sC���㪷��Iі#�qL6��B��Jƍ��G�fL�A�]�]��]����g�3� `�R�?m�����g�y����B;Z�4�'`�n\�Ʃ��7qp4F��-��E�Ѳh9��iW��"!C��|˙�m3�=�icC���/ݠ�C�Ai�1����,�!�s���o�c���jLzJ	c�T\������^j�0�!��f'n�I�*��4�SI_e��pS�[�_�)�mq&�HҍK��X2�~��jR�3V�u[���3��T��f�"��n��zl�f�mTA���@u�V_��Q'����R�e ��a�*H0�X�O#�@��O�$�͸\ς��̛��-WY�Dj�M���>�)�f�(8�A�Hcf��@	�f��Oܶ����b�(�L���L�%�<^t����Y���f��c* ��:�,�bv�t��\D�%P��s�:���&8q����8oS7���!6ߨ��1m���2La��	dc���G����C��N���7�Y�����������-d�7�L2Qf����|Y;r����uh��^w�|�C�4���3���9�!SS��)�z�(V����W�:��!��m�q�A��
ɪ�,ڝ��>���dHE���I��Ύ��âU ϝaB���ȣ��ܹG�M2+�D��>$�~��xg�P��#���l�s�E>r���s��� $k���-�r�n��8������ʉ!�ǝT��!��u�s:_��xJe�{����a@�au�ފښ����Xj�]������]9�z�T�*�ڇ��Y�%E�ѷt5�@�u �_
�Z�?��?d3X�Z9+��E�v�n�0*�,p��&e%��V}�'��8]�������H����#�Z�Ԅ8��p� ��'/t�`���f�E&��Bװ�
��bA�~��e�:Q�O�AEDR��5���0���'18�yJ��s��wO���"�~�J��;C��ȭsj2��q�$Tُ[<��>��T��Q
�:&?�PC�6n�˧-�M����{���%nI�s}�a�m��Gٹ�9�e{�����*��l��I�{0	��ۍ?�����u]�חC�+q}��n�#8K+;�`}��.a<	��:���~�������,�H}�����B=�_����9�I�,��X-/�):ni0��<Y�IÙ8�y}�ʙő%�Ȉv(�e .MQY�V��	V�qL��#��s~��
�oˣ
&�z5m�L�k_U�#��|'��!f#x���D�\��r+��S����UES�4���'�Ävv���ߍ���HH@ҡ�H��ri�����ڥN�eBZ��֦d���D��i�	�
j�3Ack/�zp0���v���}��{"RdN�p�`�o(�0��n�3>�"���ǯ��������&y5�|�9�s�O]v-�Ƒ�Z���q���餜vA,�K�[;�/y��t�������f��t�gUp93����ԅ��^��\/`�4f;�}��4�>��'��#��#����ֺK���D"��c>X'�t��bك��V�Zӳw3��[z�&�<�@���}�b���w�����3�5���7�޳��z��/����z�'��Tt�Œy$Pm���f��YR�_&��%J>��Ρ@i�z���]�o�;�i�ū�O�~��[ZL-m�74jvk�u��\��(�O�{�6��?����|�����Y��n�F���]�_�(�������E2�(DH�x�aGB�@��&p�Ggt.��t+�����Y���Ï��� �!�@4�k�BLp-s�~(jP/��ߙHU���+�Vߪ��j%'�Taif�N-�PB�&cY\��a�1�u�eU��}'�	�>n�6�n��S�t�Ɩ��M����I�m�k
W��_�"�'A�c/��O����S�t��tI��Ğ�D
FͶtڵ��/����$�`b5�����\��JqE���ƽ��sN��9b�z�g��C��ͬ��jO6�o��5�h��*D���Y�����T��+����ƊIq�du;1I�`���1t��i`�u4a�l��ߜ#��&XV�RC�3d�)�辽4`��Y��M��t��O>E&U�h�4�� �Q_R���E�	m��aO��D����h�e3����f:'Y�L�|U|bw���� �����bf=y�ؾ��8r�$"|��$o�>�ޏ9��e��n�p��)��3LGw�֪m`�����ݐ�膁�'*Hp���+:�ך��P&��XOO��W!���9vX���"u<}����$���4ן#yS��B$RJQ�̤�\��~fY�B
y.[�(��n3H�3}�	�{���`~�Ei cGD�p���-Y=�>�����E�jGR���Dm�ʈ�x�(N�~�X���ET�vQЮ#ݑJ���C"x���4���4�m�?��x=א��S�e�i4�L�����	���a[�؝�oY*"��2Q߭"	}	s� ���\���S�{N�I�ͪHD�@*���pS�s�:��*C���׹�uZR�I�(�p8>*�A��2eM��pe�W��3(����TUu� ���s�)$Co0:q�@�|�|8dc�G֚��&�a�SD=��(�� *}Wغ�v��p�t�(9���0(ݱҜ+\�A�&���hl6���YI�7
UǥQH~��D
44HN��W�^�Mh4]\l��iA��*����E����=0��߉�V��%�+��pq�J9a�?�����λԃg��S-�䞗u��*�Ah��� Y��)����p~�
��ʺ乬���RV6<�}]��s	#V�}B@"��]U�ނ�%K� ]Yl7�ࢼ�$�ޑǷ�U<Q�l�����*�L̹9kD�˛�綹|0�Ps�zf/�"+3���m�0�IK�#'�Y��q���o6��?Ƀ�(]swYrj�W�ƭl��.w����(��[<^��z<�1]��:���Z!q��)u�5�2%�U�o �gR���,T�K�l�'R��PN�m�x�O�i�m�3/����s=��X� *`�@�E�r�lO��&𻈡4cې�.:����8�]�mk� �gKZ�N� ���i��3ˉ*OF��b�s6 Y�B4~Iu^C4�x���iEZ�U�T�m�BSvCk�'ϫ�7��*�s�Jo�����Q߸�A�87��c�[P��s������/Y�)-j�#tl)�,��Fx���p���:�T'�] ��\u�%�4Y�}>��:��C(�3��@%���9��E#ޗ��A�����5�ɷ��C�R�����xu��7��+G	��%�B�%�{1��b��ɠL�	���V�9!���y�`�W�6P�<M�콿1>T�h2��΋S��""*__.�@����Fs+$�����(�b� ��SA�QL\)��Jl�O�5��v�����Ҙ�ɢ>���"/��}S�`��4 Y����Uh,n �](�K����u���ϫ�;cR�
�Ί:�QQx�W��b�%~%���1�Zko��ѳ��[ b��ܚ �b��$8RJ4�B^�۾�q�z�\�����x��Rm����9� ����߈�v����{��p�����#P~�v��^���M���u� ��ʯ<�EfE�A~7�6���(DEYrs@j�����ׂ��HX��(d��Bq�^S�&E���M��tݽ7�n�o���Up��[�а94�;Z�_1޳�.�b��4+w.W07�hܦC���ޤ�&���x�)���&N3d���^��y� �ֽUr��D�CF���� ���	��G��4D8|{�h�Ez��!��;o�똹p領8�gK��"`M�<_扱�h5�����c�y��1��r!�?�B���Q�R��(�a�tYؠ;K�7|O���L�^ ��s���s�V\���a0zOu��(���+3
R�խ<h&�w��T�϶,���|><�+��
L�%��O�
 ��͚M��\*�b�	�=1��[�h~(�V�ዸ|�"��x��N�m"8l-X������n��o)��W��܆�m��CK���P�z�0�D7xU��&\�����:��6���_=ڻ��<���=���z�}�nx�_��9�I��
~Њ8��,�̓�	�A��Y������Ŗ��"�م��T HCv�Q�	���0ףj:	��07�߰��֊k�� ގs�j�T���3x���o�g}�wf�)F�rL�cC���ݮ��݌%��ȉݱ@~hc�MB7��)��ǌ�6Sj�1~oҀY���4ׯҺ0�*���7�E��F�>
��蹪Z��&����:�*�z����EnPa��~}��*Z_�"���OvA=&�����������J�X�GRޛB���|��P�FAh��C��"8�NPÌ��ʣԺ&��K������2@li;V���ɇ��j�n�Ƭ<����J^*�۠9�8��}��žB����ݞ|y�yO���j�_x��L�n_+Y�Ix)�t��)���J�6�i�n�۸� ��b���&�A|�d��K-4n-���W<��$[��{�����&�ҟ_��.��:s[%o�|֌�*G�G��5ǚA���1�i2��|�#5FL�����1���)�B,�ԧSe_y�L�x5��j�d]4����!X�[� �X����﨤�:5��ď���D�~�)a�-�0�����x��!��33�~�}���!�%,�e��� Q��b�Y��^ҒHK<i�/Js}W���-�c�7-�?���|B����Q���~0�w� �~��z;a��}n:�Y�;]�0��i�P��`����S�;Po�Ktp�kݸ�uBͭ�b+i�W�6������ƭ�T��g�U`��5�V`�Rmb���R��g�@��ӛzr���r�}j�m�r�J��rsDx�`/T�7ԧ��W����*��>{�W�:�q*Q0v.����W���*�2����&-[kޔ�PP�nϞ�fu�mXt��do�P�@��[�>���q��_�[``6$��Y��w���O0�a���Fo8��I���q��gvs����fm�}���~�W}n�O^��Mo]S ��-b�'�"�k�p��DE��F��>�`�*��$n�W|ƜU�fw��y*�*^�=%;��hV���ᥑ��68�?d�^����#]l� ��iv��n�����i�a�T._�tq,�M˚<�iY#���.�A9n/�`ևx�箼&PeZ�8%��׵o�l5OC�6���rB>�ۋ@�1w!�.#�q�����L��î��4�9�4�D��2Q�ޯ䝽[��'�s��Q�v�W�m@w��9��<]��̆?'.����Iē��vb[�8���o{��ө��V��-}b�*� �V3L��|x/�5�i���7>�[��C ���oGp�����]i�j3#����X�5����vV�%8y~��x�
���$�����㴇(8�����n뼚���_[��[M��E.�����xʿmX�1v�/����c \���ܺ��� h�q���pƲ�s��̴�xU��J����DX����CN�	Am�Μ(6#-ġ;i3���
���>uNX�G2$3��YG���Vh�*� r�Z�͇����?Oᦦa)B�`e����}6�2�)2$�":��Gg���漙���j������}�
 �p��sr~�;���Bmc=�S/�}�hJKW�-i������Wk�@Q�(	~���}dI����[U��77372��s?uDg�	'VŜ�������к�y�c��^�	�^�c�����=����h��S��p�5,��>F��2���h�"c+%�^N���h��"�8ӱ������c�<>'?���x��u�=��uK�����oX��h�������/�W�Lofj>ź7�ͨ��V���z=�9`���
���I��>�v� H�� ����KbQ�W��N{�hP(�������K;�� �!��`���:��O��PF��mYfvZ�8l�m�����Ԇ�`���iU\���Og��&�M*nG}n'/I�CǫE]%�鹺��@h`�D��;�e�6�{�H��ں92$�%F.O5�Ht������]��;e&�չ�+11R�A�Ld�3��5~{ǻ-�M����YB���5�Y��b��ќ&)/	��v�=q��r~��̝э�
֒�l��	��ME��Z)4?_�����^vN���Q������ܠ���5.����@M5�WX	ItI��j�c6Xd\�)-�R�gfj��i�C��~�TJ�,�ӆ�~}��W^����Ձq8`:�q䦋Z`;w�R*�����H�lnYY��n���=�CWz,7�Y�����\n��!brS��i��C������xoP&���7����X���2)/�
���N�Zqa�K*0}��_�ƀ�uo�w:�~����t�J"��Un\H������LJ��0����Q��X�l\�1��m��2)�D��X��QK�Ҫv4��o�A����w��40ʹ���P-#���r�_�%��^��
�j��m`�:	��!�*H��=��NI圮��0��4�������Փؤۅ{$(j'O(��nVwp��5i6��]��N\L���K/�!��[%���#�Ј�rf�s�4�A�i�A{?�C��T�͊Q�/�C7�w-�;P[���������g��r�&g��@�C���p<^aa�͉��y��s�O]�l���PT�df���FԳ?��ٶ�RB�eP��"@e����55�/�=������������!s�H�I�e�?�s���	p�)Nɐ���������ˢ�p��$r��j���R�Ю����j;��4T-�� ��p9
�.�Ԇ7ǒP2�w�Y�v[Q�v�x�rި��� �ū�I筶��v�nHnkQ&B�U�hk��Ki-M]�cc\)>s<|�1�H�m	9ƞ�Ν�ߓ�eM]�WX�D�i|�I�y���.\ѽ�$�j�p�ɵ��ꢴ�L[[����Wa�DSS�O�a����u�e���m�8�hJb��#�a�Fϑd���VW�4��BT��W����0S핂�P�6�j_�2dY�:�3 ����<xr�
	G�)e]ŰM�l����k��
y�r�\7�� sA+'�������.e?g��h�cQ� �7��j(I ��h{��W<�嗦������}A�5cGe�i� )-��6��������P�	�
3kX>"3��a�'��*���<��.�ת�,2:�y�T��)4�w�lMD�pI-H-oШ^F�Y���s��_P�k¸�E�:f^����x��. /�G� �@���GM]=�Ǥ�Ezw����-[F@h��$�Nl��!OK�TO��:�V����pA�� (�W]ny�z�`�oV	-�2�9���yG�QQv~(H�AN�	��
�Q�)�ŵ��q%��*c0�d�U��.K���V�~�=�O�N\�./�B݇!�WkN0%q�gp6�bC�/ �:���/�ji�� պc��u)P��9r�BnȰIq�v���I�E�Z&�.�
�J'��[��w~%�R�y��}'np��b!_�c�"o����+���b5��G��txrNd�M����x��~�k� �����4R��Q�~އ��p�9��ڽ"�$%��c�R<��}���sS��v>���+#Uٸ��&WhZ��	�
�� �L��9흷5�٣�7cmA�<10m�D��}��N(]ҧ���� ��"U�P��)��4ۢPE���5���Ǜ�1wWMH��L��!���>�����B'&}9��g�|�����Q�%yͬ�GG�Jqu
O���h{j����(��:o/�0�	,ﯟ�&׉k%X����G�?���ZϪeύ�����2@z�����|v��3o2���d7V	ŭ�}뀋��^)�"�o���a�#�د�a�^�d����V�79�m(�ԭ�����f�C�y�MyU�7�0c
΋��
M,�Hm�/��%�r�����D�����5M8�@	��O&1q����K���H���Y����JP.l�U}٣����JuJ�]d{�1pPEa)h}o��CMo]4|�A*�s� m��c���}�\0�|����eq�tnUOo�R������kFu۝�����KzLtC+.1�vm}�O� T>�u���;���a�����X���'�k�d�&�;w��� t%1�q��~�������ɚ���
֪��*%��\f�"�i����^ڦ���U�L5���C
��S����ҸH�� �~Y�A�<
�Ò% ����i.�/�.1* �$O7q$x�B�}	��B9�C�E��V+�_Ԥ��E��P����u��@>F���_�$�b��UuNA	8z�������"�>FF4�E�_�p�|�eo�`; �o�.\��� A�o��yoY�KX�����%����H�N��8�Z��l3*���ø�x�l{`�5����xseq�mZ��a�i����B�������Z�e��b��i.��$ è4I�8�@�k }�s�v �d�By��%�Ґ�m�%[bW��;�)������[q��he<0x�w�t@�5������Q�+����9��3��䑀�oe:�j�	���xQj�M�ͮ4�^Ӑ�P��-��֝��&�S#��6�<~�H�Dm��1*��H��O�|0�Q�$͈a��O~������㧿��d8ک/�_lh�	L �&�v��a�*vݗ*�,d+�v�L��q�Ij�̧�	��U��M�cMp(�!�-+ζ)����Џ�1��UF�fj]��� ��Z����A�t���9y� n�Wn���e��/��F��+ֺ�6H���+�֎3�|t-���	;�l�L� �{��ѕ��Ԁ�y�?D�d据�*�O��Y����j�q�����=�p�y�S�8%�/ʍ	��S��_���ӷ���[�g��f/�sc�}I�X��r7��ǆ?����������K���[h�̿�ݛ�s�qd�;��I�h�F�[f���x�b�~���eߪ����cbNc�x�D�	F�9(�����cM�_]Ž8P�o�1�0�H ��?�?��@��%�[��8��,TTE<�:f����ڜv�:�[��I�|���+�1��d~f��l%��x�/�k*�+݌kb*�:���"ɥ�Ͻ5I�N�z����|��4i���	�))�/eSt?��RU��	?�GZ|��=�D��gª��6���� Olz�R�O���U�����Nr7{Z߶w�ʇ.���;4�/A�;EI���{��RX�>1n_<��@�hB�I��K�����V��:���5��3��J嗄�w�R�"&ĳEbIt���,D�բ�H�
�}���<1�Ό<^���r{�����<���L�v5�<�q~���J9��ޙ��7�n6��W,����zlIB�>�n��|�+Dq`
VJg�+��p�w1YB��n�İ�Ņ�]lf�;ݽ�^`cF���YE�ș��W�r1�l2}_�2�e�N{k;-YrK�k6�aLx�+u��c����t����Lm�& s@�E�����%/��#8��__� ^��8���}�j�1)��a\&ةXݦ�������ս.j\��6<
rWPՆ���.=�Ӻ;C��7xQ���� ��d�g�ʭr��ƪf�I���%Uڇ�$}p�����mq�����OD�N�[V�K��
�(���zMgH'�>����P���-���Eц�&a�c��ss9�Y����|�
η����;�Cu(ZOzUH9�k�4q��M�3���~k؉�S�>�N�Ry4��UE��]�� ޹4N�l?�w)h⡳C��N�%-�N�tx�\�-s"�W��Vλ���j^��-�ʚ6�w��I�����ŀٝ0����c��ƒ�VO��{A��΁Cx?������y`�g=�%��A]>C/�����%� \(
A��/<���F�n���L������ɀ��/�� �	LV�J��Ӫts'�r���B���+6��㛸��������q�jX(OU���\7J:/�2~-�����^;��BG�/e�l|��@L�1~�R����e�:�q
����C�������GKh�����)wI}�c�+g�X�Q#yR�w�|^�L�(����h�O���0���� �==gF-+߄b�����Ǳq%+!"f�۠K3�s7��H�f��F4
6"��e��C�\��b�c�Y����x���&���6K,�W!�L�9>s!�d����bݜ�{,�S�ۇFn۽I�:��6���΅G�,�����tq�����Uɽߺ���Ct��t/�~� �2�rT�[����(�=,��Ly��#�^
7��;m�ǜ�?�	)~pv���>(tpse�Q=_Ҁ_RI�;U��얫2�l�ܴ����ͭ����r���r��(J{��W�v�`샠���K��y՗zJ)_Lr�^���3��JM���z	q^nfҤHF��ڏ�X�_�\?��6;�$��CI�<�(�O�z�7��藖�Տ�p�3�K��<:���_����z<㼓 ��#�Gik,8�y�H)SF8���LO�Dc�
|�e��$U΂�������O�}�E�5n������H�Y�?TL���g+@Ŧ���#�,�&.j�L�P��9/+rW��sӃ:V?>���Q(�
���ƩC�����(���U��9������K�W�jA��H��F���4k_�(��
���c��>�-�6�h�Ք-�n���U�|�b�
��f��|�v^�.��#�߁o��VM��%���:�u��߶����1K����Z��tY=?��ΗGZ�(�`���tG����/nK�迋�?4��L�� ��-�VN�� cI�/�*J��8�"O$tM[��|�E-�z3kc=X�VL��`�G4<�ܾ�vID#�4$�e�O�����V.��N7Vay#�r����"n��(^��Y����W�?U$�Qpm�;G�����%w���$��R�����H�*J�rM�l'��N=�|��XbM!@��bYy-���E�{�v�p�fX��%^6S=;������NE�d@éqBu2ja�]�_��6��W��zr�h�a�/f�?$S[�5ѵ7Wi�O��h��x1�5�I��6+GV���
�S�nMZz3��RL�A��ky��W�℁�:߇F�vq��x7�T��6"a~k�Ð�giJ�3g�?�p�՞]�h�Y�L���N��q�������D�"�gn�j#X�X���O����x��v8�h��	��9�s��|���c,�����}�mNq���pݢ-����8�`V��ƤaE/t�@��
S������)�mbe*�|����i���[�ۅ���P��j"�n�xoqN��u6f$���BJ$�v��.����J�f������f�m����a3iAg_�_YG��x��]���d��Q�ˉs�'��OG��)ҫ�H���U^oec3�ǋ	`���D$��҆��D]�+f�%��&$w#�*6�%R�l��3���]9�:2�M�.Z���u��!�Y��e�(��hRJA�C��e�L'��]�m����-d����c"��y�-��ħv��M&�t�(����(��I�V�`�������^
�;�nT����]�U�O��N����VOU��)Z�9U���XR}@�Ɔ��%����Kr�|�"}��������9aҟ*����������5,����A�l
�S�2�F�|���e'�-�#4����G��"�/+J9�ǌQ@��S�h.����HQ�?-�M��H�`��W  �&�~�	�b�·��lC��l��2Gu�b�9�qv�7ꑃ�2k��+�J��)�D�����aܷ�/����hr���m�"4M�En-���\G�m�{$�Q��| !���f�� �g�d��:�wԢ���;O}�mZ�@��γJ���-�u�AlU�@1����/�`I2���۱T�y����v�S�-�i�w�߭f)0dsU��N`�F��^$��9���r2̦T	��C���6���ڤ��/qlЃ$�\��k�1a�5�M�|�{����"�~[C����M�U}���M�Y3�X�n�5�ޤ�	Y|��L���Z�WR"�ms��`Z��pe��ch����o_���X]pR��>w�D���3�c�7�8��"/��(���#��p"��	5_.��*+��^ʂ������Od1O��K}�N�95{�v+N΄�(��+{��9�0�m?�VY�k���������E2��������J��P���SDi����'GP�g�l�h�(�A�i�9KN�^'h}zR�gZ�-[�lh便��N?�K��ۣX���of_�Qv��¸2�t� cx��3��lp]�4�
6z��T�Z^��l�
��mo����*`�u`�ވ�L����t�3���z0��!��}���yVv���C#2�
��7UdA:Ve�^��l��+m	��NK�L��h�i�>��������\3;���I+̲m��U�ukp��"�x}���^����56���PT]g"���H�4t����6�:��!����`P������#��~���ZQe��	Xx�۳�&�a#��)�r%T8�z��a�����H�K4a2�V[���rn��<6�\Z/y�vL���{ܳ�%آ8��o-<^M� �E�4��=�ˬ����a�RK*=9�C?.t?�����,���ur��k�k@Z��K.8���#a$k���W�hd�.�}��Y��8�t�fq��'j�"�q������R��A5IM�j�I&���sQ8�$��,��g{�A8�,h%-�݁tJq�t3
DH9*)0����6�(���,'ؿc~�ŻLCK�������5	F9�0���G���/�0 ��V��-[m�P01v�/�a��N.�.��uVJ�2���x���*�Ms����{{�+�5�!K1Y:�XPQ��n�4�Wx(�4������z�J�'ϧ �JFD��@ ����VF�؋ĬO��^Vey��%�X#�Q87D4�A�f ��x|��00�{S.��GҶg��A�f��J��=���S�&�yS������3[�F��6���B��;&�H�^F]kyzK 5�bE�����8�3����)�0�>)B_�}<x~�������>�tA�y"���|s`1M�2��y{������Yi���������x����,T+ i�n
�0�p��Q!��M9�'OlG���ً����p4�*0_&���KfO|��,����4�����{���%Ka�q��n�5������wo����O�{��Ep���E.���F��N������l�aFU�:"�m-�7�QQ���ͪ.�8*y#����5�}t;�s��$�}0�sjna���W�ξUaU6�;���f[�A W�}�>E��l�LNӛ��v(񫗰Y�7,�sy+p��X1f�&D��ɽ���|�S��F���N2���=��w�?r��y�����T�q���^b���0���Ӵ1ǲќ���v5;�8)�B�K��̀I>//�g��� :����c{�d)���S1o�h�����]��䤨�KJƍ*1���R��j�����T�V��0d�'�HM@^��?B�_�F���A��G]0e�D�~jm��H��X�4Ll���r����>��
��4���Z������^8�;���~A1wx�=	ũ�G�d��	m��5�"��-5�U��SJ��N��w�ӹ��GI���3{^�jL;�f*��>�hp�7�fH��CCzp�����^�\�c9b����>�)&�Da�� AY��w��d]�1o��s O~�yP��}�U�6�/°�)�������`����7�s���t��l�i=�6�������<���9O/��еA��;FH0%͜O|fK,M"��7��3���z	~�MKYpNm�*�}5&3�KΏ,�������T$P���/צ_f:�Ż�����rR�"W��Yn�)ɷ�7��� �1��j���_�#�[N�_;����g��@>��th76�������x�������A���tF�ӗz�\\�=J'Bv�$���&(��5��sWG�-�^D�=�4��;"ƿ*ӏ�˟����/��J�˝kL>�pa����0R��r&�s�R�yKW �A*����(���|�f�����#�	-�иqK/l(I�S#pe���4���(����O�	a��*���*/���u��u��jܼP7���}��W ��`�nO�{T�{7U��%�{J��/i�yY�"�O
-e9.�����޳���ܯ_���r�{3:j�e~0u�OK��tPZ�H�
EEt��t���]�y��04�V)'�W��K|qZ&ueh�"��ʓ\�e8lj#Q�Eyu�k�S#�>U�4��\����)Z�����Ǟ���XV��܄�6_eʚq������V�Ե�����g�sL��|!DM߫��`�'7���x�F�s��o�^g�Jtc��B)x�r���7���.?M��\�-�]���j�<�}�^�Qc�d����~��u��2��4�0��o�$b�pN��Xu�m+藟�ZB��c���9E.����5̥V�ǀg�6N���q@��)��N���Z���h����4�J��k���181�ַ�P[[�~7��ZP�8y�߲���2���IG���kQ��B���o��\��n��q?]G�%��'�|��fj�Cty�� 	����X�۟�-��c��4�FY�}4�����*=�A'Ɔx�:JOӰ�*��k�-��E/j/�;ԍ�	�Ř�ӝd��j�v�1�C�*��;3K�	<���lpM��u|���:䈣}�Z�Ȭ����aj��b��05��t�5�cf
�Y�,��uQZ���(��olM�$�gg�K?_����>d�Y`2��U�:���7�")=F@Eǉ��񅲰��!�����A-X'G�VU~Õ*+*�ᔑB3��B�LG�p)ه����[�JM�c�� ��Z)�ŭ�3��!�M�*�ܽ�1V@,P�?7E!۾_ϨL�o܁��/R���ץ�}�Mʿ�9���Fcu��yW�d?�mED	�:p챦��a?5&2&��$ ?���M��{�N��SÏZzWA�q�^��(����*��*z���Q>M"�
�R'	����rd�I顰�`B���5�#lD��nQ7�5���5��O�u�:�X��(��AA1�#:���@`Kl�b�Hg�{��Ҝ��������^���f��i��7���?d���*�B`�O��� #A�ٯs�
i��9����:� 䂨��Q�Z�WS������q�,����c&�랫x�r( �/x=��_ՈA�&"�[�d��o�Rp���_�;R?Ip�������:���6j,[wj��e�6����Sʭ+VZa�X�p�]�]o�����ʽ�hpa}�<5��K0���Yx \�+�uP�u�q��mZ�2h�P�ODp�����rX�c�0o�^�]�t��\����%�^_+�-M��2ެ�"n=	��{Fw�;�q���x�U�
�W����^ƪ'D�nLY���2�`ʿ�	E�:����,�y����k��-;��!}0���ȹ�PpG�SOAZ�$%@�����N�"^6�]]�Y*@@�WI	�r;K8I�)D�}��.b�*-}Oc�~���-��j�GRb�����V�c�*�R�GQ��A���'���7�
g���@��~K_����;��(I����}��b�L1?��	�P6p32H�攠�����C��m����2��l�1�e8��hz���w�����P�gb�ʼ�1��g3�������toمP#V��S�>n�T�
��!�\S�����h	�J��f��s���Gʢ��y��Og������+��3�=�h� (x|��:,�F�;����"/� }dO�m�`Y�m���Vrӄ��i�c��2�/���Z `��:U2�G��ʉ�t�0/�/���F��WU^v��T1ܕH�di�5����pSi�Bn'�n�o��U��6��/ 3��	��%�z\�l�g�0Ջ�h�h'K$�� ��� �z0�?�n�pY�k)�L���Gkh�N�$ۼ������>�����cszMͶ��;�ky�(�
�3�Z�]��v�������h��g�-$<(B�����n��Z�P��|����m��ڹ��F'![��=�� E��<z�+��9ݱ���W�o�(����%�]�S'p��K�C�� ���0��~�W�=��+ٵ��.�D�_U.v�R�n���gb���s�֏��a,K(��*T&�`������'8�^�D�:.�5�W͖@9b4&cg�L������"6�$�Qw��Ȕ2CbY�9[���>��X��1k��ҁR��D�n>O���JN.�0� .��u	%�;�6��cT�R]J��*��;�Uޕ��r1�):�.�m/��&��K�������>�*�ա��{'��2��rq�Ǳ��#h������
J&�5�-�s��c��������ʟ����Ž�J&�\�8�7qA�<0��$�!����AT"4�6G�W��P����O���I��E���O|��D����-��*�ct1�gY;���F���@\G
��a���-B<,�����2-���д����)��jJ��F�Pe�K��x��S�B�&uÀ�t�����2�`��=~�HҞ�r�r��Q,�o�Of��Qh��l��Γ	uw0�2}<��Ѧ���3������6��4{Wg�fHY�ޖ�o��)�k��G���V�-� �Y8j�ٔ6�Owе��R2���{���؛���l	��)��A��&F!����6�����WFݰ�DϤ2��X��ѐ��a�����w��� ��������Zoy�Z]��rL�3��������01��S2�ُ�rYX�w#���L+#�̾J��,(-�2h<�Ʌ�K$ ��*LF���R�"֖c�����e�s}���l{|*�x���a.��܅E	Z���Su�*�ฎ{�rԡ�l�I[u
1UHH�qxx��I�g5��-�*��6�m��kva��z�; j��dT�����ʅ�Y��k(V�r���� 4��Nkc��T���%7Lګqn#`�����)�N~�о�ՉFqB�T�i'�?K��S�ըSG�0�4I�0�*�9��3������}�H��f^v<-t�&Ļ�)�ü��S�&�������敛�	���P=z��9c!&,>.��"Ղ&=���U6��3��;��*E<��� �3]�NӼ�|�����٪dy�Y��sh
�m��6,�Q_�[̰��{����Z��"�'�m�Hc(z���Y?�C��C{���Yq����m96?�2s�l:�v ��N:�oY�gP�HT�P���R�����d�y;���S�Xn��A��-���>������8X�9�7����.R]�!H��V30L�m.O�z�a*�Zq���v"ީ��I�d��MnV�oq瓵%9ټT�\���NA[�R�_��e� �ø�X_���8BK$�öKۨu� /c�u����.�!���G ��/���°�KS����*�ݜ�@j��*���Ԍ��^��F�s��P=B�|�����V޳-����9ѯkOn	sG������2�Ty�5⁂}�j�j��^fY������.�fU�R��a �r��Ӗ�56|xE��?�r�R9�.����k���]+%�z�����:�dB��h�P3j����1��"?¡�2�A�����o�5l㝽 �ieݐ`�QM�Je�w�b_��
o���朐�o	�&Ԗ��\i��LL�(�1?�хuaW�$w)�E��o+�2�-��#���q�+!�V_-�g&��x���'���
�.d-k~j����?���dí������]�1�Z�'!�M���Z`�?op lH[���S�=�H��#c�*>�W�	P��M��$�F|OL�xl1�2/ms_ªj$������j$(*yK��+��[�$�#��L���ԖK�g5�S���aD=|�l�M�6kGCJn�K��U�K�^6X�S;o��DQ�7��S��ze�X� 
|?�{׮rt��V�e2[��֦��[�tWd��-Q�wQ<Ci�>�)Y	�,�V���#�����^��b�u߅�����h�~{�qW�Ę�8N���k���c<����I����ǚ~��#�m�C��Y��R
V�K(TBN�]����q�`,5%������qʨ�9��%����^Y�ή�C�0D[����;�_3Ж1Y5�#�r��_�Oi-��4��`�Cs�_je� �ޥ�.�����VC�F�T��ԋ��6JN̚d��p��vK"p�/��~����z��[����:6��Ll����nկ��[�Y�`
��͓��xp6��;��禶1m$���TbZ���C]�)��r�s�����?��s�"�M�u*�"AQIT�ȡ��9�XBoO��Ӈ��/��'�\e��!P�5���z�׵0���4��߰[�(��7�e��Y����#p7�ܸ�	^��]o�=t�����ˍ6)+�ʬ�pE���r�*�����p�=��4َTta-^8+�3�}�K�
:Vz=�S����E��;J�ge�zi,�V�`Y���\�s��>�[��!�2ĞKC4��_`�	��ѝS�n��P�ϋ��O��"�k�dE.`2����9D/5+L����BP��?�vQJ��c��]u��>2,lн�\֗���7꽫~v���V��l�t��zȈ�����0FGwR����^J����\������9�eFȓ���klR&ȁ�]D�:�C�A��A/¥�V2��Cey�M0�˦Jmlyթj7�c�w����=l�yp�W��43�/Nck��"��=R��ieĳ� ]»�"Yuf&|[�H0�y���ȣH��a����mja6�Go�:}69���M�Y�~~�1��乖�����&^8��f�h�A��1�jj�����ٰ6՞8t;?J0�;�!��CN�&yY�f��x���(���-ZF��	�[$����2��Y(���-��.ᚂ��<NI�r"Fa�	�7Z>f��2�Ӌ]�Ƞq��ep�&Rg��>ɩ-H)���b0J7���p??�ƤB9 ��>�6��8v���1,�� %!���Sc�?k-yB]��X*��=,&����pm�	.T��%|��	`t��Ϭ�v����)	�`s�d:�w.@�[�*��t�ŕ�FĠS��j��
D�/B�l�D�Z(�;�=��[+�U��Z��t�=��8�W�wK�VH$�[�o�����i�W@73������8�t�QHTb��O���*�b�,��JOП_�()�ː}S�����}j�WÁ��a���#��=R%?��d�Ë5�G�9��y}��H%`a�� H�)��gя��d��_�TW`! pN?_l�f��q���T��a�j$h;�M�҈���:1=�#�!�'�t�Ȍ�Jg�Ɔϴ��X~z��8N��Q��~uO�T�8�Iɻo�T3��Τu��l�G��Gr��.�.-!�ӂ�ѧV�.��36h����ٽq��n�.��7���������y=R�'�נE�����X* ��MZ��Z�9������*.���]���p�޼6�B��X���|�3��w����v�(��*o�}�]�9�s^�7oEDv"�x�#���u��}O��d	R�7@ɜ�\Lof���|G���ts.4�#{L��KyI<�W�'vp��#�=��&���~M���E[���@jtJ�%h�ĸr��_��m�`7�=��Fp3&@=��??)��6�!v� �'IE��b�II�"���MI��k�+�3>nЁp��$��0f���y)���툩�7��P��/�yҸc	�I��}յ�?�@<i��x�[%� �k�Z�3�3V���9