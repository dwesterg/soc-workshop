��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>�����{I��v:?�BÅxJ�B����f�d���n�,o4ʣ�Rd2V��&����q�B��$I툒GM@�m��O�+N���K=��~���y7���{<�����(�Q�4�.�����BbLS�K�,�ݡ�&-��-��L.}��7I��L�p����U����eT�O`(+0�d����GK �<V"=����)��*������/����PY[I����n��l�è3��ML����59�ā�#k[y����%/�7��� �>�Ĕl��U�22Π���&���g_@�0�.��{�a�SE����\��N���h$������{��{�_�Z=���bxK&yd�~�����3y��4�g`�n��XnČ�:�gz��@����&�f�f�'Y�b���Ev�ҪA��N������-��AŤ��u3��T
St��yN3�Ȉ���,�jq������,��/�� ��5K,������6���zJ�!X�w��5�F�qS�������<��JY��-��iu �F����їN�k�%�é��z�L��� H~\� -x���ҍ�h���~*��!9�X��
��{�`�j,���i������tI�C4�abnh���M�?��f��;L�h���%IgNLVs�ѥ�8�fr
O���J\�D��@}������YY�@A��<��r;��R�����!s�$�2�hƐ9ql� ����k�I��ֹ�y�_���.i@}|6r�ޘ��wv�bd�N8 ^�G1��G��3���1�a��D2��"S��I«���	����*#٥�����v5�r��,ѵ"��X�������y�qK��>���q���i�!�=����O�^L���v��P��,1{��*b�0��G`-�?��Ү@�Dv��0j���<��3�O`�	��}�s]��#�Lj#����G�f|�z�]_7,q�� �}�h���~�2�8��ϛD�
����;�~���݄2D��.�o=���_���a��SV����_u�3�}(�!�l��t���A�,����kyO���#�xe�*ی��V�V���׽��T$_- � �/j��H��;PJ�h����X`=MS�\�%�u�B����V_t���;dV�	TŻ*��hy��2��~Ӝ�G�If;��?������ןȮB��M��+��kat��w��%�HVU=Ĳy�B�Ʊ����QP�V+);�)�ʦ�+$m��M�a����D,	�$ĕ�L�������.���r��$V��؛ۍ���6?NἩ��3L((]���vF1U�dp����D�1X�
��b�i�x&���2���OvZ?M/鰔}��Jt^J�ռS�~��!*�}X���!�U�?��!�%VHj���^U��*�����A^	��$�嵨�N���Ma�zOĘ�b
�c�DKkCX���Fw���)�Ǽ���ՙ�6���������&$C��V�!�k����l����}�%T��3�*���:Bm�3�~B�����!�`��ބ��Z�Q�w��������?~.	P!��5$�P�A��g��vM]߭^u$$�u��<�yԠp��<�@�R��s�!ǟ�y�V�s���>�m��H�S�>Z�\(�w"̰�8X�<b�>P�f��²��2�h���ҁ���u {��}�&,N�7$�Zr��r���˘�'��)xU��l��s!�d1^E�T:hq�r	��&xb�/pS��F��W�S�6E�v��h{�Tv���
okfƝqG-2��;8R��c��w�2����>b���@5EI�M� �^�J�OMs�8�~��ίM�z�!l��6��݋(����>`�XI���2��E�^*��=C4/Z���16�-"�Z�gktm7B�����)����w�NӐ��ވ�e���m��!L�n١s��e���N`^+g\�����}�Pp���:��׹��\�
�qFo �E��7�����޿��Ҩ#�N�2E�Kow���	�m	^
�g��lA��Y\�w���q��O��</
��{�7�.|Hۇ�
7"��9�׈n*A�H���){���	�䇑����j(7R�>z�z����B�{�\3���K
%����Wڼ�]jPݖc�m�X���]co�?���0��q��3�]M�pG�i�R�0'%����7�@(��4\�[�c������w��1A_�w��+��G����۬~`�rfxX@ �y��1����D3�=v|-מ��,������_�D�l�^��f#x��iGf�ث������C���΄�5��Y ��8�bA����.�f[��7S��6
D���Xl~�V�C'ݖ�9���j��y2Zg;o�&��mE����hٷ���&o�+�9�ve�*�!�'��&_��yM=>�)���z�N/���ܼ����X=]�=X���Y��/�\�����%�N�8:_��B�^�����j�%��=*������i���l`!f�倷 U�Gv�՗�By�����߭�$Qf�i_�5 ���q$o�6{�g�aR��j��.�zԨ@U�[�yiBnm���{�Q�=pX��#���(� �
�Dbj�1M���H��=_#�G�)�J��d�U�@/z�a��n?��Ģ��"�������e�,��i�o~Ѿӡ�|�k�����؂,�Y?�'�r��xhFS�tIȼ[��UΎ*�w��:N�K���`~G�V����/�$���'/;r�<��]F좹�y"i?�dRܜ�H�,^%֕�e�-:O�C�+���<<�^�����2hG��ұ�ÿ�F�gZ )ji7������*���䢵��i�h���|UX�X�9���F�g!�g��KK�\$�Z#�⠣'�7��v�;/04�xWf�Kx}ĵx�X�}��|'=�7:`��"�:���u�l�Ȝ+7��z0�-�t������n�����;�=�oR��v�+�'���2�T����kթ��|�gWJ��Q��dl;��}G�{�l`�
��yk~%z���P��Y6fE�2��=�^E˙���(.��� xِ�nؠ����g�>�Y'�hc^a���v<��B�|&�w�}��=6=H��2%%����}�.Ǝ%����_Г�d��Z%�'���5�q��@�����#O09��L��&�xC�D	��i'}���ND|)M-y"�:����>j��a�����U.#��Od�d�K�Pw?k�L�ǧ>5��sw8=�{�[�Li��v6���dI���Y�ii�{j)s����)0�f�P�E���W^]��D7������ǂ����E��j����l��'��F���X
t�T�K9��H�4�$�,8�W�^{��5�Ikx��egr���'{�!�/�M#k�>f���`� 1��J;U��}@m�:f_��6e��`�4����A�l^Mq�8��F&�*Áp/;�< qi.4�k;�*���E��10�i�~BcyW�ے S�F�ň<��qs��8�D�;ב�WM"��#�$�t�������-=�7�E�ӭm���j�!xӲ0�wJ
��N�0�ءK��2r ���څ�b�ދx�e*�>��F�;��:��<�X"B���/ <�y�^��u\Wrk����܏{�a�*Q�w�K�~�=���r�+z�����/e�7}H��.�g�`�[A^���
��e�F��� *�+�>� ���-��«Uh6���aǶ6}��HG��͏
Y�P�7j�ּ�J�}'�ؕ�O�q��=$N�:d���,u�{ߛ(�c��D��9VI�w�1)[�(3���"�>�,)c"�-�_�K	i�+G�����Arx1U�d����Hz!��5���۴��wף��˨eT�3�0֮�HI�w��;̷fci�r��Q�C���8��!�]� L�A�X�_�����V!�P-���'����z�9�0e�ڄEd@�̵J�Eu���r~s/�䐽�'�!KU�U���>>��ʎ�}%�..<��,>��������)��r�l�,�2�an'5tT�ĻǿЇ����,��4��E������"~f� �)�%+%�ޖ(;���O�ԯV��
:�/}��26��N��ɀ��.D����1^��JY���~����|�~m7\�濸ob��'f&څ-��G|'2��V7ِB��4q*�v�01��¥�V)���_2�򧺩� ���cض�`��X>����t]��w21��d;�ՖH���}:�@�
����qkD�����-�Nl@���L�����!�[9��h�����tw^Q"�Z��E,��%y������'y�S[�ܐt��Pyg8-i��&�~�mH���D��U�z�Y�Mׯ��C6?�Zj�W#�f��}=;�		<��A1yv��w�'��#��~4;�i`er����ۂ�s�Ĕ�0�6�8Q>TZ��9i��\�1]{��6�h�8La0~��M�/D��(��]c!?��$t*�Z ��gw���2����
ɚvA)�=s-�����,����'z���hx�Axw�UMִ��o�'s��%����h3��AT�	Bfy�X7���L�s�Rr����[�X@�FC�>\�"�k��J�g�� A2�J����>Q*#�w�TZ52�6��מ%���eA�=7��j:����oQ��;�;N��PF������ګCKC�򠋚ԣ�҇�� ������Z�'�OK�����c7V�X�}����L� �G���d�����F	�ZO��W#�s��˽��iF�[C�ֵۤ�i�P~�	�n{�z5�G{7ɠ���oZCK�7|��A�+��Lx�w*<j �����f�}F����B>�?=��4�<�q��U�/�e�x��C���0"(�4�iq�:3�)�c�V���@�~�����ͿLU+���o�"�f0�3�!��������5��cMJs��=D�U/$lv۪�	5�,˾�
�C������cT��Y�X��\Sa`A�9��o�fS�]���Ȃˀ�l�!fѱw�Gbn�gM������#$��t�iZ�����g�j����;mS���F��aI	����">���S(Y��g��;n��aGc'���Le\�G\��!E>�ߦ�j=#͈?����$
"�"��k&I��@dR	�	��7b�,�a�65U�h�_�Z<�f�΍ֵԈ������j�9�)�*>�Ԧ3L(���bWZY��!M"5qǠ�yy9^���ﮘm�ԅ��r�>؇f�m��j֔Y�M�:�b��ZG=G��oPS��?���:���n-,��J�G\�n�ȍ
�0���L�H�vf'�c��ܮ�0[m̱�5*a���r�[����U��#�<�[���h�^����5�BE�t��d��9���CՎ81��W��	T*�ʵ�r��&��p�}�i�{��k� h�������q+�M^����|<�:�^�TU�Q߼�-���!"F	6�΂}�作�G:%[�HU����oCr��8*{|;J�?����э������,��++(l#�PtO��֝4�U�aV�e���O��=�v娪:A�_�L|�2�j�Q���!�V��+7� q���s$	f�������?�&I�a�f�9'�)'�����t`_gU�����X؋��n)X:*#�<��L�l�- L�vPAN1$8��E.�q����HF������>�;�ĄU���=멖9�{2 h���0-g��*��B�
��չΈ���-ր)dE���u-�2ɩ�Uҩ~��@~�����T<\�v�Zz����M�����?y�/�PXʲ�@��Z��Ri�Y	�!3��_$������ks��A�u��8T&�gpک�h_݁�m3��8*[�U��?t��=峹�MM��ˈ�H��}���:�+]�N�q��o�]Q�z�`a3h�.`,^3�R�*��);���2�xܱ��Wj-gn��$ٟc�К�a�d�r��4R��7H�ZXw���l�,#
�ˌ�ԥ8 m������J��m��>�UQ.�.l������`��X��(�2����G���5LD��~TM8�*� �96٣ȁͥ9k	uʔ��rrs&ل��z� �T9��(�C�6�DQ~���3��7g��vꗮ
d��Լ������ �9`��yy+�x��5J	&h��=k���Z�KҶ�`P|9����h[qL�a����Gq]�/~H���z~Qp�&2�t&��k���N�YPsT��~����o���D!�5�R�o��D�P$��@Ѿ�Hwp_�� 	Mȣ׶Ԁ���F��n�|�_��4m�S���e4f��9L���,+Ci���8�N��e�S�k���^�ê��'��5�����r�i/��_c�
�,�'���1���������NS��z�|���� h!�(	B�z��x���v�ht�A�b�� ���@�c�ѧ$̓n7�ÊkՔE��X�¦�K�Y�\��.{�J3C|%3:�_?W���;e�曘��G������06k��g��4^���YXV�q��Z�x���D�]�y`�� њ�m5�4��\j��'G}z �Hf��ᓺsE{���9�|�Cn��P����A�O��@��z^��Y&�K7Φ[0d���W�6z�"8��W���8 8p!��dqr�);6s3�׼�qq$7h8����P#�3}`��JF���%�.G���}8�/L񨍗�G��fCT5��`[[�T"�@�l3w,���X�Ե�HV�DFs�ߔ�t��pp�C
,��'�&c�i��s��2� ����f�c���Gh�^�J��)8}�2YEɝM
k�]9��]��Q���1%cEP��
W��t9ӣ8�����f�Da��VM�>�桼}r�?��d��Pe�IF���J<}�3U� 랚�`���S�B?h
��"_Զ��,��I
�ʽ	����
�3�W��{�ց�޸�n=��̣ƃ�61�%F�PT��>`��E̑�`�k��U��5��Y@��O61�˽x绦�o��H�-��s+�at�H�$��lG1�w��r��Θ�te�Aq�Z��P��}��
��n�����n�XM�F�����;	�� �i��I���c#�`��]�l��)��d���B��x:��?��y�-���֡��ײ���!��_o�#?�8�-
 ���E��$���N*�ܵ.{�-��|\;(Ķm��(1J��i���r��s�d.�B�2���D�5��iHS���o��T�[����{�AAy��m�KlƂ"/��~��<���������R��"�_կ�3mj�Tob�"��r��:�_�2+Η�?B"�Kf���0���b�b:�1�&��7K�pѕk#抢�z�@��9�T�����;ʓ4-I٧�X�>`�>�Ȃ)E�s��w���:��o�Bp�Uw�?{��-�w�����&��!�� �� �O^H�H`)ل�3�*(ۈ����Ւ<�\�nrb$_+b6V2j�ϯ�Ω�,�ރ}��+~��m�m�\s4[�������)�N����أ�\�K�V���ʼi?h7�2	}9g�^�N<*Owgc�����%�>�����8�9L���V��6��H�n��llu�]��������뼚�4#�l�~��9�b��H��a�L����'��f��K�k�����$c�H[��+�:���B�X4F��l�V�W��;���#���_W����|hM;�we?M�E�Ǖ@����A����d�n��y�>L��-��� �3��H�4G���T�.���M�j�!>Q�DTo6V�W��|�M�U�ቇ��˦~��Ez)cm52˹$^bN�x^^��!Vۧ��R
C^��{ms��8O�g��$����\ ��cz���(l&�O�F���g����P񹏈���vA�v��B�ЁܬX�"�H��lJ��+XEdS	��9[~�a���1^�#`dg	p�A���wN�x���#:������K���5��:�/�W��5��%Y���Id9V��c�qt��Z��V�6�\�:[��9G�rgZ��W��_���_�X�w�{�����PcO�NU�,��Q�������N.H�~��x�ޔ����ZO�pTN���Q@��q ���X��gɌ�<][k2FL��c�O&�t�$^�S3�o%EKȬE >�:2\I��ԃ6V��?���_.kEP|�c/�i�"n�KV�;.���dS5O��`��H���qIX��@� _�#A锼Ds{@��p~��+�l��9Yp�������M��YTi�R;�x� Trvzʊ9� ��6l��/B��g�Lb�ץFbxa�'��Zp^�k�=�̨�h8�N,����vr���������,h��j�k>c�e���s��t�$�+� ��/5��� eDk�;�M��谽з�Ǜ�50�u��o��Y8UY�~Q4�y|w������ .4����.NwǙ���SQ<��g�t�(Gfj�c�ڼ�3�0<#}9�5,\��Ir'��RdN�iA?=کx�0T� ��g� �e��|
I��J6uO�h=�(I9�q!D�,'�M)�MDv�axQ�sJR�����P��g�1-QЀHb�B9�TL:ȴE��T��9�$�X��ek��
������܋ۘ)(e`�����\����FTG��Ȉ���\W�?un�&Q��[ӑ>~SH��MJuA�+a������s�4/+�:�8�맿�|"�ϻ�o��n��@�5�~����G�+@��+��z�Y��b�h���0��c���Ƙ�7ǃ��`����D0s�eY5�R|��D�qX��8\�P��^��[��W&�g��@O��L8g���>�閉��^�&�,'�|�^�p2�a�&�3b�����]��e�iX8_������ �i�z����ƴ/X���b��b!��,o�"�G.�S�!in��F���$�q��(1İ\�o����x��M�h$#�u��6�$�L���@pd��S+{4ߪ*�05�^��Èw���Ƒ7�s�j(�f�<�voqmu�O%��v�n~��:w3����:|}$���T*�"��[v���v����/�rv�
����^dB�g߫:Yٟ�oZ]�h�� a��I�z{�Cjf��v�G�)���"��EZ:E~�.:�nwBv׿�2��ퟣ�A8NP� ��=��yg�9�
���(O$5S�S������U�k3u���P�������D�r�@Oʟ���ۭC���&SB����>�F[\7)��s{�&��>�2y����?�����:K�RX�#���Y��I�b�C:ڏ��8�w����@�D�|�b��\>��G�3� �l����"���}\D=�
���� �|>�;��z&NRL-5c� pAiFԳ`�E��x�<
2�iV�
4��,t]���m��f(���H0B��-�8S�#�l�&xp��v����0�iN����(a�}�(�؛�u�qt�z��F�<~�{��2�_hT/s��ᮤ	���g�
2O��
8#욄�M����"��A�M�5���+�Zo�q1����&��\=�Qш3���n��O���fs�8��f�.�>�d��h~o��E(E)������lN�`v�0�`����,:��.^cL,�H��x�?�O� �ߩ,��p���.?�'�,�͚V��s�ҍ��A2@Ad�&Xo�g�-G����UWU&��� �7lQ<��&�5�q�8ͱ�Ͷ�up%�Z�f(�Cp�:��'�5;`-���J��|1�O������]�$��;�豀N����"�rdD���t�/&GIpZxuN�.�+�7V�@>�Z]r��\a���.��Ԣgkζ�[^��	��a��A���^ոO�H��M3v��84���������Y�SB{��̓��J�Pqnim��\�Y���Vsඐ!���� ��M��_�RI�W�H�E��G��U��}dpd]c\9�|�ݙm�kȩǁ����0�`�cK7��?H�Z��(�9?�ԡ*3�|1һ�9"k�w�oM�� ��*U,��=�iB��O��a�5���-����uY?�yG�c������א��d��_�����9�����#���)�i�{ ���ʚ������Hv;Ñ�E�Ej��;|4��:�U8M��[�[��Z4Y�h�h�ܣ������}����vAg����@�ꈰi��^Վ�q#s\"q�%ƫ�m-ȁ��&��}�[_��j�0��j�y4�c��M|�‹�����Gj&�Oոz�$U29
�so�|������3�aV�������Ӣ�Ԛ\i���("�b\��J�A�+^�<�u� �SE��: ��] �A��\(�D��e��ƎKy��G�j��u�J[�&�&����}���X+��p
f ��eC��e��3H�{8���5�?����lW|H�ʿ� yߴ��^��8��_�e���/"2������|�����E�7�&I��
����Zt�=��� c�J� o�nń�Vn��G^��e�3%��4x��1_��6e	D�����!]��$�J!��R�9�K��Y5:r�iql�q�-e��K`�f���DUB%X��j����Ě��M[47Zډ|L��1�NW�^1�l�~K�C`��
��c�Ҝ]��,��#��'����@��ز��.�"��jxG�-�"l���&L �m٤W5�����c�����i[j��x.�ǩ�������`:�3#��N9�6~���ݪ����8���ǹ{�B9"M%�ڝ���'V>�µ/Վ��ݞ�x�������NGV��~B�Y�\o�JPv��Ȅ���P��.~��%�. D3c���t�
�^�Ce������M鼀���q�bNZ�6�$C���xgZ����V8u�]V��˛�d�k�c9����p��G���'����������Z	(�E�t[���Α�e! �0�}E=X/��lh&<pSHb���%+,V�%����7�T�����FV�f9!�D&�d�UK�fluC���w��-g��2�<[��n]lB�A.Uͷb����=���2F�I�f��"L�%�Èy���K���X�Ͳra� ��H�2J�g*���?�@��)�#�qcim�]���zL����hH�d@�T���P:�S"Mx���J�@��ƓeU�_N���Z9g�J6�3x��W�����\:ɒa�a�B �;��aK�Y_^�'�7HG���/!������`&
4dS*���o���<����ٌ]��q�y��@n>�.�1����٧��WR-�ǕA��zS��|%QT���?���{�u_��s�1�����@ل�xQ��_��E�]�-�E���M�I��+��i��Y�C�S��8tgH�3�Rޓ�T��q�� -���>eJ^�
���:��k~
���:���"�zTR|X���é�,U�Q��f*�7K ���=A&��x�iJ��4�������\���	\А��`ؒhՑ�(]�<B?0,�/�#R��ʠ�v��4sDwoz�ؗQb'ĵ�C:��B�|=��� �(B|��cn���9��6�Ys,�3�y���#"��|��o,��FLO5�ڮ��o��-	zl�B\i]�0 865y�fd��?]�W�����~�� sHo��Z͞/p��\m����:\�}�����#�k+�6�u`1����[���!zUi;�:IS>M��E�gN�$-�~�R�^�y/h����r��حa�e]g�V�"�3��sʍ`ϳh8W)�Y���� �(��ye`#վnV��;����t/`6g����5dE��]r7Yoq���}�Py %����I�M��z!=�ӈO�"1�o�:�(dr���q��x��|���@�92I�8 ���P{�U�!ݝ���c����q���/+(�p�p�a1��]��9p爙���մ�soKl�W�[�Q��쾆T�`I2�~.�Ua�r� &	9/eR�>�,í<#`m8[��:c�=$*h�9���2�A�R]��,�D	�W"Z25����B���2���d��[�	��*��� �#���h1���32���XN����r�k�n�a��o>�:L7�W����P|���q�;�J����E�X�ľ���lk��5�E�jf;&�Rpxߎa��	R�����5��X�J�P���On�T�5��#tn#���.�J�1��kH��
	�Ӿ��6��l�a�p`^mxu��&�|�1+��^#.���j��8��Vw��ں����&�0a6��&�j�w>�桄^�^t�R���B ����m���?��n�<�����9O0��@6ANC&�'^sC�Jx���DU��x�����јe�("1�m������T��z� ��`�s���?ꉟ�j�8͍��D���6���,D�0@�<k������}t��;��'ltO F�?�������"�#�>��\l���y�9(V	w�쾽r�;��yQ�7�8�W�)��z�Wa`͛��p*EҀ'�O*'��N�W}��q�U[Irƀ�zb�>�׶jC艅�����s�r4�`Q�>TU�>��.��.���<hx�|[�n��߳38�ץk<tg�w��xصA�����Xy9TV^e�h����IX�=���fWi%�қf��u�9�����9&��L�k�@���/2-�׋(cJ����¢�"��mB�W,�q�&qb��ڞV�G��w��
� w&�c�6<�0JȐt��9��:;x�F%SQ�����|(�k�Οk|�}gz�b���6+c��' >�$'��>Ә1�W� ������
W�bmł&$�̈�o2C+�Ȱ�u�rO2��x���e�6��{�ދ�2΢�{�4�hT�».�3��Ӻ8���?���� �X� �K�=���g@�_ej���B������s9��I���b�^c�U!�����'@͔
3�Q(a�|��*�"K.ޤr��es�����)h5��Q���f��S�ޭ3AK%�&���bz\[�QU�$�n'��MX�X:19��mV41<����&�t�U��O�P��T��`�Y�Qŧ���6���rBm6$ᆜ��B8xk"�0��Z,��W,|T�7� ��a��g����ˏ��D��`k����������c�o."FeЪ�3[��@�8�mȏ��ԫ��8������נ�6h��{�a(�4�D|y�w�g���]e.x�)��� �G�]�먙����{���ī�-�b :�I�3C�����L�,���;#H��唟ʕ8h�C���:u�~�r�=�sW1s1\h�[� �����M�S�_cǲ8Ʃ�c�4H���Ri[�#|:�{纎��4Ly�c���4Ռֹ�J�b���Lɪ���d�\G����>7���$��Z��U�:1s[޷K������o�i�ח��N�I||����������5�W2�����I�8�K�N=U~_���\'LF'��(�Ex��.U�++4����m�r#��� ��t���76n�#�F��.���$`�
T;6�|P��j	g���"���*���]}�35� �	�lS�Z����M[iH7��)B��ùL׫ �'�jJ>�Dr���8e7J��� ]2.����+�P�\���I�X�v�s��a��&���7�)�~�"2��y�1�2��h �oKQ\"v G�(���߷M��|Ź~
���+e]H��&%;$�Z`Oa �K�f4#R�����3���yS�ԧ�]Bp��e��]�I�'��o���͕� Q�3���Aށ���[�4@nb�i�$*���\�JA`M]��DF	ǘp�&�E�2޷��&�\��	O	�*���xsv�<Njn9��OuP%i)�ۣF�6�����}.����ap���<#+ih�U�m�-TJ�񹇍d�V:���E���l�X�C���!����03��68�4-$�����m���5+�z��x�j~�s@I���t)4vZ�n��S
`	�K�3|HKtn����Fh� �p�������.�+{@�)�R�֔�QtN�r��BS��1�p�W!�ӊSq��.k,vΆV�o8W� D�Eq��=�a� ���ygؗ������h���e8B&��ڈ��G[3�<�T�O*��~!����-v�O,]����Zq=��LM�@h
���߷��Pagj\c��ǌ:wZ�o�"pEm�f~{�`4����(�Bcΐ�6�P�B�������Q!�2�F4�^�2�u���"n|B��ܣ0 lq�	������|w��p;SK�+��유e�|��Q=ݬ� �ɟ�OK�8�q3��)��"֛�i�!���"��&9g��!Y�Yޖ���h}��pboЋɉ��%5%�
��(��Mq���h�{�j�
t�KE�#�D��v�B�)���ϭ��x
3���g���]��M]�<�Q���uB���d9�k��:��EdQM�p�"l�-%*[�q&��<�t�$��� �8��qNcu;/#=�W��h|u�T��ܟ�wX3�7Ss���Y�:���G�4�k�����<�1�<e���қ�j���O=��j=��I����0k�����+�^�9�H�n+�3Z-��H&��`E��
c��7ߡ�1S����e����}&�$�N�F�/�I���"��1�X����e�J*u�t� ����י+�n���M��P��⠶��IH�(�.9J����m�P�og����+Z
脥(�>�r:Y�6o��������@i+SȂ�4�>�n� �)��9o�Gײ*Bu�n%���9�X>*�UlǜӮt�zw\�բU3��7�7x����L\���F�]i�����Wf����$&�.��4jY�ѯ�s�Od����zG~��͏�!�	�p��&ZR4^�?�/�G����YD�܆R�~���ۥ㒤ˈQ��2i�Cb�)�|(971��J������2��q	\$�rj�9 Q��&�߄H�H�K�>C�Ez����\�-����r���埧'�x��9����c8]�s��>�!T�o�*T]hGe�)�
�\7V��PE��+_!��vf;���'��lKQM�p^��R4��"^���,{gΓP�Z��Lu���P�?�3�1�Sϼ�(����%�ɢ;kM���؝�i@��x� cz:���z��P��B�b��2��pt�ߊ딟F2���
��:̺
��	֜��u�T����'�$�4Y����`����=i9�(#->�+[�&����Z��N<���@-.��Q}c�}��oj_I����Zg�\��E�$��`�3�5��������l^�fwՖ�T��1�%.�\>ڭ�S$��
O"J�0�U8�]��ު!(���R3Hy�Q��;��b�5��3�Q5q�M�4���9�{�Z�Y���5A���|�U��7�쨶8W�w5�ፘxR3m��0Rh�����ۨ�dFW*-�J�\��
�r��-h�D�@	Wj2�њ��I����93���:��H�Z۫|"�w�A�u9�A}���71^��t��]�����Ӥi�$���젬����̌�j�B�ӇQ����5�s��^���*�о®Q:W-�ѓy���X��ٷ�gKk��i_�1,%��;�v�A��Ujj�)z���&*���(7d�6��ߡϷ���Y-�jG%&*ܥ2x2Z$&mY���oHl5��i�s,șc��1��1�T6�h��8���cKz�� ���cQ��B��k��p����5H�.�/vT�Zۼ���y`n��ҹC��K;�L��sH<H&]��0��.+�o� įR��,є18��Je��/��B��l��r"3),wjڿi?�:��u��NF�v~s �)��	�IplH�;y4������9#� ���LK�� ��Җ%a��Gxl[s��� �h��f�Y̲9U�N6?��L���[���C+���x՞Qy�,��y��7WH
��3��k��Z׺[��h+\W>_:n���J~���6����
���źQ�+0l�یV'����pܻ-�O��},v}�P�h�ҵ�V����W���W��$�JU"�������hZ�[�bQ'��)g�v0ArZ��R�j����>%��fbQ�7i��'C��X�GE�� B
���ϭ��Iɱ�.MQi�|��-�5Stq�(*l�$�0޷��\�y�vnjnb5F�@jӲv�鷷	\�2��U�N�R�k=8��#G+ӱ���trB)e���Q:u�o�B�c�c�>*��⋑7�贒�����(���Ō�]B����p�]Z-�o��.Pߦ�|���م{V���2�z	��ۊh�A�m��)��av��'�������:� �/�.��n��q;�S��~"/�?�^�l'�������	Q<��Z����PZ��d�+��WɐjE�$@�ͨUI�hx��iBs�
�Ǝ�v)��;Ö�5w�mY�����
��_�x�3Y�k&�wj�ǌ�p�����b;t҂��� �"�!c襊�&�f�L�h9̚X}n���x�p�A���]m�Q���0�� ;ƹ�`��kLZ>���n����"ƺ6�E��g(U��
� l}���u��E]��;'υqꡕ5�)�:
�:Jdz�t�I<U���kg��8e�����y�,h;_#��a����O�<A��|i ��7����Xr%�`�\��q��ܮ��r����}�Љ�%
�%p���<��V��AbQ�LH�}�A4E(J�,�M�������n�'���4UsG�,��KSaؕy�xɿ����,�YЌ���kHG�x��ќx�֑+"�f���}!����sB����vf"�����2L�W��MO���H�O���M>H�ѽUr�٪I��$�U�!���W�+B�)��r�\:Ę>y����w�#._���Ӂ ���m�^�9m�J��}���J;8;�)u�L��ꂪ]8C��4���캵��ISE����K�}��7�� B`��7�T��� �$�1%�����B���b�dX�1�8��o43��?+fq�4�=��;�:W4=c��h'C��̏gf����]���+��y-a I��_�iu|^#RTh8��������$,0?�|�(�W���%��?q�q����ā�gZ[@!��z[u���6�N��h�МqB��o�9��ʗ:Z�:�1����|�-;�L��I����&l�l�m�idx��$�������.�<�y&�A_i�ۄ)��(e�?];��N|}{�}`M �,���6�pn�A%AHwٌ��W��~�tY����dj��;?��?bT�@B%��`.�:~���R}V����]S �k�}�͌:f���uB[vA��t=��J��[���[^6��2a
\��$�UAhC���(�N�댿L�)���s�~�M�`�w�T5�A�����R.�^�5a��1����)I�X��� "I㵓�yPx�#������bT��.t�?�����I�Y�9��]C�w����Qd��������}�tV�a�B�͉�HA���I2��@������݈K���#R�T�;(��w)��D\��rZSE�}WD�f$�s�L�<7y�  Ԇ�&�i�m_s����s��]yS�5pݖJg^�G�YB�'���|,ke@��'�z��~��[M�eDQ���4�2 �`ϿgC��40�UF�/r�-$����-��,�r��������^��umd/��&X1��X�#�:Jo"p@X?B(w}!�jv^�菜x�4|��;�r �8�$V���dlY�4V��`(��,�M�$L��N_D�x���F������R��8�P�"/Dp�{2Hap�e���E�I����cֽ�=P�1R��N��:�v�*O�S{��5�)�6߉�~��[�C����U����A��h6�P�P�ƧH�~��C�C��0.os��[r��?�3��C��P��ë�-��DFEF���3�L)+�:�rѮq�D�d�(�*|i:��P,=���)�<�������Gc�˭�sZ�2K�%t��	,>�ut�M"X<E0^ ����[�xm���֠�|@<�S�CPj�g0P���^�T)+�En���)3j�t�����a/���z�k��s���E_��m�m�7�.���¥�T��Ҕ���O�a�]���(������2�A��)���;��ċ [���M���n�֪������1�O_'�Մ'�h����fVמ���c��tP���j��U����[]���g3�D��ٌW������A@�\ l�l�� �D��1F��\_�_
`������M��\��P���J���Щ=3���;
�೴���]H"����CbB��K@� �������ɼ(K�-BG��xN��̵D���c�:�F}�z��+��w�;��R�'�2���a��A���2����+��PhTqvO��i�sd�YiO����|�K�N�66�i�3z�}�Q���<,��A��r�k 9F��[i(+�t�2R55���Ԕ����Ӏ�e{!$ϧsW�p��iR/Ei�.'�a��k+M$�p61k�٫	�*��SgbP�g�	&IH�ϓq2�t�z`A��'�۴5rOv� \QՖv�ٲRf���ɞ��H~˽F�8�xT�g���Q�+R�l%���+�6q��lu�{�`������\���_�:7݋���1��
�G&v�a��р7��ׂ{w��Ʒ�c�L��sU�:u(ғ�|���[$�>�q��	CQ1`TB}3��阾b}�(��cB� iʸ�if T��%"���z�����!A������hfﻵ�x.���;�v�TQ:=:X��b;��_��p�1�2�<Z[���[��5!�B��2��$9>��#yJWs�#D)Mߡ�� ���jHf�ӟ]O%Ք?�_
f�C9]=T^T��QG~�;��g�ڻ�iF�91
�dy�+������n#N��&9�̿i���CQl��+V���.��1�|�#�8z��G��F_a��Q&bג�>�9��օ@�_���waKSUA7��n%����4$������G3*�G�/�?{��q�#�O��
Y� *�eW�w8Y��F83V�������R���8%�ʭ��+H�x�s��t���뤠&�1s �bՑԥ�3����F��)����ƿ0��na��j���5ޭ��qс�7��I[ƓJqV��P98�{�spe�ܚ�s�p,��Hay�(K5WG��:��8o����zG�<��2�&�h�}[b��e%�K6��嚐 ��9A4�4�l�L�E|��i.�����jB���M���x!���Q��(y��zC/ ��滂��R��bB8��d�-��Nӹ?X���|�R��
Q�7�����:��f��~8�7�N�2���.G79�9��1�U� ��Q�7�2�<��oN����T�i� ��i�r�k&fR^�D6z{�)p�T���k��߹�j��e� cr�"q��*��EV��=�b5,�[w�~xnh|ӿr�T����yf�ǰ=�ݟ�;)��kf��N�I��,b{.�.��q�J�9�H��K-3��Es�p�P��j\Y^��	�Z�V'Б�[����;�T��#`�"�aWm� ��t�u;f�h*D����o�ͣ�.��׼إ[0�N����U�/�Lg8�i���!oto�����E��ܭ�q�����٠!?����a�+��[��6��RT�u�ma�x�Y�������;+w��U&����-5�G	�{Hhn�i�B�H��@����2%1C�	V̠_W�jY�h�����OY ����� #?�kmhc�b+)D��\���Z��fZ��<��M .��*��@�!��DN$1_6v�M2_|�s��ʪ�_b����ʡ-�,�t��*�Z��vo��{��d��)�J�D�z ��>��J#WԱ�Z؟7�f�%ty����_�������A!2�����@��5�W��l\[�0��*Sf��5����^�qO��H��G/	+�a�G4k���c�"�q��p�'Y��(	MWX��p��9F^�ݩu��c��]�N uI<t�F�8��W��k��-��w4k��KjS2��гv����Z��2�s��Y�U-�7�Su�����k�}n�!KH/ћ����E/]�Q5h�3�h��l�怡��=�e|�G>����G�0�,|��'�I�� Y�ͫ�] �}��s�T'�^�
���q����I�[4�^A����
"=H�[�]q���eȡ����~y1*���K�W��Zg����K�b����0�s��N�&���`�Ny~���߉�d7c`^~ss,l�I� y�P,}�ϰ��H񡳒 �q���b�\US���ܜ��ÿ"�wL'֬��K�+�Yx�/��ȩ�`G�=up>2Ӯ4��)㵱ϲs��>l�>�y��ٔ`��T�"�ߒ����Ul��X�I
J*�"�˝I�=����D��b#z~|帨3
؏��0 �ǔ��B@���C٨�(S-�/-o��p��������c�h׳4��{��\w��v�no�	k�>T���� n�ǂ;���� �dZ
���!�?��"z�Z^�F�h�Va�JgU�}*��Z��C`2�&L��畃A���}U���Ŋ�.C"��Ĥ^�Q�@���~�yM7xT��ɹ�r�{��\g��#E"a����� #�Z/��t�����f�Z�*����Y~CNg��}��R;i(��pDZ.�9�9��p;��}������J5�u�'�.m=!R�>_%$J�D�X�������
/���R�9����7�1�|�s�-1�e���ɳ��R*�h��9U5ﺍ�0%��!��5�4�oP�d&����~�������̓cp�1?�����Ƞ;� ������7�0����s�2bM`��
�qj}�q8q�����^9����-��p
Y�TC�%pY�x��X��3�ae��b�V'��Z���R��t�@^�kŢ��uc�ێO����}zu�IȘ��������瘒���&&�(Y��SO�)}j�f�b����Z��i��A�&��HK��ZҾ���9���_1`��
x�bT#Z�M����B�/�c�����ht���'��t�m�o��Ґ.�?l�s���W.����e,���_A��a��Ce���j�\��w�Y*����%� �3"�M{w^��%��E�~��aUQ�.w�y�ذ#h���h��%��]�hD�o�o�@Hi/�@3*3��c���E���<C�D��a���`2ʝ������ah�Y�څʴ1GS��C���ߡ�!ŵ�Q4���p�_@�By�~d�{.���C��Hҭp�c�8�� [�c|���d�o��wC�O�ǁZ��9�"����̨�7�ZZ�C�������2>�o����2�ݑ�r�9q���+#����k7o�s��n^�=}F�j�%Hk�%�6e�$����@�^�+�S��z{o��ׁ�Pbd@��Դ���X�Pİ�ᐐI`]�uX�lm6mg��_ǟQ髐L�c�8�j��oĴ �0�u��t�OLL����3�|�μ�B�.\��>?ณ��`{I����g�� 1п�lMZ٤����b��{�c���z>Dj�b�T�L�}���d�V�H�+��ם�;�M`���虸b6��|ɱ0-?�Ň�����|׵̱%Ե��B�3��ۆ����8�S��3HRj��#�7��Ԯ�O���A�aTԤѓ���P.I'4�Ue���?�K��h���"��X[vU���Ъ�n0���_'m�� B�\H,[\����W���GT�V��\�qI��ClJOf&PdG�ʆ�Dw���`Y(n�C�ǔ��ضȮX�څ���)45��\
��`w5�������@FXMT����(�Q����8�;�\Q�K��ofY/rwF�X�{�	˴`H���Uޓ9�:�w��zK��:�S]*�� �U������Z���H@h�ʡv�g�X�r�F�fo����^<&0bz�!�
J�c5^�����G�Z�}EL����*��/'�|3�:���3��{^�(��Sdr�4�.��A���γ�ڗ<����s/��4��i�1']:����!�#�E��o"L���p�v�Z~L����U��&zt��������y�/v�p�~ C0M<��9����YG� pr�����}�#_�+�Qҁ�wfՠ }�sޤ�&��w�#`�upO�J���5(@���0C����Y�{���84�]��i�u���8y��7��i΄��U�&sZ�xV�V�!������zy��q�H�����j�>��E�ؕ�t�5w]�ɸ��濪�r�/b<��E�"E{cVް���P�@�"�����']����k[қJt�ey� �D��7�������Q�n�ͮ���V/o����Q-�r��.5Ӝ�<\m�0�l���U��P
D�*��=&��{��=֗�8Ǆ���i�^yn,���i6[w�;G����&��{Z��i�rn&# W(O&�M:�J����U�}�U�(�����Q��:��MH���:��3����Y*���&J�� L����ꂭ"w�8Ȯ����e��=F^*_�;d��pNۑ���Я��i��I9�'4��?����8���k�f���-n�@	�Y��R�l}&�)̍���0���$���m\���A��1�����!C�Q|��j|GL�4IiA8C��v�;q���x*����2�w�N$��+r�xP|ox�*}�����;���ÊCF���S#O]W��z�7q�;��?���~دj���B<����箪E��}Ulѣ��f�1���恌lF�9����T��sHm���*���R���I�IzO��u��zLt��5IHh1l��DD)����D��&�K�o�sWy�0�V��l��ߙ�.C}/�.���>�9���hj�Ÿ�Cw���S���oع��	�(�{!S����ج_
_�0��&��E�G�
�>�"R^M��AUvPd�n(x�w��V�$흿����6f��2��5��!VhB��K*�Eq:?����b�k�dO�kg�s������6a��.Uz�r�ã�{f�� �:��t�1�bxfoV V�28�ŨĽO)��aR���O�ROS��?x�O�~�L������p��ww���Eh���w��5ϮFM1.�X��JA��[ �L-�>�C���_d���|����\\�ŷ�cyⷋ�`c"KU�������5�~*�@� �>ĲـM�}��kV�0�niC���6�'�bb��p�X-*�9aL&��k7�|V��1��噰ɤ>v~��V/�\&1�9'���k���S���'2ȁ"FL6��c�:O��ܰ\ڇ�3��l>�Zp�)9��*�7��n�c�