��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;����`���仢���0ɎrRV��c)`ڔ
G]����|�T�z
ly��Q�@%��qy&�>�!�\��d�1�±e��
��B�'P��h����ͻ��SZ'-��V�l�5ݱ�3F=�����i�Q��F ;�}�7֣�kB.|�a\?��,�6�񄽑�(�ЗX$���#*��-B�b�D��)$�W\�X���ck�9/g1|OV�oDz��������1�9״��Ho��G1ѱ5⫄'J7{���N�jh�n�BG��C���ʢ���W<�\����笫4Ez=�2�:
������y�5�qb�׋�N]%Y�9�%qNgO7�\F�ۈ
��`�ZZ�@`(ai( ����H�A
&
S%A@�<�];˟���5�q���W�D�+�ܺS��ci�WO5i6L���>�ʐڶtTU�$f��ߢ�T���n~;�(H���=1V&]܉x�Ǡ;�l�?jL�ayR��Ώ�^=���!hi��IF��Vi��ST�3�N�G�̾�y7��iQ�,�Cp�Ȧi�A.���W84q�-+��<�I�J�}07�])�y���=́�{�bɠ�q ٤�A��;��~A_z63�ߣ���0e����\s�z=@$�;׊�圦���;�����oS��R6�u,�'�+���9�`0�ȯ%u@�pB�/��ؙS`�~�a�H߸@O�o��z����j��E���S;eh�%.�1m3U��Y;2�?0���bh����+�G1��Sh�	6N�1��:�
�:ڇ�k��äs�sni���a��i�F֑�B#M��Md=C�3X���['
{ڳ!9)�@��ܓ���y礕6L韶��/"{���
���GY��R&���`�V�"��ʏ�oi/ψ��3"1T���Ju�#��f���3���~kO]X�����y���{y�1�BI�IW��2�t�]*�8o7�5G��ۆ������*<��U�r,hf�>qk`u5����x�x�U���s�S ���������j8�����w�"6r�/+����s�p����uG��%����-��w?�~��Sük�Q*�[����LU?�t͔�����¬SW��Η�݀�����@:���s~��C��ʗӑ���X	@GP"",�#@��- ��W��v"Aj��_��1���,�I�I3񛳢_�]4�֜��s�����V��8�g�:�nj�x�;�|��F�D���PյuZV�y���R���-2oXO����F@�:+'�� �A�)�]W��1�2�$�0���s�R���+�'�%w8���.����:0� �>+�\��i�/dQ�  �3�._tD>�j����ɐK������c�������?	�N���\����-��w��]#-��<=5�~����[���F�����q�~���~��3�㳘�P�ܓ�祥L?�2�e���p(�.�L���w���6�s��ˊe}'������s�z̰���*D�������+�DkÓ��
��yˢ*��ol	�\�0�$�8J��HM����F��$mjX=(nb����	ҩ6��c���R��r��x|������Q0#�5��z��^��G��ޟ����妀WȢ�zS+�m�e�w��6:���G��Vح1k	WR�U���<�$�Y�/�����OL�?!�3���qϊ;	M#��%!px���PS@�V�����s�}.��u����;�YnR�ӊZ�����!A��$���[S��I�}�Fފ����n5*j��%��81Tf%T��hψ�������$&sU�l���(9�4<������ԈLA���6�p ��\PE~0(�j\q�P<4��fã_�KAfi���qת%�Т�,Ʌ+P�1�;1��i*���/����ڂw��*]�O�u��i,M��x���4V�����7�)ĹpS��l�����/�w%I3�y�ӫ + D��u3��5�6ۢg�/R��s�<J^!f>�z*՘H�8�E�C(��|�R��SMM8�6|{=�}{Aq��(Y҄<%��#�}Wh���X"�rw��f�M��Mg{H:<I�~����B����%���~.ZP�v�P�E�lz�QGsl=���ɝ�wMaOh�T���'�rV�#]��]���s��\W�|�F��K7ݙS��NA����y2�{�fJX��b�&�Y���lM�fO����?�euS�b�܍	���E܌�d��L��4��_8TL�J�~Ů���>��� ��m�rXn���1��AN����ȑ�Q�Ѭ�?Fbss��[D�wq� m᩸er�ᜦJc�}Ϸ$~�		Ga��x_ĵ1�FV��ѰB���i�ů,۹�ÃJܦ,�DL	�r�2�FN̍��'%�lw�9Qf��5�k|�sy�@Rz��K*_���ja�Q�|����/�}�<T�;�Jl��Sta�kv4-]@�!��C��~�+�a���l]�c^�қ��uX���a�J�tW?���C�;U���?R�L`���^��VHȘ��7�aO�� �{�ao=\~�58�j@^-Jjxz�"��O�_�"T��.�Xm�$���\}4���7��?K�.�Zb�J�1t�Q|����k�7�7X����{����>�3�G�,t!�7
��c����hw��r��Qll�]
u~m#�̙HDhS��*fK ��DrrzP�:W��������Î1����ie1¤ʿ^U��_�Ғ�Elqn�-�Һ7d`����t�M}f+���a��$ȉ��B��F�'Ў0L.����E5ل
6\��q�J7�SoDM]U-.O(��!��:ǡ
酂���Z�P�M���j�S "F�۝��2u�`$�ej ���`��S�����YB��`���z5�bj$��e��`�/��6_p�d�m�?7w<��q���ٔ����]�8<I9�B�u&�9���hP4�)�3.�u�$t��E7b��1r1������\����oÖ)T}_���gm�~��c'I_�Q��9��w�{�R�]h(����I�rI�`�󖝷�ɟB�cp�y�)�����y_I���K,
s"T��,�ǣp�!��8��fNۂ�_8���`tOV�-���P�|?�e�CB�Mք����K���yp����ϻKSQx�,�f��t�fQ�l��]E%������ar,���"A	��*F�������	$���H/3�Μ.W5c�6s@� ���K��f��j��@h+k���w7�o)��|�����n66f�h^ل��'gܛ��`,}��x`�5PQ�N��/4.����x��3P}��4�Wa�T1)�-e4�ݲ#�6��M��í�:=��gUa+d���R��}ѾZ�W�q(OD����څ��wc�W����\��F(�`J��('	��������^S���?�'/�����c�� �e"���b*�S�,������Y��7����K����c�� R�{sRrPc�q�;���s3g���5�q�>4���_�+�n�OCV�v9
a��h�8�?2�iU��>4���G�~"s�����4V1��r�h�"<���B���ݦ��0p���l�����y�|ed�޾��$0�dCK��ɢ����ކj���Md3��{)��t�^�>pG�겤��T�PH�2�E\����RY�v}������-�ȣ-S�U�2V�zf$�O	��:�z4� �� ��l��-�@�P�f�㛡��~Db2̲���p�e�ϺQ��)W�&�`��3P,���������.]��X�#�<�(W3���g��zz��`���ׄVŸa0c�Ofth_}r��.�G{�/�ᨏ�B'�I��尻?��p���׋̂�K�h��1�3T��0
�=��β���A�F��gF�N����{g68�d�	�v<h�w�ֿ>9�
�NH6B��e���a�aT��SR0;�_��¢螑�'�������݆�ëC����ʻ����C��,!�a��;�f�ύA��֙b��Bx�>u�hR�67�b|窢� x;�����t�cz���{�q�n	�O�@�'ُ�������j&pJ�
	$D���.�g���S�3I{��:S;q��K�Q,m[�]#��U\vu�G)d?k7�Gyķ�G�@5�YT���0澺W%��Z��T��c:�qaSlxL1DC&0��3�9���Y�;�)P�+.0�e��1� T��o���
eo"�.�x�HK�Ѐ�n�Vó�76�oz��1�?ɒ�%/�z���D�����3L��4*��N��f��j�Z��:��&32�U���,|6p�C��W||��iˢ����cBӶ,,��8j��IY.n�fCkU-��pH'��`�q�Z
g���8����jd�$��4����NA#U������*>�����f��c	������F�L����橜�S��7���I�99�� �6���i"s��\�Ẉ�W���������c�n��p