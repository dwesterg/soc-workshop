��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\��?�ONy.r��h��Y)�?��v��5��4���GAXab�8?�tYj  yV�v�D�#�M�p|�E{� T"r47���PŨ���������v��6����^^�q ��$�n�Au�(��2�,A���l���ь����o���3_�.*���<c'�a�lX�tÂ(�>Y�jy��y���KEc67��`sME����g��Er�H3٩+�vꌫimJ�n)�̕T�onܢ�S��5�I���6����;��V�_5Sk}T 1~���I��+�{O��2�!�$�� }�G���B �V[����E��g�[�mEX˶��Bx���h4�e����'�?�����&t�w�bpS�d>�7���B���M�l8��J������%:W�
 �O��F6{8f+��dUQ��R�\��.�s4 ��7��B?�4z��^=g���e�#��a���,s���*_v�ns,��p筴uŽ)z��#˛�'$T���<�P�ł�Z�ةc9�.O��[��(�x���sx�H�4`rS����{V}Թ�>��|Q��Xp��3��+��EƗC���������vt�#�j�;H�J����Q�@��]��0�^�Z�y���~�
oW&�~�v-2��I Y�2t�=�,q+.�K�;��ݍ-��v��{��=d����h����7��G��u�+;��X�w�#~<b����׵��Bjq�[�X�VO����4xp4�#�5��JD_ 6ݺ�ℰ��˓vC�4GFpLjP�1�����+�{����@���-](<i�5J�#T�~�P/�����6�G,FHu��)`4��%�;2Ǫ�v��Y���W�'������>��|V!z����W�M]��n�Z�ZF��>H�zxf�r���pF�i���l����CX����M����[ܭ�:���繢x[�2�[?��yu�DI�Sn��Vt�R��Tcx��iyA�'�r�Wr�G�oL�b7���B҆�3��-�_l�+�ɫ���92�lyܨ�+?P�����o�����e��Q߂�	k�$!~�x୮�B�`���|�d9.����+w��ظy�/rmFt�"�ι��IN1(�	�l����� D<>+F#2J�����p
>�9�ڜ�����#-��3Y_
%D��SS#���HpΤ��@�J��֏��i��GZN _#�x�h6�ay���:�)�����t����|-�UN�Z[
�i��\΅z�N��ޣ0�����*Ţ����z��� 9&��"�+��_���S������� a\�V�w�|�.\]}�}5�R��U�������=N٠�"��ޜ�~��ߋ�<����h�6&/��<3���elɏn�#t�oF���3�d����]P��{��u�L�/3�~�3A����|��[,
S:6s>�1uw�c�h��$��_O��I������~ĳ����ٍxdی�ͤ[�.B6l�o[m_��3~�⤲��OW�Ѓ����'I�7Qw^2��}�kf��ɍ�F0�l+R^9�1���f�}MQ?���a/�ӕ%��ř���
��L���}���X{��o����2a��ccڹyu�ut'­xy�u��qQ9f	�Q�q���e���b}�u&��S�s�[d�E����F��qd��l {Ç��'w��Iei��52z���9}$~0��L��%焏����zU	8�0�wV��'NS�� ��G�ws�e@�����l���y{^u��i�����	+����JN4֔�r��d�Nؾ�s!���g�
)��0Hum���
*&�R���0~L�ze�i����O$��#�m�v4� �)�Kz.ԜxŻ$G�ݞ�Xps����NRB\�{4�NTlZ>9���Z���q�f���X4�q���V@��:5�cce̠�/��c��C�4O;)g*
ζ��гC�%9����������UI���N��2A�D]Ebar�>
�>me��]�8�p���1\Z�#<7��>f��PoQl�^������K�v�b�=w��@���Der�zne`��5���Z'2���;�(-O�3Rz[��E��=@��<�)�����n|v��J��9�,�!���k�L~ȥ��~qXb��~K�q�♑��N���]�넶�[?p��zA��iJ'�^����L��Щ����5>-h;�H�P��SZi	�ϊ6��;��Q~	Ev�l��}�;j�K�Σ9-����Lm�/�o�CrJ�����
�����ú2�m^c�LK�k� 4V���%�]�[��c�CΛ3s�*�w�>5F
�-3��)�
>p�H���?[����#~I`�-UC�`�q�Βd��Z�����!,Q�[�썱���Ch�m�Gc@o-―��A�%�դ�?�X����	 ���c�+w�j�?;-1�fSBs�������@p}� 5՘�Cp�,����;���w�c�e�C�A�%��]�(_$U�?�-L!�0(��������1���d�
z�d���~l���?�Z~��k��4�9�eqp���b��s2�m["
'}̤�ص�T8�H�
U�⍝K}�Uy���l�W�� H�Q����h�����Q;`��)}3������{�R��S&�Yi��Ď���m
>�@�Gѥ�:�d�H&��䚩f&���|ebx&`�/Z�6�9�+��N�7��oSWqi�~~�� ���@fU��a�`�=�4�rd��@d��<L`^T ������j���3�C�{�!)L�y���������7��
S4o��w��u1؏������b&\ ���"��a�p�P� 8.`&��C���7/Ph�Y$pY�	[|%�-Y��F�|s@��^�@�L�������sg��Z1*�����QY�yҷ��'���斡� ���b�WiZ�G��ҭ��˾O��/Y�7e�[ k���)�~�Å�R�@��V�~��q1�~�Z1%D?c��V7�[Z
�>4�{ �6� L�sH��]si�� J�k��EcZ�>`K�Z�*Z�$����C��,+��w)z0�������Ͱ�Nn�܌�S;�� �����c�~�햆n�q�>M0t�ז���6+����|l�p�:����c>kRCvaw�q�\S������p�Σ������ M��Xu3���n��`	6U#��N3�0x�a����Q�n�����\�"�e,K�z�oFJ�
��Y.��.�z����������)'t�P�tn��WϠ��?�� �����-hc,�_��`�	�(���K�."�	޺��0g`j ��~hK{!��t�7��������H��5s���~\9O�5�V ��
�j$SZ�\��rX�����{M�E��yA��.����ڪ��1`0��QL� � ݩS;3���_-r��F"b��<I��<��r��>��e1aL���$����K��2��re��o�&<�[P`�I����z������rw2��Yu��>������؁x$��E���k��%����6B���8"�)��6�k�����L��ݛr6�7!�Kg����o8Яe'�]��k(���z������Ia�!gs�gB�xb��Y=�*=�MOM�.�}?G�;�?��L�����`�~���6B�?m���V���'
� `PW�nn����]U]1�8�=��
�9��5�A�GZ�		=R�rnv;fc�LD��C%j�ЯV!|�-�b �N�7���8q��xd�����%��c���F��ө� j>t[������߯�tI[F�lo�� h���7����%^�r�^);�^O���'И#�1U�I�r�SO#z�&F���ř��,��|!�>p��1���5A٧�H�,�������+!�ah�¼~��2���A�|~D�|��M����n�������FUu1H2+��!}�%��m�T{T��l����P�۵��hk��j�S�"�]u�D.�8�2����5i"W6Ur���r% =��<½m�q�>�ǔ��{�O�7�V��\�3���0�M���Qy�ʎaa�����g�:��n�����"������CuS������e@���#�o;�j�X��Ϩ�/�J���������܈�������.���֐�US
p��9�/O;��8h_�����S���HK�f��h�I�s��:��uAO�*yg�5=,�
w˓ѳQH۔ >�'R�`�0��+\O&�C�㺑5�V�]�		'��9(Gٸ[���8Azs��-�`_;������pͱ�$AŢ�����D*��O���0d}l�,0 �d����X��udU:}S������T��E�{ۚ�8X C_l��'�Y��5��г���{q��h�rS�Y���'�&
�9u��f���ݿgϚt�
��շ�Ƴ��-�l���99����2j}XvT!m�[��y'D�K#v�[ʅ=!�G����N����������I�`_�D�!����[�ރ�i��S
��84J��
8�Y�a�P�оZ��POjȄ&��%�p��F��]w�J|1�%�-F����"����,|������9ݼx��!v����UG|܈ M�,UҲ;]���ҁ�f"�i7nيU�C����{��U���O�]W�$[�}��P�k� ��Sme��4D֎܈��5���'_��_���zQ�o��G�|7�.�h��"x{#��)-���D��K����n� C�]�lYy>�|6ʲ�"��F�W��4߫\�,?����E�jŬ�s݄�D�ٷ����TOeFXee.����Y��v���O�e��/g����}=�)��:-��p�4-�2� �������h��&K`+&�y�
p�U?8��;߇P9�۾x0�
�]�Ʈ�u,����JU��%G&֩b�?�0�l�F���a5Et�u�Kq2T8�@������:O��� ����_�uh�Af��@����5�����c���������J��f�B�Rٟ��(Cg����Fh�YS:��BK2��[7O�Q��]�>�#�r%8I��Sj#B;����� �)t�Wa"�n�c�?�{M���gg�ɨJ��y΅u_?��+�L��#�o�Xr?��]��fQ��
r|��(/���&z_6��l�a
���K�ģ�jB�9��)��l��R`qOJ���^�k�К4p��� ���"���4l����c~��P]���z�cGQW���M�;�t8|����qS��n	�B�9��r��Wץ�*JL4L��JP���~�T%Јڶ����X�/��g	U����v=B�5���L�Yr�ڨ�4�E��-�X��;t�ƫ�K�$��ᮡ�u%���8 OQ6���HpZE2�'��� rK���4a����QB�^<��1�=�}��݄kK&�ۥ�o[j��+QS��e�Q�Aɠi#��q������k9��}�V�q44���l�B���DZ��6�|��%W����Who�cHsB���C�ӴW�����z���3�bl:sZ�<GO`�ϳ�Q�Jo�iv0{
��A#��Ƣ/�C2���']��� /���az�������7�%����?��H�������H	�f�).�5�8��Bz;{~u>_sY�&@�p�-e?��W2���Zwn8��/�oSy��������DJ-���$��������E�f�`[PK.;�v��|�ìq���~/\�B簿z��鄽�a��1J%�
r��[����H��-X�@�s�)����.�H~��&Vr��/3�'��I`W�o��u�@�z��q��]�Z&w5H�y�S�kl��w%���J��"	�Yو�`��o:7��\3g��;�N�zN$tr��
���,y������<�j�3$La�\�"�+�@=|0��n�GЕO�< �>���!:�_hg������	T<�+��+L�섇D�N�u��^�e�MEN�"k�{��\S_�<C�j�lk���N�u���	Z}#iT!�,U�R3g�$�UE�K��K>D�o���e�d��4�ق��]Dv�|�/�P�y�t��3�������7�x�,�9��`�����BY��ʖ+k�*��0[(���;H�;�>�@T�	4�n�,�,(�(e��,��g{��9�b>w�ξ�؅�s_�Z&�`A[1Ze^.x!ϋ�ɠC���5��\bXƪ�V����CVM�f���U�@T�#v�Bq��m?�|�,L,�\��O!�s]���i�X�xA]���f(�@1��KB5LR%.�s���Ä�F�wu���ք����˴�-�^��ˬe-�m���¦�q:�"�,���8��|���,��h2��!�-�1RB)�]���Bl��Xz=�������� �?�pKǩ՟�ɕ�������p=h`*�|���ֱ3��*�����a7I��f+�kE�6���-�aK)\��-����	�ʦ)�Y�O�p�N��3�dJ�Aj���j���63���攱Dɥv&���>1<Ln���_p��~�G�Z~��8P��3�"���1̰π�𽑻$�&B����ndhX���)��;F��]��]',gY�g%:��Ya�:2V�����I�����-�A�]�/�=�����Fq��4[�f��0���y�\�}7�;ZOq&����a}���&S�E[�ًD������gUR���$ڄ_�]�B���_�v�E�B<a���3�������
�����7e����[��K3@��X��s1qǐ&��UB�~z��i�]�nT<@י���9{��<�w�/v] C�&�Gg�(��烠�E�ֽ�!��lBd����S"@Ј�9-A�?�JH�k�NLe�6��W��0,���6мN�n�L��a�Ӄ���~|%M��*K�G6�����������䟜&���8 '�������VU�g\�a�OD���;3������p�80	Խ$puy���]i}�@$ej����Z��]ŹL(�?�q�&�Bǳm(z���7)���]��	0�vW7R�ѿr�i���^��D0��y���-p��:�_��7�/��pܲ�a9|`\���,�9{G�T���{��ﱫ,�Ϲb��~�?�ʶm� mmȓ�	�����.�0/WＡ�����+~�D״e[e��Q��>����ܚ`�⥭�3��O�gI#�9�CC��;KU /M*�6��*\	d��I�͞VY߹3��c>3�u )��'c^��>\�^�2��Pq�"c}�uG���xnQg��F�O +����Wz�s
]>��v�a�^!�0�t��٢6wE2KTx�zΐ���F�o��6#n��]�J��d��-T�_�̊M��e	�3�M�\����FQ��2s�U�>GA�Eu~�o��`ո3-)�5zB���_r�k��`R{���rbMw���gɢ3&�r7�B�!b���r-�H��l���re[��aeB����%֚o�&�a���/����'ׄ��9	@:�moob��2o�6��砏�V��*$C�
Gf�*�?�tK4���{��o9s�:�g�Dt޽�Be7���e;�E���F�(�熬� ����*�P��ݯL�|������-t���գ�����Oc��Ⱦ�x��y�p��F�QT�;#�ɫҟ�>r��2��.�4t��W��,�N�Dۉ��%���w�z���+S���&�4��=�O4�T_����Sl,nz%6
���ɋ�/W*ݔ�^�~)��-h;��������.�����#����QD�P�� T�js՜>7�,~I���2_�}���z�ߡ�A��-��-n��v��Ζ|\�Zfuy}��� j����^�'=[�V>���^\Bw6��1L�R�HV�o$A������@s����^�M�;3�v��.ס��b)�t���[T�=|�!��H�߿c������"0o���u&A9�=sp���ZzX*bS3��ݞ��&���*8�^:b�)#m��6G��A�X� ��]���qܵ�gE��	d+��3]��4�(����g�Z��n�P�/e+�OE��	�in� T�9��N�Y:c���FX�����"<��������xT�}���,����?�� �;D������� ���PU�3U|uB>���JI*YxC�q/n� �C�.�&'�t����_�R`�|��(�)(Qx=T�Y����ٞ����$��c��b�j+���:��
J椷����;��~��x-����a�9��U��N�߱��1�t��� _�J��)6�Xp��%�R����p�F���F|��o�_ 6�/��G��2`��������w0��E�?D��ȟ��B��=ۃ�'�YM��hф�������g;�N�z�%�� ���#3���?�|��Ň0��N�L�=�;��q^�y��i�b��=2c�N�A^�Hr�?�����K���{	ځ�/@�M�z���n�o{��ށ�a"��|\�;� .ni���q�R*b�߸B�~�.ȍ�yD$�H�o1���/�o�����sVT�0G�m�X�p�}�F���&Z`���})��ꭿC��T�?�wb��A�p+h/j��@��@�T�m�,P����qԪbC����G�H���;�&ۄ�����x������<1�wCHE+O���kN���H�|�:H�q��ƴNq�l��Wy�a�F����B���&�����*Bn���ӳ_9���8�x|���8��زXr�C��Q1=F��xP�����ddPVc�)��a:�4�E.54	[���.�L �A���}&����": Ͻ���8;��ι�y;c���:�C���z�}�s�dd��Y����I4��.�'���!"4�C�S,x��:�t�e�mq�T	�:?�?B�o*KV ^U��a ����� J0�s�����<-c���"������e���9�D����'��ƋC�^x!�N����a�YTXH�Ӄ��
vJ��T����7{�N=����CQ���BtD��s,�Q޹�䂗�<�0���K�v�.X�Y�@7�ꯉnL�2�u�%��aɈ󡄃�{���ń��\�M�n=��k�����XR $A�N��/���� �
?#3��k�I���"���M.�\��{)*���#|��f1�1��y��tܠ�v����H����Ǐ*�<9�"ͼ �`��ā�"�]�z1h�/1�d������ ~#�����`�^�@6ʏb�M��4�,c �g����:�T,���|'u&�B8~����좽d�.�݌�a#�����-{� ���A=��,��|�d��0dC�GkLlT����H	G���s���2���Q �Ⱏ1��V���p�E1��̒�������ݛeƈ���@{$�ͺ�J�Yc�,Fg����is�j��B�(��B��񧤉������WbG$$w�p��F����y���%�yF]e��������4/'T��L��8���Ӗ��n<^B]��Of�ͻ��V�h���2f��/����B��Jjݟ��h�bv V�~L���a��(���֢�n6��*!JQmS�e�׳m�?��;H�om��m��}m�B/R�o���t������.�ԏ�i;&,��#�x]��@��r�úT��U= �~j<���#V�[1 <hs
]g;��3�3���@IMd#w��4��E7�!�Y�4�<�]*CHK��n���Y�Y4?[2w�/�bVI������\�&��?3Ǜ�՛%v�jE}(@6����ưfoU�KN�1�v�PoV��&���$����d`:�ͣ�RƑO��{c�/��B�P+�i �� Ճ �2���e��_{6&ݦ�����=�) [d�*�ܠ����F��x��k�9"��ڋ�{ݑ�x�'���*�f?�^N�Xٜgλ!��Z����*&�JdSN�[���K�L���4�*w����ps{�&GeIS|�e�f"�Y�|JM�)�W5�A`ƥS���8K#B��&':�Tl�	b�/�]�,�6:���n���V�����B�Tc��A՗p0P|��U&��(���6�>崰:�LW��?6������%���8`ҏ�n��v�Gw'�&�����=���1�;�\�ȣ�$�1�K�w�w�����g��R�l~�Q�ң��W�W� #�.���{?�H��cZ��5��"VmrB����P�Q�*�	a�D�mJ=�x�� (~�[���_�v-�GKJ'�Ƚxb����?�pEI�]B�WOC�$'6N�
M"Zlk/��Bӟ�.�'s|�:Z�����\������ 𑵌��\L���N��n�;1�8F��]cHz��C��N#>J�&��Ş���\��]�d|^���,�ݻ��&��qW�90²	"� o}|mvg`䋏��|pɎm�n���B�W8Sw�(��%ڕ`1��';��+�f}n�/oE�(�P�ױ֌L���ê���5;�Iݺ�wk�y�*�q$�G��n����Iy�s{'7
b�0C@2�\�b�kн���
wO�[��'��p���Kn�P��xÏ��eͶ�p��
�	V�����H�E�m����<ǉ�hx]�j����_�$��N�ϗ���MK|�r%�Q��g�?���^.p���ݓ�k���QUF�'���۶�J��lYpFm�o��$���d�Ͻ����OL�:���T�v4vԧ���N���P*H��<ϲ|��j��%`u�Mn1��/~���!�~yx���:2E�v�^�8��֩�CVM&�,�k�7��s(��~2Ǒ�F0s��r�20��:"�,��>����-5Cm
�&v�3�hq*��ܜ\�k�m��t�c��}A(#�z�����%x������� dJ�����vQ&N�Q��8)�h�����Y�r�����ɗ�M唝��s�� �i�|��;���J��_�u�3y�cH��X�����S`�+�n�$��_�O����Z�nH*o��l[h��q�0�4��6��	�*���q[��%S��b�.H�|��-�6��
�c��	z�xU'G^^A����_Z���
���D����U��4�+��߃~�+xь�˭�8�iB�>@HQ���S�R]⃝�%G��Qב�qŖh73`��i�����<l&���%~/z�y�j�%�[�NlU��hr|�Y���W�y�j�J5ܚ��i�Q���/<�����^�ky(G�o2��BO8��)�I��{���K��g2%5��^�h�р�r��5���[ �,Q.�<u2n��6���������⨴ҽ�5���_K�˄�>/�ܘ�W^���C��!+y�J D���C��S�Pd��5��sl�p\Q+�SD� �GYt1�g@���/����jsY2g�~�M4q��V��u .B3oTD�w��{��i�����_Z%'F���i�9mEH`4#M�O�[ݹՏ- �y��!Y>�^�� �eh �����~��iQ�������U�����w��^�Ze��S����"��H+��p_�/Μ��MEU�zT���i2��F�ӣ�c��b�J�������ɋ+�=�e����움\�߼-��������C�GXv��b��6:yZ�SwO��hA{�$,�e:�+��Kl��
�,� ��ȐF�[5�6�e���xZ6	�Dy�w�����d>��X�<�9_�;?���m��ūR�Φ^�)6f��#�,m�k�(0��\I𫪻	#@<��Dpo�0�K�٪���]H�#L��RY��:$�����:X�����2�{�9HyEJ]^�Po�8�Ȃ�x|<t�5 }��ˮ�;>�dP�f�����S&A��}��m�7��i�����m�'K��������}`��b�>���j��zDy��7�x��4�6E� NNG�Y-�w�$�Z��+��.$���Ȫݎ�!7�ΰ����uB�ލ���X:M���]9�Ā.�P���L�V R��B'���rN�aIs2ʝ�ֻ#���KHAY�gt��C(چ�M����G�I�!�[h&K��{'��9�H�8���b܎������j�g�_�N>?�ݰ�T�C�%4|��͛ʡ�+�l�_n\�Rƃ�bʜ����{����w
6�.g�ݚ���ĺ|���O{k�E����D �JR,q��fg�%���Ki�c5�*�S�,�s� w��6�D�-�r*+ڃ���9h�:On �t�+�j�s#���;F��y��C�խ>ٿl�ɬ_�k�9E���)4/3�7$$Ki�T���MVį����+"4Tw�`Ĳ�tI������w~Oj	�@�䳙��]ݛ�f3�t`�&���K�������9�Å�d���#��Y=F�_����)�JF�o#ŏ6�[�)��$�P} �x��S��}��	!�H�i�*�wt��eT<��g�L��G�V2�^�G܊m��a�w���M�"_`�q��܌�.R���u�o h(�;��\7�Š����~�����H�Wphl�#lL�mmvtgm��EO������*��疧d�A�F7����\�%�*�+uj�6���/0&8q2UlA�1�Y�qH��uWZЂ���K���.6x~A�����tw�|X�ϠL�4�[س�!gBq��9q�ta��PH����C���+��|������!^�/�����Ix�����˵��Tʀ-�~�q��as��C~�G]2����#�. R�-���)���6@Wn77۳b ��~%�5�����f�\%�"� 1�,�p��z���B�R�m\+�#ʧ3C�ʝ/����aʦ��S,�^���ԓW�����oso���H[̸fz���5���(��M�{|c8 �ş�m��Awʳ�Q�^�H��*&5C��1&Z�N�B�4@�&/�{D�e*�U����=���s�8�Y~�;�Ad��X��G�kjt^7�{}�k>��k�K�֡Z�5�����`�k��y��cK�䗏}̫~��-�ֱ�Ö�{���8y� ��-������
`խ1eì���x�*6�9���߈�Bc�F�(��F�Ի��7uReH"�O ��+�
��x�"ϖR���6Ұ z��¸���=�7�:�Ձ2�f8�le�#�PM-Mx��d��4��@�Q9G����x�rU�v��\�F5s|�y���J��n�f��`G~�I�f^�_�O�f�{�=��ݘ㐨�Fd|�/�)iCA���������D֙`��Ϭ?Тeh������1�F�к( >O<mT��v��U�¼̠X����#�<[�y��Ib��G���LN�9*-/��֧��+��ݏ�2�Nx����e�v̭m�]%5���}�|�tv��}j�no�{�/��bԿ���� ��6c��2�-��_I��Zx�>���M��^Q�G�VV�^-���I��*ԕD:h,� %eB_��\�[:&�zj?��-�7v:,���u�a�U be1>�q����a1�7�?Zo.�5�x��;�%h�=�#���6a*xt���<�(��@�h���]Hh��+��.��~�<�F1�Y~����R���ծ	�����e�'Y�Y�x�B�O�@�J���m?�j�5]s%��#x�}[6��$E�ݖ�,��W�����c�߭p�\v��v�����?˛:��gی�b��'B$?v�Hb��ʭ��0�Q b�t�O0q@�M�ϙ
�{��ɮ�Vm��L5��	_j�o�g5�I�Gܽ���$[]w�۷�	�ne�<�y��P�kW����uX�H{G��1V�P=�S%噬-bt�T'J�)C��B�&тck��GU?��F�k��,!��M/"�3���˴X� 7�F��������1SĐ3OO�(Y�sN#{0V�tT�\S�3ғ5��xn|�ybeR�N�ϥ0�9^����7�zG���^�o�2ǜ6x�"HA��:��o`!t��]��0����%d�k�ٙJ�(�v�b�5h k�ݕ��L��j�vm�0�����|ws�t�i���o���#��
dƼ���F��R�R�]%%9��i�ox�2��V0$�N�<�'�_��wV)u�X�����f���b�VA.���T(���d��=��p	(�T�=Os�c�H!W04C�g�^`9Bf���vӛ�s�X�R^����Z�a!~����FsL�a!%�D��j��R�o� �E$/����fC�����"Z7,?CrޚR�'���29!��Zi�1���P}��I������8���`�iS6��]e�b����X��J�D��&߶o��n�A���D��&�7yRd��.��c�-d�:(Sp,(�5=��e֓�Tf�v�"+:�fAU5z47#�>2��@]��EdƐ�Uy��lSd���*�Bw���гz�mA���{.Zmm~��{�L�@͊��x��q��ce����2_'��گ�=,����FI;��{���J	��9��{�7�hN�tj�ٶ���6�/k��J곻ҳ�,	�s��>��S����~y��7��۠Ye��J�kꍧ����I���`�x�9��5�Ѵ�E4�X�l{���;M�n74����`<�G=ȶw��qq�="���T@�����	l�R��N�0��ly�H���j���!J��J��U�>�rv�3���..��t���I�-H�xk�C�p.�Jg3:x���+#V���KW+x�O��z14)�F�T>h
.]5�fv�����E���Ư�z-��/����K��b���{r���a'du$"&���w�� �dwG���o\�(PP��d��/g���q�I,݂�3� O�4�G��w�:��4|�$��8�c����V��B������ۿ8�s����ߡ�B�ϡ&]�H�G~}} !fZF���3��`B!ETZ!�V���b���� ��:i�I��{�k��B���<,/��a)F�7��h�h�C��I��!i�����F��!]*�(-��#PaJ����\�9jA*>@�UK3��<��F5q�@$V���L�5U]�g�D]k�C'q�>G���F��k��O���M1V�«�T�Q@���?���U�D醲?*),t^�\9�կ�#�K�1q��W!&~}��d	Pӊ�` ��)}�zg��c���
c�-31ԉ�gԟ�$,;C�p��o-��e_J��U�����X�޳q��=bO�[&w6��p��xF�r"��& �h$��h�����7�x��f\���xŭ�f7�`ˎr7�p���/;�~^�>�l:��W&3�G�84E��ƻ�b8��K�+]�"%|�/���푤�W�[UE�H���]S��z�T�e0��9\,e/�"�-��oQ�t�O��Z��rg�8ܲ�:��ē⟴�,�կb���74 �����D%Z�R4��n�'韛O��@�+{R-��_�TV�`P���*�g�XRE���#m_���o���+&q��tX���91�O^BՊ�� ��N��a�A��G��I�;��U2���^�_��R��F��?Kex^mrJ���h�r��a�� .F�v��Q��͓�l��6c����8�|������JM^Wp:$�l���L��Z��&L�t�1�=�:�X����Ȟ�pE�|<i[r�Ԗ"='^�M\^~9*8��9����
���y�D�񩠕F����ɜچӻ� bٲ%S����i?�p�q�+��,����&��U_�	%j�qj8��2u�Lօ$��cW��+�iw� �3�a�e��d�4��Z��i1����8��
s��j�̓����.%�R�i�ql���K�Px�B�g��mwR��e���	%�l�ꃬ6���Hx�Ba7�W� �� �+�/H$�ܟ3�j��N��zS����c�ٕ)OCSi2�W2�)Z��:3�1g��ʵ�V��$��Ւp��{��w.���(��r���;�=}�Fr�2ś�E���?�[��R�����1�U�����vL;t�iUmr�먿1Fف���v-
�v�L�k������H�H#a�����D��/Y/eqŬaR|o�T6�����b��d����	t�02��Y�!Z��1����F��=�����&��q�Zj}>�ܸ65\��[e��ϒ�Xg�E��G��h-K����0(�w�#�scLu��'�&[B('F�k?EJ����8ɭ�v�ؖ������s�W�C'�Uh��fz�`r��t�4 �ȁ>o���0�-
�`�e uGj�ǖ��ץn�xRw����"~
=�2���"����oC�F+��̩���I�E�:RJo� �~s$�q�Č��=��ż����M��wȆs���/|����?Rp~�i�\�Gpa�8Yo<.���O�Sg��b	1�*R�$���o��ƳU}=�w>Ϩ�O�.�������"EQ#l��j]z����1&�������r�̩���i�d=��'	����7FbE����u�!��S���X���x� `q��Q^I�Wޘ�a���:�R�zJ(��k�O\�oM�L�w���w �-s������J��on����Pχ݃�!�.i~M�5ne?p4}D�����AP߯���c�v��F��ę�����jb-Z���M�z��?	������6E�ux�p��2�I�{�����pĘ�jz�ګWh��pL�GW�b݀�/5��aY��F�xZ�hD*БɈ&�)
l,D|4�S��$S�!�}V&��w�|���+<&�zl���bY�����>�j{ۺ-oH4��;7d�<xb�o�V+�p���4n1�d�ͽ�e��3��!�B>r���U}�0���J�B��s��rZ��m�C��#o�x�����S�R��^Mc����-)�Dp�$T҂%<Ţ�<N�^�@����f�+GS����8���2n`B�r��ɪ��h	�Zn؅*�]!��@�	�Z�]��Mh>�ו����k麍ّ�Q|R�6)ZKAg���iqf�;'U��O�)�J�x�rL��߹�v���4�؋�iTX?�ŏ�0u�2�Z��#l1q�!�]�c�����8&�-N���G֙��k���pG�},�!