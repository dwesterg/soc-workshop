��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���۰X�cr��	ɹ�U�����60=�ܱ2��-utTXfϕ,��r�ҍIz/k�T"̴�2��o>�a���1�.��n�~�ZIc��\�2��,���Vj
-�NU��&�m�T��剤��&(?\�i��V�ӌ@�I4���vd�����,if�Q��3|�]tw��7(��zzݮ�CO{�դ�L�h;8،�ֿg�v����ӄ�9R�*�R5_2pw?�_���{rf�V)�2�;p1�Z�Ŗ ��T�ߧ3}_� ��O��I#�m��o�O��kxv��ި��3���ӡz^�-$Ǟ�ʶ�皘�u0t$����z��jSU�J=t��8�cF�.��\�4�Q1���Iv|%����e��	��g@��2yb��+�k�+>��PπjtMܥ�Ξ�$�	�����*��.�g7��V�R�N���3W��'��Ga�5��u@�e�D�v��.���5�΢�ˮ"�$WՃ��k�B|�����ל��WbR�= �d�_��W���Ii{�ed򊗿NQ��kP�����_e_콆Jc�T���,�ب&��AS�8����y%��v�7�|0�ێA�
�J����μ �A��F��8���Wb1�=n58�O�ep�F	��\��'Nҥ@�&G�� ���{SzQ3▸��ce����ɖ� wKhRX��m�I)���8���
a�1�z���դc3� sC���������؋�ՉΞ=E��њY��g�}%�ܷ�Әo��o����H ��4����u��G��J��&�]�]��>Wm@b՘�:@~�l��ݟ~�eq�	��TRw��,��a��^9�gr���!�j7��;V;I1(����֐�������5x�0)k����1$���<��CHI��gq����v<�a�Ly1�㈰v;ٔ�v-�bT��)[@����@�dfz ��2�� �����d��PgM�nͽ�#'�k^�oJ{��)���O�Nۍ[�n���ٴ��?�e&+��֤��s�M��?�/�!��z��X}���:Y(U�S�Y@�S :k�2Č�rN�-���:���X�f�`�!�����72�Y�&ܱ��J���D=��C����T������s���`Kx�f���/p�����S�jE��z�*��*��c�3�h�B�p�q��=��ᢵy��i9H�+c¼KlV��}�%Q��F ���ٞ��׋@�ֹ^m�\���^�ǱGn�QBP�
ma�l-:��,�5��r���\���q~v	#br`!�d�){ E���1b$J�˪6!<�|XfL
�WSE��	>Eo�\����G�3�1@ƴ	�)q�-$�����(����3��Y�`:�f��f�	�c��e�G�����IX�>Rz7�T[���C�ms�k����H�����n.����2�#��,������V:#Z�ڕI�g�5�n��%0qY�)��mI��$A�l�-9HU�<�(u6a7N>�[QCr(�EX+����eP�_K2����=#ic�}}�g�q�x>lSNl�o��9V�j�/'���� �-i"C�F3c�of�d�|)��<^H�TXS����?,eL�
N!l�vGf��T̶���!�>ye��'��p��6;��ap|_��]�B]��
4�~�J9�b��9V���O���:�5@��D+��h�k!Mٌ��9�>�R�߂N�aR��#~�Kj�ƥ����)4x��4c��o�:J�_��<�=���u�q���h�BS�<<93���K�����Z�p��2Ru�hPb�7W���H��d*���:10��qv(P�ڪU�j|���H/���!̌���c���",�>L�`Q(A��UnöF�H �c��`̓�w\��w���n�.�!��-�`�T��}]_��_}�4���I����.�3F�F�׷���
΢�����](UԷ�yRn�*�¥�Rsq��*l�tem���;}V��I\@�&5<�d�ɐtI�J_F`�f�RL]|���JrWO��P1B����=�=���S���m+�8>���
	�b�k�q��G���$�7�e�P�W����-�nR"D���Jz��qZ��
!*IpzG4�P'
u�(��&��_�λ�ޑV�%�<�~�V�e��"�!r��f�r��м��ǒq�������a��x��F>��	J)���ڛɸ%N=}�+����-J�n�:ɷ�mN0���Vi�%#g����J�ֲ�|�g�����W��K{{ ����7m,�Qy�M�[��k*��b�����E�=����g�WR��`cx�`

���ҍ m~�b�p5�O�I��Aj�s�;e�kz��"@��;�k�{�cP?�jLuf�hn�&�?B��yk�=g�cd�6�u�JF�׊��ԩ]J�n�q��,&D՘�.OpΔ�j�{D�M��u�f�r2�LB�Q�Z�<�z�:'��UQ�HL1�Ҍ x�'5�u���sunD���|�%���x��&�:�<�eo�����V�:S��|��X�x�}B_�����|hsy_=�V:��u!�Y~�[P��! V�<��A�X*&���hFp�H0��]�F0b�_〴rF��]�2�K�&i�N:k��C���v����5A+�W��h'sA�!4��X�a�`��J�uHI�YI�A%��Th�@���DK>.���p5蟓�ЮÔ(��Z�Ŵ=j�2���@5V�>�����Lږ�{g�Η�����ȴ�њ�$��(/W��X)�&Z" �����,Y�`����-T�qĤ>�ysȧ����Wu�'���JHV���@�$�f8�T�� �T0-L�bW�������E�O^��Df�T�	�Yj�.��^l�/P�)����{A��/����&�z���	K�-sJ�BP6KnL
|Ƽ�S� �Kj�M�j���a�JR��aR̕�����/�g����㻈@����D�N� �\���/�ͳ�����ʓ�	DV(G�N��~{5�_���MYh���܅�z%��sԦ6��ꙿy<�;��e�]�����1��Dߌ?'����L��7<Ah*�ܡ��H�
�$�\�M&_�%S�☩[��3A��g��V�D�d�y�d;����WwZ{X:6p��|��h��'����&T����H���*�]� q)rh������;,��Ǥ%��
�v��Xbȓ��6wh�u>�M�]����Tft���LS�<���[�Ӎ�0�����/�S,Q���/�L0�U������j0�T.�`DE�O~>�b�����p�p2/@�R uX��u|w��0�b��xS��qDD�����7�?�vQw��6��'�"r��l�
b��P�ŗ���ݲlQ��0����}��4�j��v�g1j���O>���H����@;y͗���1�1q82�v;+�S��b2�4�Tl�f;�ϯhG�~̄Sy��
�/��,�,���5U�K�_؄���}؁�A4��Pl��=�<n"�6
K�vUbUA�#������?k2�T��<)�J�=�"�M#�.��y��i�-�����s��\if��0�*���6 +}��_Ȏ���_u-���?�g���י@SSL�>��=6q 9v��^.<��//%�
�u�r�;8~�7G)E�f�
�]��:#�2��}�� �!�A�f�d��nW��v�>N����ľt�gA~1�S^�h��G�UmH1'�«t<�[3��~�q�o$�9��o��꺊���ڏ��קx�(eo�0 %-�Y�B�X	�o����zĳ�gj�"x�9�v���P�:\->��~F7x7PB�+?����콐�Y�y5O��+�y����,�+ss�i�a֭PI�)���"$i�;U�r�k��xoU�c(h �#E�@�{���~?��W�U��S�&�q�\�D�ڀ�n�^�{�\��2F�m��Ժ?���m27�+ߋ��ם�A��S�c��9q�����C]!.�^Ss��8��I��I������̆9�f���&��&�_��T�u��q";�F4�}���g����[��L��e�VZ�a)��� �-�5ZR|�繥x��>!�9;1	��ape���g?��u��b���C����ɸ��ȃ��z&���oF�@�G�je���,�3�pL�4�������Fݢ���$.1M5��aaI���o4�b��L�E��g�:h��u͎Dy\�������aG
d7f'B�%&;�)&���������O��^�C(�ҽbM�U S���kT��b��.���<C"� 	(1��\�����gQ@p�4��2k?�//.t��kMW��<r��1��赵�B�rø����	��Y�����T+Nl4-�h9I2�u��Z�S�rv7�\LW���@��$�f�%�zÚ�;}���dFS<��VUd��mD`�6w�$�4v�h��"����>3��F�'oj˅��'=Q)�euN�\u�!�Zu%�*ˉ��Wu��v�����Rl��,�[��j?o~�y��_��7P�|��컒�Mz���Q��(��͸G^)���6�z�ҹ���Ɠb_���G~"�Ǖ�?���r	3�NN2��+�	��Ya�~����^��'Pé��������p�m���M��{��>�؂iGV1�򔸞@JfA��ԺR{Z�l�}���p�X�E�^"�N'q~v!Z���!�qi�韈�O��И�DB�m�ư|pY���.YPearc�U��l9��ӿm����N&�}��絺�c��!�[Z�h�5�� �}�}>�F9ީ��Oӂ��gM\[�~���̷��	�Et;A��!�b��ʪ)$"�d�<���K;!\��#`��QEx���M�dS8]3դͮ��Q^~�W�)f��3�C���9
p�ۓ�+��7Do����K8V}*�"=����>��q�1���^V�`|��H8l���c۪�8u�o:|�%Q:����t�:��7�]�󖴦᭚H%������[$X�#dOjh�Uq��2W" �n��q�꛵n�E���M����NYhÿ�SPӮK<<;�`mp�p��Q1�	 ����R|�1�`>)}�+���o���J(��Tɏ�~9&����*��ӺF�4��)��48��e��^}��ˉK��AG��ԷYc�յ�cU0�N]<����� \���������Q�ϡt�T4.E/~tY���;����4�W�PK\�P�
B���pZLEcB��O��Q	7������D��������P8E�
���v��,�4����#�hO��e7;Yɇ|(x���c��bb��g��+5���0��.�ӊ=���4���W1��:��D<b�z"%`"W1Q`]]��sC��o�2����ƬZ�-�{!T��sAiK�f�㉑澠�������#�ߩ����$*:e�����p��ox}�r���H
��<��j��X�MB���O'�7_�ʧ�ƺ�-Iz��s{,���FB^�l�@�,��#W��1iТx�<��
��|:��|b�i��V�X�w͑<�Ʃ]j��~�#*�~�;���yq��ƌ.�AE��Mj��KĲ��:�N�����ɒ@�[�.�T=/�����:�9�@��h��#�Gm�{Z�ԉ��
xȩn�����6pU��4-Q�M�>V(�R��Tv��X���� ��}�$R��!*ߺ�`�ݯEz�6D��9q���f�%��8�Ŭ� �����
1u��
��O�����8�\���Й��p��xA�\�I�3Su�ɜhs�dr�}O�Q��b��P^��f�	g�N�6��Ъ����a8������� ?��>/V�d11���RF��q�?J@����֋1��x�u�}H�k)h?vJ����}sЊ���]�1�_��� ���Bbal����qd��9��ej�@ާʽ@��}A{X�XMΛG˳��E	��~�4d�Ґ�j����|"�
�l�����\���aOa�)��t�v���J� �H�qz7K�PW2���}}���R*���f?��d���3n�:a���ŤŮq�T����)��D�ַI��]�^��[�^�SHpN� �c�(�"�"��A��6'���B}�5c肆і%�rc=��iL5(�w+�x�y��m'g�����������Tje����MEm|F������x&X(�!`�V��oYC�&��?�4�5�=4����w��U9��������%�]��3�hS��'Nh�����"e��2XcC��'����rj�7�|WZ���r>7�f3Z�(�%��ޫ{�y2}6�pΎK*nm��l௾c�$����2={��R�?6PFW���m�cn�	�4��8�b��~�N׋A�i����mP�L�II@*i���A���+�AZ�|Q��Jkh�\�W_�;+i�WU~R�@�%(�B�ü�s������wz��� )�I�C����﷟h�"ʮ��q��`�Y���K߳wn�;��%��n��Nd0�]8f�=�O������v+:���#���úڃ3Z��\N:��SQ��5n^�V^O�rUu'\k���cBI�W��K�
���C���_=�c�.�O=�pc�ȇ�d���IT-���W㵀Ä��)n�������AG��<)���vJ�aX�^AȔ�� ���v�82(���GH3M���	����K�D�Q}�7�K��TG�=�(��c,L�ܗJ:de��f4<�b�����=D�~��D���p�g�*�c O�W{W��9�Pqc2}@�}�e>�S	��:���UB��x�)B�<ʰ"՗��MB���_(@�ѫ���o)�>��~X	�oI�є�zI�Q�Q�8 �l5I�&y������q��6��*�O�E�>'����{uz�w�$яV&3�"�Hp�N �)!還Z
��>2d�W��_y7�y��t&�k�ڀ.R0QY��t�ܵ� ����HZ�t �4��{�gFs�KM`����z)��Z
�� t^��F�R6�T�{Z��1s����l[���v<=�ȄV�g��+���X�^D�@�[�2�+/Վ�t�6Pm�? ���[�g��18m_���陭����a[�,*@�3�^@�Ry��Y�j�v��j��
�1�l��?ݺG�N�%�CR����?��B)q��x��9.��5��9~�$�����2k���
N�ق1�I��[�
/v3��6�H���ڕ�������($oW�Uwf�N��~��1[��e.��5�S�#����\��Lt\��6� �YSѦv�V�V��@T������*"/.9�ũ�?�#7�DG$C����|&�Ɍԍb[Ҳ������О\?���ҧ{�����[K�v--�H���g�9�����#�]����W��!$(�P��RxY���*�����{�K".E�*kk�z���4T��D�@c�);y��^Rﾵ�� ޥ5�̮�td���(�c��b����>�i�mEs��e�h<�W�r�k{���5�,3`b�n��\���~��K����z�0�������w���"8��A�&9Go�s��t����,��Ԛ���C.|�@d��P*��T�q����� yb|6'�q����K� ����z"$\T�]��?L�O=\� kQ�=���ʧ� b��h�3�A������]��f��tڞۈ؟�����P鐠��(	]̞[��K�O$y�r��x�9�A�;j�s껇g�h��\�k5Y�|jqC�Z��waTQ��`Xm{
��)��W8u)s�d��<})?��V�
b�yY�1$*�!��t���U�p;0��+۹�f�wx���+�/�����4�J5-ۜ�8S?qNꅍ&z��s/F��	�ͮu��D$�C�9B IP��ˋ��+ܭ�	��v�U�ϊNu'�W��L�?������Q6	]��-����ě��jו�T���$X8��+�o]���O��/��u��t�SJ���D�O�>�3r�G���k�5ϙ2�M�OY	(o�����Ch�U���A��3䵾.i����l�k��J$�룃�޹�����J��c������
OgH��q�Y?�_ruK5�\��.�N2eZ� ���Q���Sh˛��x��U�,{��ӵr�-zZ�i?E�}8W(�	�$P�e��*��RPb1���N��� O��64
�\K鸂HT�0��g&*?�vL;!j��h*]�����4���9I<��=v|bsFM�=�vt��t�G87���јF�G��SqJtߴv�![�p��aD|x��jT5�k��[���!jZt`*n#E�[��f��i��t~�Y¯�g���0���T/�����`ݤ|Z2���nቧ��T��t�M�#��c����Wn\�aVL´��`-IS�c(O�$H_1 ��$r�*�F����i�g=�e��v4]����sT�gC��^2���i:2�LJ���(V�,9�� �m�3TOpq��!��C�� P��>�K27s��6k�~�=v���Gj��-��sz������\�mu�f_g��A�Ϩ������r��瀵�p��v1%�V��jP-Y�Z����>���xV�U�e��U+rڴzGư��.�L���$Ŝ�B�����������p�^u�[3�~��qn|��_M��t�1�i��3���Y@\���[�W�|�.Ew���n�=,�5t*O=�(�����&�Z+ue��w�Q@�����p��%��/Y�D���g����T�E��!��!��r�q'U��k�l�|^NC�5��nb�s:M�z�T�=�<b�.X�C�|_A}��S�]�/�2�
z�|�����s�
B;�c,̕�bŎX�[	(�x�U�u��s�˄�}H��jl,>��D'���x��Z)�g��}ɦT=ڜhu�!���.����nK�;�u�Vt4��Z����@�t��bz#��Ĺ���km_GM1��j|�)�hv �[9!�M��.a/��&�͓GY��W8Z��(�t��S0I��m�d��e0���.$-���Ɓu ]|�d�;#ìÅ���
�Bl{�3�1�0�.�7Y,���6��i�r�l��	h�S*I��ѰvRf��v:�;�^%w��B�������\0!��jrЎ9|�"�i�vJ�;���/�\�"B�#AA�{��oKaC�0��M�\�:�=�ߑb���:�����(-�-j\��ѫLm�`�=O��ė��,� K��XVq���*oi��	���u�w��o���@�K�>#9!�;�\�5I|yEi�F�A�7˃����p�J�c�`��t�`�?Ǿ2X��L���]�a��g1�K+����B#�'#��3��S��- ��_[1����`9 �M1�pb,������C��@�T���OmH��Â0g�ָ͜.��m��8�r����{��FC/S���T�%���8�IUcZaE;;FȊx'X��*��:ALFZ�N�{D�s \�؀��J��Xw��\nC'_㐭'y� ��I������@&On�3�E���@w�2`NC�p�x�d�O��joh^}�p�Ufc �->��k&���I��h��b���|H=bTέ�}j��	�C�vÈ3$��櫞�o�]����������E,%�R:�L;�j��`�{N���aVD����}����"LQN�o���cҭ$�	���T³�f���(�Gb~ݳ_ʩ��e*��Ȉ>+�i�TE�a��-f!*&|���p�KGqT�B|��-�S/�85�
Ɂ9�� ��M㘌%k��YS�!B��Lb!	C�Ù�ϭ���RS���.�S��� ��?�]��9�1��?y�F��[52�N��蚉q:�8fx �$PCCz&4-����<c�	�8�T<�$�f�)YIPs?�����-�MNsG���[̋�2���E:c�Z����)�
��� i"��K�%Q��@�bTz����T�槞`O�=�C	1�y�$s������
�T��N�� ʹ����[<�X{ӧ�59u@�'�C�*�n��b������=T��~4��Op�:+���4�	�Sa��8c1�=��44�S'����Y� �v���Mъ��8�Z}��|�۝[�$��ܶ<^>"9�E��3�jԯ�Vk��?n����	�ul�QU;Z�kp%���OAQ_��v��ݾl���0��� ħ?HUm�]Hb	}�L�m*�~o? z÷������6���k�:�8��@����ղ�ޔ5�v��6V
��\R��P5�����]����	��5���_���+�w�%������1�	����{��c��Lt�����Ü<��7||[��?�� �3r�}J'��8b��?����4����<[m�#9z4�-E/���п�l
X��ʌ�8�{��j�m�!'o8ұ/U��ɰ�L���ё�\�W��)WDf\��uH���RI���j��щA�����U��t�NG�7gtcٝ����]������ *��u��l�uƴ��2ֳZ�71������d ����Iks�P�,�GI*��m��"«�}�&��	ǝ�