��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g7#���m���4�2�%j�[g�{��-��Y�\'�6��`<!Cu��l~��`�Ķ�������x�#]��b��^��B(�������>�[0��?�<c,�#P1[ݬ���Ak[��߮��h��%����6�O��W1+ x�=�`����0- ���KMM>bBS濳]�1�}�{t��f�%���4�[�F��.y�x�6|��;���9N�ˢ�eN��TݟΚ�YO#"�!�&D�f���/�_�a���|ܾ��U�f��V�{j�l�Gu���P���"E$�ջ��eo��2-]5��nR�<4
`��R=��R�?�Ų+�tvKˏ�](�/Ы�v[��-��������.��.ن����?�~'+*����U?R�5�D?(��z�)dEdᅇ�+����J�[�K����l��ҳl��ۀ�%�y��w<hD0'W[d�Ҟ8J�����k�SZ�F�>2�%!�T Ud��2��b����)�GX�'Z@+���4ETj�/s���������������|�g�s�x������W��ki��F�M"��&s���uɹh��r�|~��Sm�[z����[F��r֧ٙ���!�7PvkQG�2��+��CG��!̢��f��%~L��K�2�ٜ/�t���޲\�vd�mT4Q��BO�Cʐ�(�����H�@!
xa�dk���,���1��#�ϧ�#�%�<��]�LM��2M����XEnϲ\���͚7�PE���W�Ti}q7�㙦ݞO��Ի�<|�����y[�+��E�deMR���5�K��;����?��ԞQ�I�ݑ��c�3�˗�|&y��'Ux,�P5�]��n`gA�8�͇Vy�O\��rl��U�0��Y#�1�O	s�)���ƫ>��"i#�mD�|����x����]��a���Y��8"&�T��i+3�?�w,�K�.m#��8��|"�?��+��#}�o��N8��/�&�V��!N˰��3ĸY��V�D����ExWvrTPm���[a9�G5�nc��T9v>�?�7��J%�V�;��"]�y�u�Z�A4f_�>!�G�\qJ���>UT$�T�H�軈*W��5S�7!�����3���Dg��ٸ�7��Q��(��H���j<I���{.)!����6�8�Ψ);8e���m��Nk��1���
�3��~��E��f"q���m}A�e��ĒK��:͖�S��(w��l}I��ЭT��C�Z+�l؉����[^�I��i��O`6Su7AOU6�A�&R
�aW���5Q2(��u$5�`��j�8R��W��8�@x�;d�J�s��\Ӯ�vQ�9q���`�.��Z��|�����TjP���9�"&�W�Ao�x�<�t�s���j=C�%O�~ŏ�_d27x
���q9T~�9���o�A���r}[X<��P׌Д�=*c3G6o�h���jY�rQsmW�-�������,��`�8 ]Ӕ�Y-)���8��M��@8��yg���^zwOQ��Ңv���P�d��6�����%vU����m�&�3������Ǚ9q�,����ix����~2��*�.�$����7i~�T���2�j;®�U^�;�!)�e���J>�3�F�-&3��R��#�'��S7�e'��oUjK��������6�"@TAk��6����[��� �*K�R����Iewq�>�MyD^7����ty���#�h�F�k��b��6)O䖮�[' x�+Yi�Mj�j>��%T;@�U����.�C��8�a[����´�7焪�Hq��ۯ�"�Ϧ��MnF�Ӑ2=��7,�Z� 9a�,PEB����z����8d��k�yvH����X�{�R �X(�?�e<NTBD�P��E�iW���%�c����}�i�y�uE�~FjD	"$&E��:�ˑ�Ɲ�A��9<NMg�#�YM�����$��e���I�	�"�Y�V��й�AE�NG��}^�l�&o��.���bA�	k�c�ٵr�rD�?7��9>ɼ��fp�ft/f4��"�k���+mUb�W�(=$>���b]���1א����֋6�ˏ�b�e�9�����B�G��d��JudeB)�dj���@�;�>5�?cu��#b2=Y�4�n�{�g��ǅ�)�O��e�B�ˎf4-t�s�nm��b�ZS��E�1HWƱ�q+z����
�8y��#82s��\$/�t[;_�>������M?!y���ҷO'���wA�2�e�n1���Vb�r��M�
A��Rƅ�X������ɒ9���Ǳ���8�$�l������%�� D������
v���\>�)�Y&J<�^�m���R�Ds����@��V�"������t�}ί3�2'��ctT�z�ë:����s; {2�k#A�<9� b�g*���?���MY<'� ���7����E��·"D�����c3[�8��1�E�HT���x��wc��-Z�Y]���WG1>�"*T6�f$k��3��zc>�I�f��;+f�z^B�U�Lѫ�#��F_ �)�9c�ε�YP����z��u-Kh":��af��"*���!eh�䒚�ߘ����|[�q-�T�R�B�[�^�q����5���|�y�Nɞ�m�S�3�P+��4����5DF�c
���td�k�ָ���2Ty�-���W'�Uy��{�%��'^౼oR��o�y��
/���vɏ�1�+�	S�\������ϱkuP9h������e)�.���B��t�x�K<�!�V�۵)|��u[R�`�5^�I�=O��n~�a����6ԇ�Ȫ�P�=���g���̯���g'�~�W�Zy�RM��ي&�|��nXpe ��V��<��F[�[�/~�5� E0��[���6�D�i��X��4�Ӗ��#[E�H=��l�ҚMq�J��9��1�b��0���bFRݞPjXn��F���JM�۫%��l�8�U$����=a�*jV|?���F��C��Ȃ��2;?xY�Rd����X���g/Ėҳ>b�E�1f������~q�Ô��G�wg���N�aoܨ���v�"%w켗8��_O�1�:��e����S�?=�f_/�x�~>X:(]�ǂ�o���N����4.̝�D<���Io��r�GWYQg�Hk9����Oٹ�����G��@�|O�U���0�Ai�w�
�K~�`ϗ��s���8.o^��{I$g��W Y�b��+|ݘ�|[S,�� =�g������~���Y�nR͈u��P+��?���4x� *�{�1@�b���T�:"�~����ѥ��}~�>*�7���sx��s�3	�!;_���Q�׻ǭE��5�N�d�
�LY�_3�`�M��E�5k�5]6(�P�����oIި�-u5�Cp(��wd����Z�AJ<�0�?���":��i�b����I��"lK�Tte�
9���d�#*uM7i����h�v�Aea@��#/��M�|����T��!�j(DuӯZ��6��>!VX��pC��<�"�Qn/)t���7�m\ѐ�	v/V��:~�s�"��K~�V�'�����3�W��_��Υ�T��-d��tg��&�-��K��h5�� ��<=������T���ƅ�*,0�V�Fj�̪��A�-�����/�w�VJ�wV2;g�BSD�p��0>�Y�T?���gN�#�.��́�²�PG�4�7n��{�T�VI�zbqT8�vd��'���h��O<#�ޫZ]g��S��|�'��F9�9���hdG������I͜?wO5.���RK�ӕRl�%Ȣ�>Z?��y숾��j�YI[lM6)����d�1a��W���m)W8�~��Ǵ���ŤDJG��nb�=c�
�#W��U��T����:����yK�fA�r��[���	f�cui��`���L!litm����*�0<eL�+!��q쐘2��[�Ut$�Aԧ��w	T�_Ў�d��
��o3�I�F=�NXSgC��=�T2�^�)9SO4���!�pSI�j�S�7���A(Bu%[WQc}�r��S�m۳V*6l��D?#_E��D>w�ԟ�QG%T�,-�]��7kYa��H������֘�]�3���fTri-8/}2��xQ+/��Q6�u�T�F���jX��&��Α�b'��6~���r����<���:HX�r�h����t���{���5�UdE'�;+�2�w�e��d�f�� V�I����>e���H/��洠�mKShq� ���ҋR�-9s��Y�"�-�
�x?�d�=7	,�k��o{��J�Y-���ym�&���#�*}8#�Ź#�qS�k��\�W6���)�q:���F�qɶ�)C��=N[_��u3�flB>@��yۖ�:!B'������:�,���xL3�1�#g�of�*�+=ng����ZY�B=�4��Y��]�1����B7��P8�$^-04Qǲ���?�����,z�RJ�ǌf��eD���8�n_�	�4!���S� ��2��]Sf��?8�rp�U��tHL1������`��X��׷fW�Ԓ��V,F3OCr��ڷ���k�m��W�ĩ����P@pq�e����g� �*�ؤ��J)�.�	8�-�҃F�������+�4K����`�ɰ��Af�A��M<04�r1��H2KH~��F����!iKOw���ho��dG�� �%��d�A�4�w��=�5K��X��n�y����������!T,1n4 �]�{�4}�4� ��a݌<�ŝG6k�G��쑚i��XM�J��������³�q���gkd_?V4�'u��R~)h�g����[�#�BK�����G�xip�H��p��t{���؏Y̡/�	��km;�b�^�ď�����-�gW�a.�X��/�;?�>�[��A�HO`{զ�i����Tl�.`I~����G-߷zcc��3��-5�Pk�h��>D��<��Ib:6�z�]��Ca�.qT�M%�������^�=�$y�+���	,ŵ��5�Ա�<��3�?��~oh4x����p��IL��A�RZ��m��Y�;��8G�vY9���A���
Bō'?�79l��N��&����N����Q��l�C^&�d��RSͣsצ.N�7omH�~s㼑�{1,�M���b0C^����K �P3��9k׊Ǽ-:(��8b#	W�x��
P�8i+�Z���C��ɖeZ�q�=�'���9�5�������0���Y#Y����s![ol\�{S�@D�)M�0E�ߣr�V�j��IzH��i�@�����Acծ`rL���A�|B1�u ��$�5����	�h#~��m���Ԏ����p�7��ŉ�q�uyqy��Y꾐5�BSyۛ@{����q�v�q�D�A��%U($�X8!^����3O�<U/�D0r�o�4a���D��u���^��(ؕԯ*Ѡ��(-7"X�ت|� �L'�PS�Ӳ� I"�c▃�$�dWŠ(�sk 2�/�i�-�o��6�T��#[a��2rw	�X�?�� �S���4��~���<����YX6o0��=�1}`Sгv��,�+�4#Op����!B�K�=�Sv���b�uQ���>k3��5&8yD�-��C��^q�(ݮ�f-�p�a`e��r��w��)�Aq�'�LA,
��_G�L��R���ڍL1A6�f&~/�/2����]��Git/b��J���ᇵtj��Mh��<�Ɲȟ�<-rnm��~����6��Z��"hO��C39`�H?
��E9�AS����K��.�b��g"�dg��D�x������W��ZP��<PZn���¤�k����5iG#�%v���^�0�LJl�����^��^%}�t��a
��'��}���4_#@�/�<�q�
~I�������$f�A���GB�%�Ѩ�+�!��
���!�t-���@�*CF~�h���ϋx��N]]�oO�l�"g��~�9�Y}�^^�IHM~=(��8A�UM:$v��������]'LS��Z"?P�q���������AEE���Yf-�2�Lt��F��4*{�7蒏6T|�3FZK�9�d���	������iV��*�4��^|44�}�"�Y@��W�bv
t!~Db�
b M��܆�1�[�~u��,S{�x�ɬ�Ie�|����}D1�����-1���-�{���١麲K��J(/j�SW�(ܪ���d���)b/%$�N����҆��GVL%'���j���(��y��ll�R g�5P�M9_��ui��b�B#�(��$>,��0�'N�^%�����5������J��42ET6V�Z�p0�SX�"٦�]� o�7�V��c������l�������,b97���Np��p�e��b�iI��7�0�B:�{u2���±E��2s�(縚� ����|�1a��:	+��	�Yb��zu<�+M6�7�+wj�**]������׵�z��i�E�C�
��0�-Z�����:�at�n;��\&n��Z�X��b�;3�T�Φ���x�/D],�����`��/�	�	���N�meY�.�)�>��>����bHJ���f�qJ H�je��=_�LIgupP������U!������E��6td���x��܅.���\��Ӳ��+�]*��t�O̘ZLܙ�gO�=��}�{����ˏ�C�lH���z�i�?ba,d�zΈl��7֏T� N?�H˵[����}��̂j�6�%�����uغԿ82+�c������wJ�t���5����&��{r�s����Dg�[�[6 �֬6�kb�o}Cܐ˲6	�G�<�愌$�����}@�Y��3��|=�*�j�|��z�C���t:���g���j��=Rg��� 56,�J�������e$��b|
H�7�9��}��bLo`�{�?��x3_�T���a@Y��)����1��<��."����ʉ�b�`�x�zо��*���bs�W�aTm��N��2�n�����;ސE���j�w��|�T���|m�oF@>.�s�#�j�ef�$&{:��$��K�u��cѩ�V �L�C=�pg�`�w�(Dt��%c^I{����T���?Lax�p������dK1希��;߮��eea������N�k�]�+ww�A#ܧ4�+-$��׾��`(���gVE��-����p��.��ċ^��k�"�?�[�����`��
�G�u*9�J*�P&�H)k�U����`�A�wAߌ�JH�6ӑ�f`�Xus0]�V�n���|�nL�Ӽ�Ug��<�_C�����FӔL� ˴zC\*�5�\�T�ҙ�p$}����%�mF>�,�X��ow�&U�Ȋ-�l&u���NOj/9�%�C@_+�c#�p�s��+V�W�PԼ��2&u�5�TZh�)��d֦x^���+�vM�.#z��ڗta���0AN�fΧ��̴�_<Վl�˞�Owխɸ��og�6���ޝ˿��A,��e�����}y���i~3@�Y5 kLYa.=#�h;#�Ʋ$Y���>���8n��h�UV3Y�+�JLkX|������V`A��q�,�6/�Q������\	f]�V;>���g�g��*����g�s��߮K�/���G��O�{ρ���XS!�R�"��+{l�.������U��,ۓ\=3�����n�t�\�]s�p,P� U�)���[ᨳ,z79�#���:P�`��h$F�hW[KQ���?�`�7+D�`�:e�����0�sj�/�
F��,��pA�̓�]�	s��UCO�Ѵ�=��%��Q�
}����f��Dn���)r��^d�	n�Վ�Շi)׻H�6�����t��zh
6t�`�
�b�UkCmBX�0�O��
�l��a�������Au�~U��w�iNu�~N	�P*�;�tH4*gz�_b�z��VKɵ��Sy-qCe�����D��K��;q��\e��]�x�����XC��������w�K��x�Kkje��u��8h�"�E.ڍ���7@����\��(mե߸�I�RW��^��n��@h8� ��8�3>RV �����麩P�aRM�<w����ϑ'�k�Q�i�FȜ�o��|�>�PT5C`�.�9Y1r����0+ہj�c�)�~	�6����*(ٳ��S�N�@IO�a�D�?��J�*+�Ǔ$/?���"�4�����ٔ>�E�P�N�N?�B�f.�Z��p9�˛hB���,��"c���z�JJ	�����mV�W��*����M�G2&� �� d��?�΀c�4�� J�k0�C�P+3AA� �>1j��酤�Ex�9��V��ٛ�J@�dS���6>g,�� $j^E����MI�]1��'?���j���ɽ������]T�Ք��aI�).(r��V|̔�x宐8�0ڇ���	v�0�������Y�س1^�8�{�w	!����B���F���7ΘȾ�7��{�MA8#�г���k�Y��ﭼ����+ip�uݺ�f��*���cV+��������I2�1��5Yck�&$&h<�tVjiQƙsơgy�x�'�q���3%6��	�D�b��pnU�!Qn/�G��E��3��!�^*�V�p#��6AQ%|�6������u��С�mh�T����az�Ǥ����t;�e/'6`R�n��E���Oyi�9%5p����v�\��(��8�,��d|�T�ImB�^c(Ɂ6���س��H�����g"5(�Fu�UGs�Յ�*��E��KU��_	�������v7%E�n,��!bO���L��t+*$[q�4�C���,�?@�AX���P'<B	�)�܇<�.��YAqr�Z�r����KK>���[����K�?�7�%x��br2}�`;�����H�F�MR/�f#a$�])A)�a��&(���]�����O��~����R�A?Hu��h�Pm3�T�>̎B�Q�8
����z�UV�X����p���d8*M�ų��.z��<wߓB�xTT��fo*�1ӡ�H�y��i���T���ɉ`��8NG���Z�Q��$�C-)������VAj��!�0�.+���֓�eṐ��}�.��Ӿ��������`��M_!eco��L�:D&���b�4�Z�����+4/BVP,+=A��$��*��:��+Pb�n��ZJ_��{R����`7���y`E$�FKO�� �G4�>����3���kW1� ��DDN�ů��E�H^<��d9��6�r����j=n�V���Q� �V*T�