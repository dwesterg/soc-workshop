��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���=�Âe�����L����D�ޛ0��&��ތ_X`�+`�:!�
�"F��A��x�m+����{��6�c���g�>�*�J�p�K.���_�=�8���#��D��p���1��~
�X$�R�tD�/�Iij-��V[Q.yF�]}�~��[���N)���vT���Y��6<��R��P"�{�̧t� !fP�'J��ԐN"!i���w&����u�11NӪ`�����빇��Ђ��sGL�%~�۵(9���$�{�z++`�1%���N
�Jd�k`A
��o������-��Kz�ג^&O9��P`�]S�oab�%腟�)�~�_L$8��aC�+�щ?��#��%9"����z��n��f����O����S5h��`S���y���H��I3hS�{�4m�e��5!Ff���ߌ6���Ylȥ��x�!�)*�5��XH�q�
}x�O`?�Dt<~S�����Ӑ��^�s+���扚*k嘠{����JSj[�n}J%��O_Џ����<v�x�=p�N�{����������TD�EaA�bW���~��V#�����
���E��>j��݅�((b���z`AW��A(�u�l������8Zl� ��(�T#Jؗ��	Ǒ̄�g��aJA$!�מ�����l�Y����u}�¶M�;��2"0�9�*|��Q83��3IP�1��2�K�`	~Ǎ#��c�B�E���X�$�i��A�4����q��)�XGa)�.po�s,��E�W_C����!��g+tc��s�v�%�3]���$���@)����&�1`*��ou7?��pDZݗB�78<!(�7�6��I��*�[&�G:��,|�;g՞�"���z��@֕D�,���$�Q�龊�12Kq[<y����sk0�i�S�ͰXK	�a����f|�{����ޚ�:Q @�'R���}���w�i'���f���*^�iu�9+INm����s��~zl�����8L��y����j�Vt��+�Fo#W���f��-	(U�����4����m=uOl���!v'dN�qk�ۮ�	��tQ�)��n�zE���n%=���eGX��b��!k���%���ӿѮ����������w*���w84��v��Ԫ,Y)j��-V�o`8n C0֦�I}��.���m���(�I�)�3d�).#���sӁd���v_}���1�n���������?��P�f�U�<��6��Sn�s�4hs��;�w�_1Qp�L�����������C�)Y��Q�L3U;�����fL	����ajv����tB�i��+�����t�<b�ݩɑ�
�">wy�4���Ϙ��.�Qzx�5����M���b�1�H�9�,�fBe+��F���F�a�M&�8\$��Y yu��h�������.h��`4o������z{�m���I�����f!��v/L$2����j�W0 ��1r�����[P��A�4)���铥؝�J)�Y �5b8T<M�e�����O]eeR{;���a��C���x5��U.�C8=_)�a^��c�+���*m�/���i��^�Q�"wF�% ���Ut|��I"�.�-tS���V�K<G�y�r�hP��-=��G*f�Z�m�C��5�ߥe��n�JvH�Q��'�A��Xk�.�؃&k������̝��� ���D���:����=�"m�z�$Q�@	o�7
��v���n��
�?�<R��1��at��l�@��o����H�/X]#t�*
"�CFW,"E-��|����t��~�g�����q�k�gsd�\��A}S}����^��"E��h�n�4�TCAr3'��_�j�� ���6�`h�
ZL^��p�1?q�\�z��5|���g\��is�9�;�?�O�[ �.pܤ3�-��5�����|�unQ�:��@�a��Ӌ��C��Wʐ��j
�-!/�x���r|S>O���Bc�ŝu��h;����{h���B/UR�Ģ�.�-}he�X�O�e=8����/L�V0K�$_|�n�
O�&�Hh��"�J]w�W���MP����$]e_�G]�Ir�s������1h-�`=~�;�3ְ�7<{�5�΂����z�L9�y5�2��)���₌�LyŃ2�ٕPR�R1���v*j���Ѯ��_%�[uC�[���ܝ����pQ�x���[�w�J(� ��pV��J���U@�|<.܈�� ����o%1�9�[,���u�)���]-����o�]�Y��)�þ�;��J�d��T����"�`�\c�2t=e������RE�d�%��V]��3.�y�a�Zt���i"1OH���𧓨?0�;�6|v<{y��c��_���pU����x��ٽN�r��4����
f�h��A�wDA0���!w.���R`:�zb�3QJRo Xz��8/��]�R���#�7���>�`�g�\���W���Ca[ ��������o�ʟZ
�L:~6INs7L`*�$�X�=1�*�4��%{�j�I���2��jp��+6�����f#KDx/Ha�򸈩��~����9�� ���5�����o�O&W��gܾ/c����q�M�ZA�/�-óXE^�*��$ڇ[���E���ՉY?ͳ�)�$���h�[J��r����G���L��|��i����<�R�r1�y�� @����Ҽ��[��'��th�zQ�����`���/�GYcGɡ��c{N��l��%��Z<L�����|n�WՊ� �Q��/Q��3���<e��DNM��vZ�ƅ6��u��jM�AB�5�m0\%��;��J<��_�C9��z���Q�f�O��������w�Š.�X'��y�p��б�y�Ⱥ�?�(ķ��)[~8����6y�s7��ۖuD�N�2@����2���NZ��R�g%6J��-cN �3Ϲ�RǗ)��A��HW����_��"�v����,�IH�?�f�q0�m� D0T���rk�!�̙o  ��ŋ_'��҃�V����jb�~bv���R)!=��Y'@�����ɜ$�'�b�B.�J��P9��:|	�?�%�,�'Ky��ui͎f*�֍Z�!E��ɠ�d�Υ-��.���Cb�_�� �Q$���$����1�����x-�p���U���:�&>�~�Ɖ��^c<#Bl����H��F@r��~xt5(�GsK��^�e$e$UOŁ�A���H�$�������h?)S��Y�QR@T9h�1z��=��Xw��Y��/V���}��5d�4V����'g^�ϔ0lk��Ri�k��I4bOe
��t���:��l��V0��ڼ���yy��u{nr9m2��Vh�]��s�p�$�~�~ohE�?��V�U���s����$%��%ޅ	�z����Cϯz�=R�=w#�B�*@�Cc�5��m�`���88��)HR�=h.S߱�bL�c�ݖ*�r�������~F�F��ω3�w������v{Hڽ�)P���>��񆷥6����ҏ��A�&1�4����3��,� ����VqR�L󪚢|�?jD��*�ѽߐ$B��/�����=��6й8ٞ\v��d�[Eܰ�]{rm������/�y�L�3��m�0�{ݤ��Ґ������7�#�HK-jUOD�W_r�K��X��?�Gq�<� �ȯ�@����R����ZC�'S�f��n������1?��7�4�]���Z�-�M]�sh+c�7���B�~� �(��&Rk�H�	+Y����1.��HJf�t��wJ��ǭv|1�j��2e�Nm��ܦ�42j��gQ}��&p�����V���Т��G�/�ж\��Ρ`�0Z2����[�3(�҅�6��� CBȻ��&���n�D�Ζt�ܓ��>�7I�JT�pH������{ȫ�iο��6j�N � ����t��{��PTyМ=]�j�dX5٘x���Y"�*�_<�Y�Bq:>������WX1���'ĳ!�q+u▥��c#�MO ����dݺ���- ���Ki��}e�ي���D�q8�������Z�]1]�[(��a�\d�ИtK���B��m��������ss�Ң��,��J�Ij�,�X�A���Z�o��Ǉ�'-�F���lc*�n��=/�n��F�B��F�;0���&�j.�;��r"�+�,}Ǵ�a�����������)A{���q��F�Ӵ�G�{U�_�i� ���p�<��W"e��Q#��a��2k�;���[��)/����z��x�3�/Pd)�@��b��3*����#O�>}c`��p�Ȣ��@BU�}(Mچ"�W���~iR�S���Id_��k/�x���Չ�6*�:��"VP�DJ�y�����y�g����/�GT�j��P���B��ZNe��3�����F��"��>����^y�����w�͋87�x$�6���<ӏ��EżU�D)≮�?��6�%��(�zH�}���Ы��A*<g��丗�)Қ!���Y3+�Ed�dq<��L�SI��F�K��5�0�)�\�V��BM�t�8�'��_�Ľ�I[$��x{.3�M0�hz����ay2�zxg hF��JL9
���ʖ
�� �%s�� P���$���aߔW��S"gNU��E�]���q���1���tѽL����#�x	��ڋ!�p/�@������|�^ŗ�����V'�h�A�7o. �nZ�L��
��s�Ӏ5�+W�ue�sFDw�KWC���4i�j�^��|�#;yR��(ܹ�����-5f�A?f2]�5�%�~9�@"
��N@��̜�E�V�~a��9�Ma������J}� $Lj�AE��&�6�Te0E�#M��4���_�nῴ��l�C�7'�S��d�����h���!�Ƅ�L6n�C4�ݯ����8�F��р|��'�`��=62�(Ĝ��4"�C"P�Em��9J<z�Zw6=I)}F�xIJ�:���:��cE"�J�(y-��j�C�bx�ۄ��$�s��9�R��>�L˴B���E��VqaYof.RRYy.}�sVg�TS�H���g/�B�hV����o�䃕t���Q�ܧ�[T��ʰ�Ж��sJ`Q3��xڲW��m*|�>���Ċ�j��(�ܨ��ο��[�d,�֓����-,PpY�n���?�F�H�� �I��r<�ny�i#�.a��*�>���Dš�*�P����3Np"Bj\��+�
78�W�2#�Ql�Ep���9#���t[>�핫��*^C�&iG�.�z�����*�.�E���c2����e}��G* vsJKW�����'���'��Ɍ%�U���g���Ű
{�\08ûq��7���>~��2]�V4�܄K܊	���t��L�u��Ϊۍ��3pL����Ù��H��>������bM�x-�ԟ;���ZY��<[�G�� 尲hh��loNTԊ�o=����Wѐ6i_�\��	�1X{N���3tt�����>�I���w��ta8awby>����k���;�@�j2�buN���0`�/@&[=q�Ya�} $P�y<<*�;��#�N5p0��t�%�0��Q煖ƙQ�;��������j1�PD�� �8�}��?.ظ����=�����i���^Ż��ƻ����O��+q>���c� �O��d~.���^�͛�v	�(��:+��1���n�	7����Xo�~t��ئ1g��T�F@�)��~����ǡ��x�iմs��?�A+o����D@�iP�����>��=�	"�P��W��@	gK��T�\V���h~��k1A~־��ݠ�T�N�E���J99~�����k՞�~�6��٣6�Q��F�q��W�Zu��!tM홝09�)°4ȡj�=s�O#���E,��z3LVN��#���`f�]����탔d�Ĉ�K�u���q���gK�A �/��&�������{-���;N|*L�ޖ��H��,���(�AiW��+�s��PMn)vdKǴ�g*yMY2�ڢDYqx#W�cX�e!B��jpŠ�'���I�!k���RDtcU� �w�+�m8^��Ss����E5h��1E¥�gk
�9D(����9j���NhN�TPj���$�D(��,?�3����N����C3�q�RF�g�t�ŷ:pծ%tN�x�'F<�S��M�ώDZ��ٵU�X_ע�������I��5��I���ĉ�J��B�R��ZkD�C����ʑ�}8�P8��81���A�,����$�H}&'�ӑ[�,�?����)��7���?��F�.�0������4�3��ڙ _�.�u����7fh=(F�\��$�!!��9; �W6!	?R���M�F�J'���ʻ<���@�a���ωVREd�<Ժ�kW併��D�k3�$ކ"�X�t��0��t4��_M�Ώ ���T��Tv��@ܪ:b�Y�J������hj���7�4*���W�<.;Ï�u��h���4�[�_�#�a���x�@? ^xq-� �5��9X�8-wgYq*���/��BP4\����T'��Y�G2V��H����<��16�oQ�Z�HE0���\:LPH�>E���T~x Ӿr��/�s�*�� ��A�i��"�Ge^�����%�%�G�K���y��0���m��P	��k�*��;��҃�d�"YJMo�%I��#�֗�z���Z�U]�����0���N,`{�'ӌ�#�4%d�ƑJ@��q3��l��qz9��w.�Yt ����i@�+�����+Ω!g`ds��<@1��^��n���KƲ�"g�B��n,� zې_�|���6�s&A=5"������ֻl{S>��?�Q�o0G
nB�H��z�Bx'�Ŷ�j�|�'���˸7�E����ޓs$l*�ˠj������d�n_�h ���Yjn����~�J�f��Kp�,\���2[j����2CA�*��n�7<�m���&M0f?w nV���B�9�+	R8�Q�?��^Su�ZDN���_+c^��u}�2���̜_�#�
љ`�����R��A$P9��B��r�1?�Tn_�-�E���c��g�ũ�z_��k�圐.�m�*��c���(�E���r"�o]�60�f���d��X�@=�i����=2�+��
�h��.\�-v\�}x�9[�N�/���佁��z-'D��'X3��	9F4�TH:u�j���y&����ߜ�k�䭘��6Z�.�����;�O�O�O��|�+a=�!�D�އq-N�1;�U�9��fLHʩ3 ��I�U�C����c��{duT�^��z�n=	eN�ƝK;X�[5���ĥ AJ^���|��x�6V�KO��+�����X��⎆h?[���Q���%-����;O�B�߆��q��t^���ҾqK�ڠu���AU�_���Y����a	���kA���L��MBN^ދZ8��=��g}��D��N��俸+�΋!C�-��n�9J0�����n�F!f�v�c��B��O[���e�W?#vB��nկ fe�� `��6;��kys%v���Z�#�"��z9��<�My�=AF�-%��Õ���b�0��;P���D�8�P��*��uKU/�N:*���������Жg�L��5�l����P/�ʺZ ��&ߒ���j@�2$f�`)+e���馗!�H=�G@]�D�$�v�v�U.�1�����c����di6cnXQ|X�hI,$����H�+�/j�Z�;��n���#�����w-wB��:n�*�8�iKL"�;ҏ��M(w[�����VuS�炔�"���4M��
W���7�a���g�0�G�bj����{<��~pS,���}[9�%��:�h�����yG���������nT���اS�l�'$���$�5`�Q�i{[?۳�)gz�[ѱ2�p�A91DsD�>����ͅ�����D���[<x-��* �������GSC�`VblS;����F��9��u��L{�	2�WW�����\%3B��W�=�Ɍ�;�¥.;�_��긶�՝�:ﻂ�Н�}���|����gh/b@�z�C�6UK�(� �~k��vY<��F	�y�z-O�u+;�Q�L42��,Y
-$�vOܵc���U����S�9���vhy'�:�h5Jm�q�l��Z��@v@*w���31� ��N���]p��_ľ?�OFxރv��7�)�}M[�Tȣ�I�o�t-Eh���\��w�pZj��e�����7])��N���P-���LŒe*
s?�+q�.�S���M�t�d3"pbUMjt�0!�(�M��{P�!�!l��H� �J�R�T� �I�k�	�=~�z�3�|�҂yQ�D*+�d�O�$~]0⧫��iN�G
��V��{���Z{0��vH�z��>v��=:�COP'aL��Q��|"Ѣm�s�3yXJ�{Ǔ�ǎ�V�H�h��R�x>�Ԝ�0"�N����QhZ�d�&bp���2�3�f,� �Ț��"x��&�C�(�@�ȏ�?_��؞�!ßZ�Ǘ��9�1���?�|�3 ����9CJO3�HqώJZ�{���gA]]&x.�X������V�S&Â��ҴcJO&����|�?���{��X4�8�H����S��������(��M"�ϋ����86�����*C�-`w�?8Ɯ��6Z�'�9�����TuB��q/+طb��o�"����>�
�l	4�Sf� �]9Xb�8�Qb |�߯C�B��n�c��������)�O������d]�M
	�2�������HjyR<aQ�eO7�w"k9b�tU	5<;FKm9���j�XK�]��8.|aZ�4���0�/��ץ¾���(�b��E`� ���ހ�̖f�����M��KckسACk��e^h�b���o��]~^�H���p1���~���P$/}�h�c�;R����	뿓�<X���1�y�t�O:T;��7C2m����[��	"D�'.V��o��g���X>�Lu�'�2Ϗx���])n�E�<(�#�V�`���v�ڭ�l�z���e��<f�hO�y_B��"(@���.����2��B�'O
�<^�:	�Ii��
x"k���ap�V_�V�?�d�/J������ؐ�e`������yJ�B}RD��KO ��2�7���/,$�$c1U�G�k?��ªc� �=z��uf��`Vƿ=���&-��:���1*i�Qf��xA���[�>m�����Q��.2�G�b�;{�J��W��up�!!G���>�$}$����Q��?P��er��xz�
�*
�f���B�RU=�i��P&8���\��AĐ�_-R7� XփF�m��*S����Y���~�A��)ML����	��`)���ӷ��=��&sfU
6�����Q����f�B)���}�L�#�����F@�щh31��N�]sy_�����_�O�iL��6K��/3�GjI�E��Ij+VLT��`�� ��6e:�3���	<Z��q6 6ė't��L8�L��T�`���f�/Ix�Y���t�7$�M�ԅ ��~GѠ�0��,B(;h���;� 𥧧1ѷ0Wsa�-���7�����d�a���s���O�'�β��K/��P��2�g��ۥ����A���e'���f�m+g���a?5*K,.=~��dC9H���ofc���^ 1@��!��W7�0�����D��Ŝ�ܣ�A���ྒྷ��6 LMB��8¢���T�ۛ��/�2��g�5�eV�̓�ƮX�8��G�A $��!�̴����N�\EL��!�q�� ��6
Z<�-t��L"#���ۨ=ׅk�9� -ti�� ��n�~���KVH��yS�^����^T	�m
������B������z�����K�)!<�;�<Ԇػ�9�$]pc$�����|JX�c9��2A��hc��S�$��S�8������B6�B8�6��|v½���p�瘌H��Z����&�*��9��ۢ(d(��a���j��?�	z�rPL��~̋�.��Pք�]Z{+�Z����
06�QҬr%�\�T�Q-P`��~>�� *GG4�Ԓ)|��<�G����̜�����TZӇ	c_�.�}9L�{��ET�K4fN��`��<�w��Q*�,��oD�6���/k	Lo��yo1�uwR���	�����/p��ɁO��"F�]����RYFB����HMH��1�nA{��%y���B��e��P*�-+�,E��E���/V{�Q��,Q���J��4)k�xͽ��ۖ�J�0=;�zQ��k4�*�
��7�%�K�����F����҆I�.��M<n3�S�������9�>{��ϥ�.�6i�a*��*��Zo77|��.�$*�uw|h�(J�r�`#8a�ܬ�Z�SM�'��}>pQez�K�M��,-O�lx?]��RW�f�1�'��t�p���ҬdO..D�Yt2�����G����߂��_O�K��D0-�p�&MD�\�h�8��(�/U��W�v�M7��\�,³�^�UڟG��2*-]�+��|�;GX��XI�jQ�}��C�ݲ��A!�,Wl�C�#]s�B�*��R��{@]2���%�Z�,�t�k��T;��S�01s����cRF�K��Qr`h�����ة=�L�irW���
�2凶��j�P�|����{	�E0�z*�~����e(��x��;#Hf^
���<�V���b���f)�*/R���R��Q_}&����ْj��T�Jt)�k"�7��]�P�?�cl ����@%Ťj�s�3�8����'
�ݢ�"^8���Ɠ�������5�3�&g;�G��9��������������U+�����ä�IG��^K���g��$� e�P],[�jx���jUC�Q^��-f���$��e��a���=�5�$$��l�yH$�#��4�����l���>��2�>c,��W��5����I�b�f��oґ��9�[���Z�����0���0�k�|��6ô���U�m����
�m����ïO��t��q"���=/
��^�iE�Ho�ܯ�^b:5�h��o�ބ�TJ��鹩�q[<��@���JC�Df�gE{gU�^��+*Y�"h�����8z�� 0x,r��Z?��3Y��L~���Cw������C��O��y!!���R9@���^��Բ(��7JgN�π��-H!>�0�6b�|aC>����}�J8���5�E/��L)6�T��ܱ�����ocR�m��]��?�R�ҥMV�V`s��s �ȿ�
�[�ǯ�6C�>�ޟ���q��@��YL���IF�!�z�9]EHM�W��.��Q�ު�!��
�2)�\�8�%=	��}�����n�l��c���b�lI�5�Ū>}M��¶��M����H8zʞ��-R|T�g�(f��a-�7� ��$�p��ߺm��E)�T�	P�H	lq����t�8Ug"*d3�j)��,jܶ��ɗ�UC�rι���!�_�'��7�s~�P�s�ŋ�4%��x�4H-�w:Jdb�D{�~��uW����c"7_��+�Q���>"��RZ�MCE�q��ɤ&ٺ��1bxKp�G:��М^o������0Ay��!���v���J�%�����*4Y�A��U�6TG�j{�^����/���K�t�3�U��V�8'Ce����%�?��
'6���\�����t2��w9wgO,�ecśi���V� ��HJ	ڠs���£F�B���'l�\S2�'��u���Y;��T�bҗHo*��"�g /��i��Qy�����m'"������1����E��C�vJ�'F�2r���m?)i�S�}�mҼ���XA�7oc��`J��Q�DB�=�ӣ��#t�=�),��q��h��|)L�Tg�J�r�=����ҠH��3{|L�,��Jm���nv�|s�c�+�!��c1_S�_�Ćiz��P��	��i`�ѐ��a���D?�U� �>�����b>1>���_��Дܼ���^	��q%�,%���w�����p��R�AM�4����A�����p���;���r�BL��!>R`'�x�ˀ�#M[F��;h:���Y���8G嬩Lg����W	���H}�T��4��+�����]B�%P��i䂼�(y<0�a`t�VO`h�?�f�?l�7nC$O���fV���@mcьN��$쎏%�Qy"7#�q���4�\���6� �?]�0�&��������OK��쟃��^C�/%4���	����X\T�uB�b�]I��X2"���kOݳK��Q�-��/i�!%M:3��̕�F���zq�,��.Z�c�i�BY5UД��>f�ߐ�M���,�=�8�T.N��Ҷ�&�1ƍ���f����*m�9x%��0�>NW�]L��ˠ>�iiR�����i [��/w��yHV�����3�Q��j��_9u4�I~;CYX��+���X�@�l��J��da��~��|!(Ĉt�Yz�H�m5�"�?��4�W�l��	��dB�������E��~�;|gO���ƺ^�-mv��d4�[#��j�"�r8<B��p)�]@b��G�߬�h|J�"'�'��ӥ���r��p���`9[<?za�g�=�A?6�D�!���7�T��y���(��I�@���Z�l]7L('�₭ת�������W8<�=�X�*O� �{2@�7����H�<��"S\�����Х�-��n3KU�7���v5��_N�\b�\�n�� �YCZm�8X��3ZB��j��x�ى[	�GN�w�cǞ��޶s�J)�?���g�h^*n���ޘ�y��͋%�VpRĚ��Mٳ��p,�vh�u_��i�����Y�:=`V�-�{v!`M���U���y$�}$'�Pr�6T���!ƒx<�X:S�8H :wƴ	;,��6:��ZP��nv������S���L��ԉ�*��U�\7kh�$�!B�������I[z�� 5%m)u����b�ބNƿ{�~:����M\S�{��v�`��������r�;*Ʋ���p�d[<�o1�r������Y�!UޅeK����n�د����9r��nk�<��A��1	ck�e]���@�}h�5p��)�8"��o[\�ғyP�K'�0�P�`���|�e�MC��w�>}{/ff0�ai)��.�3#Q3.�CrIE݃���$�p�q�5�vj��	G�PD�'���'[⠪r5$�.��=�+�]2�<�qm�uƂ�l����&%.Áks���d���4���v�0]��q�C�Iv���y��S~��O7M�=!�������R�v�>�䫱��'ӡ}��ZT������F+۬��{�^�7��Y&�[�8�� �)�Q��e_.xE��F�Ue��rXj���h^��*��}�kqE@�Z�v�!��T�,�-��B�8B{yC��'i����|5�:���r?��p�܎6��͔^7>�Q�4�� i��N�K�`�;�GP��d�
�JG���MX�%� �: o��
��Λ�jWc�ߴ>����SsyH�߽蝅������x1�z}��dK<�׫�SOia��b{���i�<�'�*�ě�s&� @n��%9�;�dc����d:�Z���Xn0�����ˊ0�9ގr��%���0u��ɔ��ᖇ��&n�.��A%n��u�5R���a|RF-Q����*�P�P� M;�/�h�Q�+�����/M�zh3��M�F��K_��N�n�1�59ٿ��٦#S����^yH�t�9�F�Ɏь�A��t��6�L�	?z@%�o~�E��Z\�=��j��4J�@�,�.i��6�R�M�\��<�۵�Xc��E���ݑw��������`]C��S�V�Z-���oN_3�9K�y�jE0�)�Qhm��p:�ʗt�Mu��y���k)�i�0�.���&��;�mHs����P,_��%Xa�V���Bvn�|Y�҂H�DD2�1���'p�EZg���:1��p��~7�U�������3@���
���Ɠ�a�o���j��Sh�D�����VXov�<TrW}b:�+J�h*�j�)�n���ʹ��֑NxeV$�{eܑE��:���D�ɖ[�99h+�'�=���Q�3v2+~����"���P�����RȄ�Qf�\�"�e�����}B���T�wK��t[��1'��t������W7d�8?b�٧O�C�+�%�F��(���7r�\Q�� �9ηr�v�*$�s�D��=�)�\+Z�+�0uXU�	��/��ƤGQ=�x���o��~��ۂ�/ÛH���	U����
+��W�4u1�OCg4�JZΆ<����,U~� �]KWQX� ����6�C�����I�b��*���C���t�Gro�%����AS�ș��7Q>���x�	A��=*�Hge�N�J�jw6�-���pV�n{�`+������� ���KT!���(XK�EP:44IA�w=���t E���U�L�<q%_[�Ӝ�F����O,�S�`�T�gO�Y`]G��6Mrx<���3"��y�'Ѳ�9PD�3<��%�t����<5�u0���=#`�A�;la�	2�q%�-��Y ��0磵�vHn>�{AOJx�"�E��]y͓�!0i�$W�{w�GӖ��+�d��/�i���6�=^��֦y��Bq��������+������:���ӑ�Y��b~�A䜔��.c�c��-�B[����������e_{Yg��G�a�#_�ǎ�i��%������-����ۜYsW<-�����#�P���֭���o!ݦ�+��!y�$�@���b� �ڌ���T.Lά��:Օ U^']����Qf ���,��B�"