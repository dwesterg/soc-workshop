��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bdy��AS7ijm�׼�ă$��*�(��-��)V�+�w�r"�/.�_���50��,�)p[m,j1��(�!� `�$�;	!t��c�e[����<��[�]��	Mg���^��?�?\7b���Ъ"m��A
�L����F�pn�n��3��=�����ҡZ�9��T�a��*[09��9H�곜Q�$����y���߮��R�JT��N��/�5��nH�ߛ���i+�Ήл*���w�2��K��p ��9��h���F\�tˢ��bCE��9m��p�d� )9��J�ЦO��q'��ST�xN�dj��B��I��0����i�dʶ��*��Ԭ�a�c���]��v���r��UI�^R��9��d�?�J]DD�ue�x��9�ý[2� ���6��
9L4�9�OD��4jNlb�n��+%Sp
D��*���:������2CqBYRg����1/_*Bp+J�祮�b������&�������~���:�wv�qZ��2h����7NL��8F�������zɘ6bӱDυ��gR�+���.2��igG����鎱	C�5c�h���&��B��93%�� @z�gÂ��ur��(�w�-�����q��67����@ٸ����I�qM��������G i�y8�r�}����H�B��z
���G�.���S^��ğ'C®��X�G�Q	� }��������S�hg]T��G�#nx�0��v�`�e���VJtY�����V [�Ɛl��'��=(��1�g�k���c��>�b�V��ئpA�u�yua`k�u/X`�0Dq�s�x)%J<6b�ϼ�7�=0.B�=ZC9��\}���9��%B�	M�rv���f�I4,.9�T؉b��vf:���ܘ�PSu�R�G�E�"�+�ǧ��F�r�. g�ӷ^Y�%��M\�*� ���]�z:���'
�et���ב!�����S��ڱ��^�h������KΨ�g2�G��bC���7&
�T/v���V1l �����T�+ىYN���x��Áw2��/
������l��lb ���������	�,\>��q�9��km�~�ɒ�B>�g�d�b=�7��0B�V��uN��L�e�(�<)�Wh1��`�5�Š��Ê���ZC������V����2��<��F̴���G��Yy�{�� I�H@�����h/���%�d�vF�������+���d�{n�0�.,�)3���:�2�]����Zn"4�c>�N@X�$��w�9G��F}L=iݮ����42r��V���qb��0L��*]�K�\�3�1jN�ztK�`���H�������!#�;?�s�L��z�@�5naHc��t�+�!��W�T��#�ϲĻO�4����[�!&��P����G�|��Fw���&
2�bW��3���<L�ko	?.`:bf�����i�\LB�����;� u���"�i9��sY��7sx�$_Rn�b�g;���(L7߀�-v+v�F����ݝ�*F�rJ�:K����0�ntn(�)-�檐E�8�� ��Х�s�,C�����V��m�S���忩챔�b+��v9r7�Q]7zQr%M��J�Reqt#�́�wP�et���ҨRh�i�o�
-z?=��Y�/��2�w>�銤�4�a ��g_U� G_MZ�a 0�����^u�^=��BPB-����lq3�I�u�y�\2�LR�{����$kjݤ�Z]��8��U��н=�l��c���rI*Xmgd/a�߳���� ��c3��s�1�ӕ�8Y�/ք�R8� zQ�b^S�2ճ�/���Z-�H�L䁠T����=J����,t��������M7C����=Ӽl|�zc �^H����Y+uĉ;E �a�M�s��ː�"!kP.��������A�!�S�Ϝ��}њ�^E*޳ߺR��O�U��nw�Y�W���`��m�8��e!���9��(k��)�����vpr#n�mm_k��$�ʢm��
%�wP�|�T��j.&�[*��3�|R��$�.\ڏfm䱖�/xѲN*'�Z�����4��w$���(A�ުqas��~�Y>Ci����pb�����Ѫk�ϻ�B6��'_�A�/�����qc)q�@��	#�G�N�?�l՗!�t��������ɺ���r��G����v~���b~�y���AG�B���BD�W�T� K'�5-"U���l�t8�uQ��g�K���4�/��'�@^���_{O��}8�{���Hѻj��q��,kM��_at����*ڀ6��V+]ٱ\Oe6�22��Ѽ(���C�7^�L�� �/t���\q��0ċ�Y��jD&�S��e�;Yu�K�~ϩQ����R6�u�bB���7Q	��)�[S1$�c������?J5����ͱ?W�nq�Y��u~�ʥ��7�0� 	�%��UE��=��-�j?#���0��I�K0�YREqN�8B�<V�W���d�9A���zuRȃ�����'L���[��:Jx�ܔ)d7�h۾i�����J�7;.X�(���y%���k���ũl�f=ث5�X?n���ןy`��\Q"]�EۼjM�$)��a}Ҽ����������iF�V��X��P9��T�DH�\Y�ǼM���n.���� ���,	�QZB �J� (��w&9iv��֐��϶o��Șz87�
�O9�y;+h�k��n�Aa�� �|��_��I��,�����f�%�r{
�R5%?�9��"�fCn��7(!8�(w�*@L�w�1�/����C��Dk>'�,���ޙ��8�E*�G���Q��A�g���)���U����Ex$10��^_�W�u�/�~"����(4�^��<�C��Z챍 /� b�S����<b��_/�9YW�z���~�f�I}�x�a���0���	�@��*&��脠�y/K!V��.f)�+h��9Q%�.�U_���Rm?��X��x��}q�ïc6�H�)J�5̼+LS����&3���x���*��`�|��^3m,!�� 3�ם�0����y����4=Ie���ξ�+􆐲��Û�����7<?�n���7�i��������<�1o���������Oh~��	X���$_*��3��{�ڽO<2�'d�r�%���8Y��{�T�� Q9��Z��VsP~4����f@_�N��&�sx��L^Qr>�n��E0r�S�����;j�g4���_�(�����rK�WVf�<
�(}��#�N@U��n�����~g|S�-�"������G%��d	P� Wņk���ܘG��46���ꡄ�o	�;c����i��ʾq��_{r�bf�B�)J"�9v-�GF�ˡ��4k��+��s�|�6���'�<�F����g���*(r~��ԥ8#�ɻ�[�����n2nC�:�)��H�v_����cV�B�W7+c�s��O&�gw%�E�
{�"{a8F�F�+�]]*���G�j�F4���PH 	��^�|^�O+�����zf�Q�\q���w֣�l� 򳵅���HR�>ȼ�j�:�ݕ�<�bk4�9�/�&[ �Υ�[br[����Yc�f�q�Ĺ9bt�qB@,O(���ɸ��EG ��-���S�c��<�)�M��40�i��Y�	$��0}MnRR�KP~@�����vf5XQ�,Lʃ]�j!�SiD���A�K �9сU����/�w���L���������'c�[|@�z�>Jn�Z����ι��rd޼	�k�T�	hٱ��;���K���-�CV�00#�q�j���Nѽ�������xB"7�g�%}=��2/T�j8[Y�Xh��=X.�@,:�Q��J�a"����`���:'$��ɫ���^|���ר�շ����&ͼ��oؾg��4]���ByI�u�lF�)n�sC�A6w���k��1;ˏ�uB )��#5B��(_�a��*7��+K�!�AݩQk��c7��	��.L%A+��vJM�0e7�=�L~d��V����ӻ�!��H֖-�M�G��T�sR"�.r�Փ�"L4�dZ^��"��p��'&�%&�@�X*>P�����E�C���Z�&IdP����k�-m�zI�A��� $�a��ʾ�Q#�g�����.� n/�zht�U~E�㽃�[8l�G,�X��X-�%y��Gx�(_��;X��&ك���{��`��e��^�clW�߇�t�2~��s����Mv���H��Db�(�&M�����1���EG�Z�C�wCgDՀ��Ʋa��?j*6���ʯE�<5�4F�,�A�A����yl��[)D����l�^�h�K��ߏ[=9��B��NRQ��.��.���+޽�A
�B�S����`8�ˇ}���+w
c����y���s���\:��EN'�t�?	Ov���)}&m7I5�=
�+�i����#���{�$x��î<��|9¦�`��~_m��(�
����=����J�K&�F"Q�Y��7%��MaF)���=K��̘f��NBQ�s5Ij'�S^qqD�2nL��6Ǹ��t,�>��ÛAH�ۮto��C�{V��y)1)��Փ?�Cd��X�I�����#G�A`B����L��
m\����W[�9��B����\>�
T�3�]v)-���3<���;�l���j���üǗJɷjW�1�^�j=��M��T���x[���T}ӄ��!!�߄��[�&Egуjy'�İּ�>��#�`΀&R�u�,�izPbi����u��˛&؅TW5`�)����
׍�C�p����,'�Ү�MD��Ӂ��ҙr&��|^}`�h��}���S@0�$�Eb���}�<�R��Ģ���R)ur�NK/w�T׀:6e�h�j0�~��*d��GO��;�LZ�U͑��W�Uɔ�~������(M� �MW�L�`mx�68eOl��;q�B�������U?�4^��y.�s#��4\Y�ܛ��9.]~���O���)Fzr�8v�+A�v_>��ȍ��,f��2 �<_�TbX��e��I<7Yd��������>k������O�X����m�ak��xkߕ�y�H�(������:�����0ud ���?�1��=�����I#�Ii�sG:24���c��;�T�N,���+���.P�j�&���(jlCS�w)�h'�f}:�uy
����I�P��I��x��qտw!��ݜ'����{��Hu�f��a��ZU�
B��\����Aѽ
��OX <�Q�b��J?�M�CG��-�O	��	�g2��پ��i%��N��u��xo�9�9�X�GD�����.,�����*e�p�<�-��l�i���}Z�]"t2�CQ��nA[���\ʟ���SR��90	�}
�����/�h������*X�B��:�E�_����HH�C�����ˢ�ύ93@}j�
�s
wM� l�p����q(A(4�/��.� �D��t���La���O�z\R���S�O6����_���J���\��G��I1#)A��)<d`r��o�.����&��~ڋ�o{$����3<G4B������W��N��Rv��ҹ��[��l��͂������@���`�q���a��]�,�.�c�j�A:��#/z�Ju��2�Q�ޙ�U�%���;��������e��Ѯ��m�^(l�k���l�ul�}�Y3����c�I����,Q�����h��W����3�8F�f���A,��g���*�b�U���[w�Ly����J��wk�ʳ��P�m�eٮ�o*���a`���E���.�J`�����r�k|�x�8�n��H�n��� ��hD��
���/:�A<�۫���t@��(IK���j���J3�����A� ��Q��ȴ��BG�L&{�z��d��-���'KBx)3��k�_6`�l�`��r��a�!��B���dӹ����͡�ӆ��ڂw��8Tĕ�(��f	��~9��\B�����Mdh�0��,����V��dEIX ���!��)�#���Е^�lm����\��К��w3O�4@��n���_J��^q\�O;a?��i��_�����'�;���i)ش��;g[͎��w*&�a��F�o�8[�~嵱����@8�#�iC>p-�Mp�`U05�
�5!�q��֣��F��_��2+z��u��U�J�_|֏YO�WpQh�V�N�m�]����3�9]_�{��~L����~=�L���L�(���j�g�-�f��ނ��d�L:�W�L�07q��y�&��ĆZ�?"��Z+��֧���ڙ��V�Q��J�==e�R4��BK's\^
a�9��g�fW�GX�jhzni�sqAm�6_�z8_��2�ی�o�c�Q>�z<}�׿K<�Ζ4S�V�e�O�q������${�+'z��3�C�� -]2�k���1�6�׫~�£���X���� ���Π4kM�9���P7���^P�X�5��^k�8	6@���Db ��֎����&h\|�]�I���1�� ^�g�O����Z�9M�]C�g�8ْ�6j��X�j9� e��_�� �,��E��Wa+~�Nh��e�#7�L$-y��旃*!4ݚ�F%ʮ��Ĩ>��+eyU��*��⟨j)�"�V��R�GtΡ��d��"����� �!%��+M�x;9�[�W?68nX��p)�ᅘ�s�ow/U�6!���j�Z�Sd�=�����c)j�֠0�:1��4E����2�ߓP7&�-�o_�jզr�(��)������F&���9���޵q��&?uL\��P�