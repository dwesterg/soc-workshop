��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��a�gR?{N	[��_ �Q�Ej��W��f����*�'�.Ǧ�5uL�B<
BIO������F`9
B���(&/l��ˬ�B(7h�E��5���	�Nh*��Pwdį�
������gp�-�QXD���p�E�s��[�.-K����i�n�ZM�s�-K�kK�I��^*g�T��:F���I�$�v^*�������3�2uT�J��_b����Z99D��v��	���1Xh���lT!_=�_`,Gz��_������%�m%����s�����Ug��q�/���S*,�#��:�X�R`�k�xT#�]�f�b�%~�A�>[wj�~���<�pZ
1���:��?�$R8m1
�$�@�^�fc��3L�ą��Eɐ�KH�\~�=k~��cu�`0!W/�d�����i!+"��+�K���jn���=	|"cZ{��ր�X(n8.ݩ&$������D��.�k�PՒ���&
��6�ذB����n	������\����9���Nd�������t�nWS凾U�>V�.�+̴�P�/���)p�n�V]ī�9�$m���2�[_��Է	c��͗���W�E}���Wc���w���%�&�k߃�����奒:;eq�[��.��)���b �/�>��K�W�%����d6�z(V:J��W�,u�)r��"�!�
�̹�mu!�ˌ �Z5Q뎣l���'�(��Wl�k�M�3���z;����CXEW^�
D��L7����̌{�w��5�	�c��`�L���稨L�m��Ң�_�GG��D���>��K�1�-�i({�#��)F1�%Uڐ������@�b����<�(�?B�g�7��	�ԗ�B}��gK%9R�)V�q��k�Pq�wp��EŚ��Ę1�͐^Ъ��͈/�����|ð2�-�6�T+'�d�{�`�@�f�w�.(V{�z���Դ�9[��g<A���?����,e��$��-y?��D��o�g�h0�i�\`mM.fg]�灥�𑟜`E�x݃߅kls���1'6��Ɛ��E�'�Q�8�f��DʭRҩ��mmU�ME'P�h��r���Y �Qe�6n=���3`���Vh��	Sy饵�Rـrl1�����)N�e�4��$ي��Q�&
�'��	c必�Pc�o���f��	N��2O�5ÝDJmk�z�o�(��9�%]�Ws嵉ׄDn���S~8svb	>Ɠ�<ۣa�e>ouޫ�^.��T�FfKUE����!�)>���qgǇ#���>�H0����;_�Ì��V�}��d�`8�KC>�'�ҽ�#l�@�׃-��WP���B^7+X���rc���IS�̳�Ň�5��yT,�ng������[�!A>�U��7�י�Gp�޶sե��s�B8ͩ�>�.�u[	%���^��~��(u4�%^�Q�M!(�"��C't�p'l,W�<�!%��y]ʎ����mE�`�����JPU�LC���{S|�t�����D���؈������:�l}jb������؅ho'�=��Ԅ�Ķ�����Ly�f�I�6�B��ǣu�Zb���J��{��:�T��y.8�f�vb����3?�,ݡ��'|o�8/}mI�ҥ���-�G��5��#g^��5��H��VŦ
8�p�E��F�J�p"��q_����N�P���VD���.��j��z5D-�V�gT����#6m���V�y�����I[�A����\e���������6�2
U�i��F��������gv�C�e��/a���ʘK��1|
��a}�l�K�u�0�����[�,����J[���(�ӏ���{�U��䧒�B���u�
�@�IFE�7� �����D�������Ř*2
�g-SD������J헸�6�յF?=��q����F��M�#<�s�mp��x�X�g��v�!=p��n���a\4���Nl&B�dw��k�Ml���Ok���w�j���#�r���+�Tf���LTky"婵죸hmg(���PQ,ȹW��s7.U:��c�R���o�F�=p#Ў�h��ڤ|j��PY�O�L8.�t�w"A5!\ ��'�k�G�g�^Vu�;�y�WA��3/d�u���@�����zK��~�CbN���4$��dCN�a��:U�%�ܬČۡ��8�E�@n7�]������U�}wD����=q�_���ϕ�����Ǹ��n���k8;���H��d����b�VHL��'���$�E�˃���V8�����ʆ�|�7���2�'3����j@'��&�K5����/P��eP�_ ��u����h�-�"j�
@}�/�UN�L��n5#q�.m���ݟ%���*U�D�@+����39�Uvߏynў$��#e�5���;��M��!��m�
���0Wx���Q*�P�mk���}naQ!��We��y��n�!�\Z��E ng�C�%)'�W�
����t�w_8��5��2�J��y6�Y���8��(�`}�R��k� Sm���d�(md=�-�}��5�Mq�C)�1��(�!�f�2�
�k�^��[�ArT�'����VhM+���W�:��#���^~�q�&�^9G9�X��^ȍ�e��!}�8���x�F�:��C���8�P�u�o\S��Ր�T�����0b��_�m����O$�U�#�C���\��������d�mq��Ǧ��;��I�G�S��������#��̐0D�(�%��w(��}������qp%���i�9��u���K���U��}���X��~��Z���z��泇���~c8��:^-\�i�쫞, ������p������:�/��_6>^�����E�Ϯ�R��2�b~��P<Ʌ��C��6�X��������NF	��v�n��'��y9ʳ3��ޞ
6�(��`�_P��0&�Y�F�qQ�4YG��6�1$���� �Kx- ��I0S���w��9��P�(��=9yWa�����ax0{�g�{�RV�g��8\G�j���z2�ZH4A���X�/L���?$��_�����,�\�_�I���vz��b�i3G��+�6~����c�3�\��%3�q�����TM�^y���?�I�.}"��1�x