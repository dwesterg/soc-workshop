��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<�⚂��	 �G.�S���bA���)Y-�
ѯ��qG;���iO>Tz`f�J G�x�}Mq�G�|�
��$z?�/y_;?=��:����TS2-,�׶+W�>Te��/x�>�U���j�b���0'h�AK�Z49���(D��L�E�4/�OZ�|��/nm�O�v���L��?��D�ȝ�7��O�ܱ�SY�-\�q#����`�S =��&��� �IV�leCFp�g�0��6;��(�wM�j~�0,'�C�Ox�S��;��8�3��pElA9�'�.���0m�8�]� or$X�9UOV��隽P�}��h4��Q��I��Edj��f������8^}��VA����j!��汯Ҭ��y���7{��i��#�*�=Q�p������.QfL&24�.b���@�\��O���� 0d�t��X��I�*?C��-�J�tp�M�wM�#7�s��v�Y��b0�����fLb<q]�hN��O��&O�ԡ!oF�_�&�6$gJ��+m��Y�+XP;j�^<��ڷ�&�?�iXY�偙7�qB��vN��Z!��,�ĊPh�=�|�2Y�\v��~4:�c�����&��~՝�0�4nqޠ�dP-��I���ņ�K�;�6]�Q�1�YL<R� PrhSoG٤=�=�����=��u/����O�qo��'�<�����D.�<��Ҟ�����Ď�/��*������Z�>A��(XQ�[v2�V9	�d�%�ᣳt,:���#-|J=xS‏b�����w*�k����?4N~ �4��� +$՟!A�Hʬ�Xˢ|�B��_�tf熞R�ghK����!�=�p<����K^{v�l�>�<y �W:)k��+����+����\�i��m@�h���A�E���J?q�U[� ]Ԙ>�.����!l=��H5���ڠ��5�^�3�Q��e� �5��NW�1-�Z��T�o�ژT�4H#8�c#;�Bj�G�V㚤;�|�w�6tR���m��;���ύ-hS�I������U`#T櫅~>����ֵVT3|ľ/}�!�n�"��c�K�Do=y&����}Hj�'�Zo<� ���<�&��4�tWFX$%?{�?'���U�x����y�4#yv8�#�Q��*�R2�wb���kc�I�m9��'�A�� DnKT'4���b�?���v\�z�|jH|~�s#�'����wQ��&�b�b��?�b�I6s	�{M�P'ߞ\0Ϩ��v��Eo�͡��7�荌��%1��.��q@�+�=�jb�1Q�Y=� qZ�T�/���r��2�p�y<N1�������<'C���/р�"��X�/ �Ð��Vo���E����!1�&#���ju��3q��n=� 9T��P7�/"�K��3���:�h%M�u�u&m� ����h
"�o�=Y���ؼ.sm�����TsS��5���cZ��m�4�$�K{�i�
����ڶ��"��X��Z-%�����t��#��"�Р}�m����b9�yBO_{����s����|w�Y	Q"��y��M�U'໹���P��20���w�� WY(�m�&`������h�.���y6U���v����!��C����1�%т<�ڧي���ӂE`�D��7���:�P�k+x�:���*<^�%�#0K���?'�D�d���i-�{��:HB�c��@�:��Y��bC�f���%3^ z��٥��G�k�[����e[��V�Y�h����Wx��6�}��܎a��Z}<$6n؋�;pd��9�E�� ��r���N���ZS��ٌGX}{���ˤA��8�L
��7l��[�]�@�����=y܄��'�J&���A7��zl������$e͇�Z�y!Y�[��wI��"]�1_�e-frl՗����V��I��p��Xk�qMԺk�)��J�J��v�L9J���ws�<��8�8!�$�D��o���[-�CV|�uX�Z��ko���R3jqq��|-��u�9��M�P�C�/�\U�TO�n8�X3/����)�?3#$������t�oV��l�i���6%İ��`Yz��#x�5��:=��G��V!���7?�h��̪������}>`��O>��T��A�@��V���(�:�%՛�U�ht0��Yk�sQ,�O[�.�&qD��p]A�u嗼��R�B���8�26�3R\z��c��YDج죂�_�~?HmK&uP
�?���뾅0�p��4��<��Ӣx��C�T�_֖��8^ l,|�h��0ę." EQ�H�gCSO*kur��A�⟀5�8SL�f�0��I��U--�g��u�E׿e��
�3����; �Q0��+Z�Ȋ0+�!���l��\\�7k�\�c��i=��L_�?��t�����1��vL
��Z��
�?�T��D����;'c
�/�Bx=G�C�'Ub:f�!(��f�������Tihgj��j5���_�f?����wD\�	V�=vE����vC� sS C~a-+h�e������۝T��s
3R���Q����{t LJ�8l�h��i��&��\��z�M�\+nbtĢ��Y�%]$��u���������E?�*a�=��
#rO��;���By|6�*]����i�>�gi�"�M��þ�Wt�N!����0���&�V��,����K���~ �<�n�;y1�E�.b��VI;���'��e���"(��cKC>�5<(�Ǜ��5�z<`������� '؉k;[�����3���aCQG]�` �3Rns�]�{H���޶0�3b�__mw�)��ژ,y��V��5��XT
W���}�Ć'G���N3��[z|� 7�x=tT�j<	c�7'���RW?��	�67d�ՂfB�� �jXQ~k����c�q�ؠs/$i|bs�`_�V4�+޷���~����/�p�þ���(J@�x�ڷ�q��^��		^(d��b���N��Ov��x��̜�,�)��6Z��W�**�ߕa��"hF."���� �&c��/���(��:�e��Vg�W�P�r�{M�Q]���3���Z���Y����W7��C����d㔠��Fy]U1�����ǊU��mD�~sJ$)�m*|�X!Jt�<=}�a�ɫ���3e�J��5����D��n������t����9�y��Ε����v�r�ZRqe9�[/Hs�87��j=�'���$�4'�8K#+.������[]��Up��;�;[���禀�r�e�F�U�#�%�1�h������˜�ӫP���Eu>��:Hi�H)S�cab �1�?ɏ�s{U7�buÞ��Y�!�p{7[ǐ��6�T2C��|Q���C�/bP�'��
�H���TK��xs6^�\M���>�TJ:��F�����AZ��\xW](q����4l�*ʠg��$a '�3�CL�����C��l���va������FI���E��n^zJO�e����30��_<4fj|㉈hÉ�#�&�����C���),*�����kލڒU���u'`[�NPd�`��X��� �����j�ݐ&6�=��]��ҕ�߁0�],4k"���0P�!R�z��-1��^�u���=/�� ;���Ŷ�afr=X�c�-�i�H�����4��S�*��=�#7R�Q{ڨb쟺c�LԂ����$S�GS���f��P���6<cnv��i�T��6���4��@�rV�^HjEŰ��65�B8_�/K%��<���l��}�԰�Y�`�a�ٕAΪ.	�]�d���2:��φyL�n��4i���sШB+0~Н)�qD]-�v�g&[+���hV ��*5�y�G�y�-Ez �h�����(��(�@�o3�V�*����{mug�	y&(�A�<˚�:�||w�Y�8��$��G�Q@���YK�^_�@�#�}5��q4�>�M=G[SFDE��'Ӆ�����N�`^׊��6���ohq�G�g��cY�g�#���c��S�Um�EL`ٮ�2I,O�~�1�[� A�to-+�>���
�$���*���P�i0�e#���7q����$b��x5�y��6���d|�Y�� z:�Ν�Ra�#�ٻ���v�q[�~�e%�<.��onO�5��˼�!�	(¶�!Uzc��}�z5�\��wl�Ӵs*��N��^�{"����ī�0�6��3�KL�9{�^N���u<M� xp5q��@��-�V~����FQ��1�����,��Ј��?�3�S0�^"!�[�c��1�%v�w*�NG��uS��٭S��j�;i��w���+�v�9iq�]:Z���lF�R��R�?�ɬ��~�
ȭ��'�h'�i���#�>�%�>&N�g�uU�xu����bt#�Ć��F���ץ��~��9��U����ą�vS.{�8�^�;QSg������02.��N��BR����ɭ+G�"����f�d^6.��L����V�� >=�j"ӻ��!�\0�Uqs�u*�$0	i|��pp���m5H��bu�D9�<�E���0E
�Ϣx�{�b�1�Ǌq%�ОP
2�O�H�7���L?��'��:N��~��+���%[u7�Mo���uȯ7�s< ���SqN�{�.�cV�:B��/W�k�����C�kiΚ�F
��L=��
����m�g��n�_u��%J�M��
X(���l'W"(O-�U�5s��-Qå]�*�	��׻c���#IR[	x%ԭ�/e.����{,�B0%��\[;���x��-�����X8�¾w3�J�g�]�m�r���������ȕyaM��M:�����B��<�;=�!mU�W B�mX�j='���^,�����0^c6����7z�ӆ4��"���*@v��p.��Z���Tؓv���:�no椼�;�ô��Dt��(�Zf�Q^^��08�5�H�y���d�������q��[�@D�Q|�\�+���\-��=��00H:��]�8	�S��eJ#�U�U��K��H��m��jI� �jT�2�p!��nT��3tbM���pp	�~�"�å�?
aϟW��S���r��ޜf�!G���ab0N�!+
�@��S����8�)��3��Ђ�5p�=> ����n�grhZ������M%<�e!P'��Y�;w� ���K73\��C����q��&;-��a�	FH(�)����$1�t��a>�"_����O>�8|?z���j8��S���W��Ã1?����T���|�`�Y�����g R���P�J[�ȋ�MyD����1L�*0�<��#���,3��H~Ip�#��'#3l�HjM�]�0V"��%�ʤS�'���5	79�!���a��Fv�Fm'�38�X�>�1n��xa8�֪���&�ߞ���!�����^���]���9���]�����e��5��4R��2<�M��q�?xoi��?�0k�t��w%~g^��n�` &k��܆�6�Dƞ���q�D�U�<��K1�|�LYma*�ɅcA����m�MR�';M��p�j��m�,��L�^�s�6[�˝���%dP�Y�8�Q2G0;FEd��C�o�.��ط���"<��dի;~*R���zQ���O��,�_QJ��gE��YKY�Uw��?��7�xՠ� d}^�=s�o����mC,��� /|1�����_W=?	�X�Ҹt�u��!K��pœ��Zw<��O��X�1�y�Kcm
#�ع�2��|>�lC���j��7��e��W۪Qf��������"��I�ղ��u��5�;C|��^[I�k����[�ɐ�W�}�-KfG�=�v�k})R{3?!6���O��}���2��m��t6��^M��_�3/}�}XW�s��;�ӧ#���G��f��FS�Tu�,�C�L��TM��,М�4�l6��#!�������p�λ�`f�
K<0�j&CI
�ؖ �@�*��Xț�)��eܹ���?ƚ6�?���<Skl�֠����
��O��6g/�+`SY�ȋ>%)�������2���1�Q����T��n:|����	��x�|3�8;��nIjy�m_(���,%Yd¿�Q�E6���X� �h.��Ҁ��x����D`���jl��zzN���h�a5��9���~g��0�S�V�Z���)�3Іx���H� �W -J���͒m��S�_%���^��:-G�`[d�����8�k��v�����0!\tl��|����J0S7�	b��G=�L�� U�`�履 P��B=OY�cQZ����2��竫�ˠ6����>���\,���Mq�pᙊ6�?�C�#{����As:��~���a����@��}�ә�ơ��=���Q�(|o\�G�����+%.�[�����Iep߉����K��m�&SD��l��{,��V
��Z`��9]��*H��w�)*lCf��ߒ�c��)�BҞT�K�R�!�"b�X�U5�m����xj#W����c��c)!��T�"�>�Ͽ��`��l�40�����h�!T�)]�1Ks���>�X�/�%��l�y�Ꟊ=\�W�UZ��(�BT��~|�-X�2�~�����N���J� E���pp�^�j\�V7�l��^���ɪH
��3W1Ec��"��l�� �K����&VA{5ҥ>p�L��ktɉ�5+O�4��7k'�w��^StӋ�cD�X!�Z���y�֎g�[A�w��.{*/���3�K�����Y[5WfՅ�.��J��#a�Xt����q�Si!�M��d�mЎI�2_�Q���C����E��]?T����~�Z%м���G��DQNh0�S8
�;0�z"��bE<S`.�YyȟQ�Y�A����󂧭|3o�����A(r+�vFx%+�E���P�� ��������z�9����y��J�(	B���6��X�zk6A�|n�{<Uw(b�)0�����8;3�TP'0�X�_��p~��.G��ڽ�7� �}@�?1� $����S]�{�	\�f�t�.�&��dK����S�毎0����:���ur�R�'��x��I��������)�F��E��q���A�$�����7:�/^i�����C����b�Ѓ�?i���w�֊��4I堍5X�XAJ�@��}��6����Jqe�}�r�� ;��5�[ O�6r% ���W�sP��1���_�L}O���k�[Ia�D���8Ny�f�m��Kj+������>���.ژ�#�39M�ك1��T2e�ã^;������QF�m+��Y��T�CR{a3]��1�k&���� XN��ǀ�,�	�3-�}�eX���l�&n���y��r>��1�]��A�L�F�u�[�61���7�Kp��5\�h��^� UCGgHC����x�?�1��;�F(�Z�w�#CF�v�d�8�ֶ��$���6���s�=�C���& �N�TH���#j/�|2��Mn�;:�
��i�D��.C��Jf;FR<0v���5ݺ�^x;�b��*���m��bVF����9;��ÁB��"^.�b�K`Խf}v�vK��=b'!�����N�{�d������K>����Ɍ(y���)��!�W${G%3cO��6�7�&�,�����������T�#���`G
�'X���[�p�DEz�F�|��B���8�:F�q�Ab�G�W� �Yq� �8zC��xڦ�K��e`�#]>��&�>C�g'���������>a����@�q�-�
8�ʳ��y���7��ZϫU!��#��{�&�������^��qy�#+�k�;�n ��綦|HǎR�h�^�����UօXE�ͼwĕ~�u�P��t��ߚ����*m��L�|�pyj0S�
�l��cU?qB[�Ɂ��`�����Gp�L�"٦�+[�E�=��H2�Y�[��l!���i�Xc~�BD�=����ʷĢ	O+�q);�o�`3���۪��d�j�����ƻhC5{:���'QH��y��&�D���O{/�&�$}��%?�Q��5u�!����`�x��=up@��?4���_��R?���z2���L�������DEH��x��`a��ϯv�wj���8��ŕc����m��|��=���d2H1j�`��ze���}8�s�x�%�Y��7����� B����苈��m-MT��x͇�N���mgYOz��\�M:�䎾����| X����D���.�Jg+Z
���[�R�vY渮��e߿[�R&{�J^�!W�`\����[�v�z62/[2��q�As��:�@���c��h�e�g��R~Sճ��?[�9��5؂JȐH��$�^�P�Ԧ�m�r% �9A�.'�Kb�S�ts���h�+$	~�*�` �@�*�󎨅��� ,�����s������7���� ���S�ml�����z�����V����_�1C�;Dm$�u�Ρ[m�UI���{#Pj�R0O#ƌ�d�>Iٽ8|��0�ovYq����$"ՆZєf=�`i`>��'� ~��� !{Pv�B~��-�^�@�g�G�v��<�$��o"�(GI{�虏����#=��$�7��3�2��*2͗�C)�����0Dx� cHlJ�t0W[G�����z����=�\/����1:Bk���|M�5���x��P�Z�����`ȇ����������]>~-94Q�M[q 鮇o�t�vW��艥�9�gm\�/9�-��.Ö�X��I¼�q#��49F�����ů�N����}��;(�j{/]�M �cRK����I�����5��[/��a�:�`��_�Q����I��R�9��cަ0U`� �#��/�ԍp���|h��$��fz׹�@jӳ���/��.��xR����ǯ�5ܩ��ok�]v��7�q����32��`%hŶ�	��#���	���;��eZ�&<2?��C�Z��=�#'P�O6�5���Y^ǮYՌ�^���s?�kC��90Ȥ�YU��V��V���H�ω@�J�X�Y�l9���=�X"�~*C8O\nI���E���]�V��n�����EÙ�D?�)��?�D�k�=�J� �p<%Y���mO�U&H�n<�`��@��9��7��6c9�*��ҩK����,�Z��t?Q��&�4����Y	!t&F�kDtS�i�D��B�#��������N=���kL�����<�}�s���Y ֳ;��r�uc�A�H��[]��n��SO��L��
C�m���5��<gsV�M�,���I�dnӭ��4�vM]�L�ŀ�N�
�r��g �u'$�<��R�ЏC���U��O�+�v���D쥱�5j�C��2���}F�6:P�f+)
�{�"v3�*�2�c�Z_OJX�ԥ�,,06�\����{�iܖ6ܐb͇���I���+�V}��g3��z�q��ӡ�1e>��"�.%�����[qu���楬�}��A:�O��@Í��w�B`������맮s��9֨ _���}X�*u�@	�9�Ɓ���c��>�q��x��?�ߒc�Z�1������JM>a�D3ģ��\����:�}�s� �I;m�\�~�O�b��f���N{�ز)����kR"Rȭ6���"@t��t��@�3:�"z�7s{`�g)�_GE�7�n���5Γ���a"�4���u�0?P�ci]�C͍�T����;::m8�������#|6�[{`�0I�'�n",Z&����9h�/��WP��@-����|K��B���1o�eC��_��h���g~�VP���ut����fE��~���I����g��pݧ�jB��%Tă����W��Y�� 4ղ?j`�	*�'���k��
�Q�@�#]L�K2��x�����1���Au�oן"�����`���)�Ĺ�p�{�@��eS|��J�����l8��=d_]q�H�����lI�u~J���3ѽ\�k6��1nu���kL!�;�����ѽ&�Z�@^����_6�#��u�$����T�H���{�[xn6��g6�l��9F��v��l��%���m��K�cr�* ��� ��[�� t������ _ƶ$b��[}"�ҡT=�}T���9�i���y&U-��uI�keE����9��q� )x.=�7�`b��q�g,Bp�UM|85�jr���~����:1�b��h[/04 tO��a�w��D�]�v�!&Z��
�� ��Fj<�� ��couv?Z�yMr����&�����`� Q�B��B�>{��ܜ��l�mE��Ϧ^�<"��v�N/-�
�zF�fT�߭I�ZH�:cc��`w��n1�ih��q� HN8�s�7��9;&$7>&�!3����o�x����*�;[ZM�w����qQ�~4���	��ɬ��K>�F1�=w�;���E�>�5hC\�l$"%ςNP��S]$�/j�S=֓ʋ]�a�.����v�A37.�pK�2��lӨS�:��j&�D۩�~?���H�(��0�w����GH��Ww�a�:�xO
��� ;jc���}L2 ����Ӏ=�mm�L��NZ�T���|fl�^�9��+^�G����_:��@�C��]*d��@�Y��\�4t��'�?g>\,<b��c�f^��(:�B���8#%��K��k]lb���so��9Y�Wp���� w �hU���o)4���oq�4��Q���Zy쁰��Z��t*���Oč�f���|⣶���o�V,Ϥ@u���z�/e���]����R�0%�C�{�y�������e����� ig+�t��>=�W��Q�*�%�1�NM^�Yݗd��a����gsV"����$��YD�4K&�)S��G���>q��k�)��w��.t+��0Sy�a��u����I�ze�ߗ����XaL�
F O��qL�6�n=��"�lbz�i���%�B��v}mr��.@�>܇E�µ�`[���G��_.F�j�;��q/:������;�(Q�#��O_"4\p��q+��\��\������Z��=Y�}��i��e���Dw"Q�N��	�XL���o�����W���܏&��T{ߕX�ٮ6��R��^\85u�\��prҕ^�)u~�����^�&����`~̉c�ѻ~��V໨�<_��z�ӆ��}�a>$�()^6AzѰb%�Z{얛����9�_>�wR��'��z������!�jnP��n��ť��3с�.�C�*���*LY}4~a.[��&za�Ze�-?7����@���e{Џt[�s�������Q���7��O�?�Մ'��U��S~��hne�>����[�5ft�.�ږ
v�<S��J�(���>�"P)s���43,�Q�#1܂�cԢ��H=�6����`��ɂ�q*��ʅ�`P_'2E�Q��Y?s�g��u^���R�J|�9ho�S1�k)� ��Z</<� e��%���2���=��=q�_햤�To[����|E�@O��{�Y�<���2��i5!�۸(ċoZ��Qe�o��$ω�Z��%�F�
��|C;�����	#��?�p��c5n���ܬNÖ,h�i9����ϭVD�п�U�ܒJr�3û0��'k�9ߟ�
<�V+E�!z0�x\)�L����U-)���e?_e�NA�%��U��`:ݖc�M��X݋B�P�N����ob#� �N9�f6t��(����CF�����ȧ	)k�d�8_�R�V��ra+\∃�P��/7�uZ��q�s��˺�.S�WZ���L���[)/'k��}Ur'�u�i;\0�*M��@Wրu�lλ�l��#�����	%w��P�aL}\�3�[�`�-��c��y�F?�1ٯ_\x�����3ܣrq�M}�G��w����5���$��?&P�^~[��p�㜲B�k#��j�Y]J$h��%�-J3��eL����H��Z��v!��Fև���!��áƅ>��㧣r\@�ϒ������w������vTgV��/���-����b�q!έUz.�!Bz�;�o�[`�m�|�x�S8ê�_ �Í�Q�Ԏ�E�μ9��=�Pn[���Ց�����pΒl�ZD%*�7~�0�¤��5�Vf!�]d��ì�i�0	�� F�R[�^����s^A�" Z#�$��]>�@��d?�p���%E�7�?$63�Q�@Et�-��a��({ߟs�\�y]�(�=�ʚf��ëڗ�8�(�
�b/Z��Sw8��}���?'I���L~>�yM�����������a�vj:�9Ⱦ(��� �n�*c�7� d���vTv�_�01���LJ��n�A�y̓5i��y�m��Ӏ�f��]8'�2n�wUq~;��b�?�qj�_2����[��z�}(1��E�U�&=��|�I-���:�+T�����h ���S���~��f��� r2AN5�|��s�xɈ�D��J=�ia�L�¢��Av֗r���:�
LDmD�DsX�I]��{&���9]�V����+!��;܋�Ͱ�i;n�H��Xa,E�׶��hM��L�]�����9��i�t x���ɢ�dq��/w��䭁��F��%�I
1�����>mY���F��
�����9ef
���C�����V0��8����u���7��
+�a��֤d����r���ka[<p�����_���[}�ˎ�A f4v�e@����o\���r�d��0��ʭlg�O#�Ý�lv����آ4Q,Д� �0�0j���
��SQ�վ�vA�]]Ơ���л�b�;��_�t4Q��n�:���1������o �WF-�ڗ�i�4q�o|����n�ΆD-|�,ui�۔�:7¾ߥ�T>}���z=�Jlv{�K�UG$�PgR��A�߽�h��H���2��z����m�����Ox��;3`�yX�Z�t��1�	
�F���lQ�+���ײ�L\�i9+~=�`�A��Kn#ĵT�1����W*��;q��fN����JF[�pw���� v�pӀf�����w6{/�}\��*���k�����n�KQmČW�{phx�en���r��w�ek �{�D��Y� ���î�K�n�v��g9g����<���� US\�[������%���F�o�\M�%~�Q����*Oe������0��+�M)���{|Q����,�ɵ��	�>Hm�噦Ba��S%Ay�2�X��ˮ��<��R�����F��/�1#{����M�<�>���dWn@[�hW�����kp>��~(�G����8�[����:� ���NہǇ����$�	���ZAޗE6�+jc̽#�������,�n0��V�}�hL(�:��>�BgH+�p�F�
�:9$�j�{%�S,�?IE�0*af�P��'N'��{ ���3�:Ut�'�P}2h�dP��/��N6(�"+,�����v��Գ�/M1��-��+�V,M�6ø�����Z���j�<�^A��RV~|vA�\�
Ѕ��=Hv��<�IQ؇
�I�HVH�o��ldT�9�1B���eq�Ӊ�-�O���38�r�����L�A�+�Ks��Y�fC��S�Ia�+�C̻�\X4�8QH��8R�q%^:�?���gb����Z�
�O����$���`D����i�(
�*a�<~<~7�]N��/�-8�Q�����
	VUb�Z��K25��W�B����Ŧ�ε�X��X�fN-�X{+�{���1an�K�a�ϝ���B�^����ζ��2��;��{�՛�-����T=�A!
(s�����`�.���J�rC8���8���,N�F���}��Đb�i�U�2 6�P%�B���7I0ٿ�s�z�X�����:�ܢ�z4]�����{@��9}��*M��K�$ɏ{�Vr<}1$ 1�y5�+���	ZE� PCu���=Q'�b�+�rM"��挴����9��7�y�1���?�1���jmb\��}���'Px���7�j�m�@��f�� �A�_�5I�FC�|1�V���S���Aw���M>0(�K�⌣���(.� ��%Ps9��!hK2�v���h�;^��a�y=��8��|���T�+���9�>���yբ�D$����`��9�b�q�ں�&�4����]���a���\5��v1g����ݏ�e������1�C	3����x�b�I� ��L�]AxF6��^&�!�T]R�׎ǭ��P���%��BH����,���2�@��NU:���L(�ZP�H8u[�;j�+��Ɗ��x_���*�2�����b�U��
9�l�Tu��vA���
ʍ(\xi�Y��U̪��mX�����rA"���Er03�+5�!�k0���*h�Y�c��,c��c{�j�R-���hs �X����{i%�f�2��5;���v��D��I�?=-΀W���a��~�
|(����;�j|�e�<��Y 3��Zm.B0���!�������6u�����"Fq�����9g��@nˈ��nF�jٿ���*W�?�m��~�jzV��@/I�y8̹bL�z�=)�B�W�*�(r��lt��ʄ���_�2c�bOb
Չf4�b�c�5��k��� �1qT�|�
1�-����-�)j�"��Y��&�+�y���rC�FW��y�������r�12a"ٶ�3��͢uB>�C�:-Y���OY��Y'�N�����s��TП~"�QM��_����W��J���ؘ2n��Rou������N�����>�PO�p��^m��� E����b@���
W~O�K6'Q?Y'���2��  �淈zbnV�2N�����C�)�鯋P{��'D��(Q�nm�]�2?(�˰}�2�	'F�t�'M�ɞ��pq3�h�o�1�����gsM�R�ŝ�+-�����Y�Evیl
u�$��k�ObʶT(Y��e��q��ȹƜ ��f����!��8���O�`UGD�U����;�;��R_��i@��
� �S�+֤t�BM��i�
&&�����B�ŕ�6��%��,�O�.�����t�t��I�ؤ������	�����w���H�XunI�����N)8DO*�+�1��"B-z��i�e��K��O(?/6��p4��M+|�*�R#��EB� ���!p���|T�c}���J!! �.�_C�gB�������XD���/;�4�Nwt$�n�їU���� 5���\!<_�J7ŷ��'��nK���e�
T�IT�֛�fp*�;qY:,ҝO5d���Y"Q^Ad�xr'fX�'�6q���m�hKQQ�|���]�8=��Rơ�T������t@��le�5 (�_���x�*nI?�6��y��^�
T��qb�
l�j�k�Ȕ7P�|q�g{�o_j+ɣ��QӁ�ǒ6Mʷ�g;^���y�7�	�w���摍X� [?��`��
�>�#��ϛ�	_��M���h;�E�u=�w������rF:�^]�vt�űm P�jc�yC��H虐93�a�����<��Y��<��;��
E�S�a�����YX��a�,�}]���tFI@~���f}N��jX ���J�y��U�t����lq�٥��8&��4P��vTkba�����^�!���=6���Ϲ�b(?�9�]�pV`�T�/����V��@��w�P�'y�
.P���ɇ�KC�hZ��FO�n=
�h�d��]�T��B �/z-ݎ,8=���e(���P]5\�D}�-��^S��,:v��+ÞH���q!u��o�������"�|��8�G[�HC�$�oS`�9����������ImEV�����;^�;:���Z��:�L �:lH��b Nį~!�?B��^�d;oͥ���(;�N���=a��ҁ�7ѡ��#SI{�Q�؀@��aq@���B�zEVk��Ν?sN�5�Bc'�h�@��V%6���0�x
	���/�vlG��g;��4��D n��g1���-�ԥUhG���8�[��LM�u�v/��r�=�k���7���*���"heM7ƥ}[@-[��,�"�=��_@��&@��WP{e�~EL�����Du��8OۘEo��b|�}���3^� I�*Cuo�b��fW�t�fu���ȕ2�,���M��!{+nZxHĠ�R�-�����@/���C�K�����P�fW����GE+va�vƆ'7D7[[�!7Yh��J�A/��P2cy���*oz��e��!m×�3�~ˌ-6/�r�1Aڮ�_�����1��!�Q!�w9+Bu�藩�8�&Ki }GT4�\[�O��R�%"�:�|"��@��B����Q��ɏMs��F���j_��9&�]�'r^�~&��i�����$��,ӅC��RV��� ��\�U`����K臒�G#���^>U-�tk 
�A^���gX�iV�ΡӚ�Z��0QM��Q�<���CÙ]���e�y�P�{f"����1�*.&���hߛ��hIx��]#D��g�^��ȯ��'��/aފ'���ξ�\�ZKA�# �U1.8�t∢�o.\ى�t�X�~űs�jRKE	S&�����D������6��5��`vڢ��_^� �,Q;���>w���.�	)���O��ŝ#0z��8�m�#Z�"��IjפH�WIn
cG�[*i�7q��&zÌp��o�^��q���\��p�M&F��IF��� P*�z�����yI�Ͳ*[��!w=ϧ���h^����L`B�������f��ن�G��
'J�����0pݨH��A�;��Vi[���l�unޏ]�A*�7�5wϣ���lBM<(��+�{׼[����:��),mQ��C���vT{D�lb�����}&�L���1r�%w��H���ڻ�����%�O�W(�[�s����\��r�n�_�CI��4�؉*��w�}�O��`?���'㫜��_��BJ\Δ�R��E~�Ow(�u����G�J���1Cr}p)u����E*�-�!��Z��ß��_���}�;��A��f�}}�c�U�(n����Pbf���f��Ы��\>s�<ż[�x���r���i:�.x�?��{�w�iΩ�t�)�znt�@/��C���AvʳT_
���>��iu��������_�礋���c��F�/�vT[�"�ݍza=�bio�X_v-�HX8�H$P���u �\�?�%�l��H���0�R��Lh<����8�AՎ?�q S�t��~�(�MV!���yr�B���?�����49<<�+M
qߙ��̜��0+L ������<�l�Bt��9��*���~���_sr= %��~��ŏ�d��!H�6��s?���P��Ș����R��Bň� ���ԣ�}4zI���1"�ZZy:�����?�g�7��^�V�Kj���D���Ú����;��(�Y�E�1ªc�,P��	�[Cٛ�����6~�PW �����{���)\f��i��cNIx�Ȫ;F��w/;�'���y��
�vS�Ow�n����%8��G���ߧ�jg�J�i�vsI�����q�9��%QA�Ǭ��ҁ���V������ڏ�.'�y��@[";�mm�$c1!�c؅�����}����� l��!��P��=�� ���ܪ���z�o<U3xmf���`-�^��x$�Y]Z��7�H����o$͡�9d�~\�O��'�^ �����8x�V�%�w(GJuE&�qF��\R*��4�p�س�{+43���X.��+��ll�S�Ks[ZB�J�W�y%;�V�O���o�����H�FϠ�W?����M�.��a`��8���|�)�3��X$P~��+��z2ƍ�TYD�	��'ǳ$&a?��L.zH�;�!�*������_��R�M�58�g���k�1ac��<�?r����+I@_��Ҋ�n�7�fyP��v�rK��m��������m�xW0:�f�^F�������R��oy�T����� ��.=�m��P*S�5r>ʶJq�qA��3j6��|�h�$˦���v5ض�}��v<-L�&��kc�|T��N	����=*�P�$>�=:���X$v�d|�Ɯ��?���֤�s��:uHA ��߂7?p��s,[��m��ri��;����\��Vkd�>�s,�&�yBݾ�<�k��Y�M�G�$�u*g����:!{Y�(�Bc-Is��gg���CHn#V��F4��8�f��9'�d畯gf8'�ɤ��^��Jk��-��O�Ƅ7t�`y?T��֓�`+J��o�u�7��u}�Y�&p*|]Y�)ץ�.j�a�M���_|˲㋤��%ȗ�_T�Bmq������9�	��U����RJ�d,��Q�a5�X�8yw�g&~X�k_>����F���w���<�M�����|���bJ��Q�_�r6[E����.֟�f%c�N"ƭ�ƴ�'�G���2����> ���}�g�@�h��`-����%�r�NN@T�`;�M]Ir�&F�$I�~M-j(P�ʴN���g�k8`E'��OA��ح��$;BP���L����a���ռY�=&{ڀ6p�=�W�h��!�����Ss�!�LA�H!��`����ה�/JBJ�X�m���)�u`�[i3�v��|�ĥ8��J�r;
g�;;l[�݀ L�]���๾�L�o-5�UlY ��Wzl�wP�$�M��ٙ���<D�Z� `>��!�pʯ��tjo��S�H���(����ݼ3��3�kx���\ ��ʍ������"��
b�%_�F���a��"��X[+	���|9��gN-�Y{{qMr4e����5?������[-��͐6\9)H}
j�C"����yL'����r[��9������GG�%���w�=���Ĝ���$�x"?X��/��(}� r��	v=��v�,��x�Y��0��h�|R6.��2�ˣӊ.�f���~���~��|�L�	�s�~D��{�fAa�7_�ȿ(�)��w�HG]��1[�y����
0#V:��FR�@?oɎ\c�"	r�p5�)[���H-�}J{�b�_,�_X��?���xQ�	jD����m��_��.!�[D��*	���RK���x��|�>VE&��K���n⍭!gc4A^-T/�0I�B��9�8�E
 Y�έX�S�)��u��c��7;N�R)/�� RD9��G���͖��bI�#���g5��)!t�2#�B����Aa�(�7�e��o���qD�����k6\��"M��"�!�	�x�J\/zl|��}m��j���EN�m,����u`\�K��t�6�{%�^�~tK^%�-�3�Lό���Md^O��G�x}G�rHR��Vx�WË���.�IT.�^��v1a���} �����Ɓ���Ɂ6x�8��������$ջv��x=7��
%�-�PE�1$P倫*v�]d���W��O[��_�m{�>����ÿ_W����f�9�z��;�����E����<_�����yS��*�*�����p�~q���n�^����<��}�D��JEn� 1?���%̵SR	�����4Y��0t$���l�p���J�5|dט^����,)h[�ـ���S���({�S�?�x"���_@lW�,�U�s�x���hr_�wp*2\�@�!8�wPg�ؾ�-����a+�o�L�5���6+lpF�'���Ҵiy��?orZ�a"��=������<ǽ�Y�R�55��j�&*�@d���/(��*�sab@�i���s;�?;��_���a'v_XF��p�5�#cC�0���]( taQ����8m�->툺4
�u��\,�UZûÄ�}�����jY͉�Õ�pke����25���>JHA~1IP�V��>�cM�`�L����I3z%74���$d�����f/��uDx�mj�p�i�����R&����'Ӥ�z�-q7w}-�8C
~��̞���+4G���`-dp�'�ӗ鬨���tʮvt���Ii�����|@!IV�
��(
�\�d���R����.0@��R�n���k$/S$i{�J8ɇ��@�xጹf�c�!y���>�.P74Z�X�Yt��U�]%)H^�m��C�2��� ���Q����N��X*���zD�%���]��ݳr%7�_&���_��o�x����s��@P4%DO�+�3�s�Z\	�L��I�qn��m䌯��a��M��N������!ޱ܁W�ʮ��,IB�񦔐`�Yu��7;�*=��ˢۻ�v�u��ٖ�ISD�����OT�o )�j�(Ŏ�-P����R�B����=g�g���H���N�Vo��i?	��g��V�UIqXY��.+�m��2Xǹ�����lzUhݯH)qb��� �o=�A�ϼ�/J���@��9y�&�Ff�k4�h��*b��W��m�j$���`=����6]�Wd��i�>a���o:����W�fG��A��Y�I���ގ�*r^рȥ��D��b?��!�G�ǂ=������
Ơ��js�8���D�>{�(.7��w��D@�g��(�[Z]�a�=��nS�$6���11@r��`5����!�Q���>��A��&�����7��j~^%��f��'sm�m�u�a���&g�4��3,�
���2)r���h�߳�ݸ�r�xx3lDo�Z���$�|G�����1	A�l����}��j���k�H5���QnK&-��k��Y=����!nX"��F�?u�։P�J���'C��c Ի���4�2��?-b�9�!����&�2�_�-���jˀȾ)͂>���������a� �1������]�t��ƾ�L��c����0�G}:¨�hj@\)&����P='�m�#�:������:�\��@9b� �� ;�t{�C ���E�@,�zо����Y�l���-Ӳ�lPG��Zr�����j�5�J�X�,��tn��n�5*�86�.�A�6����A%���w���P+C����`@o����]|#7&ⵧ,���5��V��!����u�_�Z��/VE<�3c��-Z%귯j`���[EX�V|"7n���Qz�����dV�̰k'��g<��7A�xe����{��̢�;�S���b9T��k��{���#����	!P�����_�/�xT�z�[��>p4���X�(��p'< W��$��q���J�(�-���b����f���$s���Pupr/o�.TzݱDM�b��e��v���掚�(s85'\'��H��s+���a��u��w�M�?ȗ���J{������[M�c�e�2�G�ǰ��~�2�Ų�@�1{Y��Ǎ��&�~ų��y��L�<e���V��2��V�C�t��T���� y����P4��> $g4��ئ�֌��dނ��@�W,T=�.�?c%�4h�E��%o����&GvN��!	nW:�}�J`r�i���aC�.PD&dduY!���A�F-F���X_�)�!���8��	���rS*Ϸ�ek�%���X��8��^ �/�i����	}����@m�BY\���C3CK����j�v 2�>����$;T����H�(��9p�OzO]�����~b"q�f��0=��<� �7�;v*!A"�V���E�0SC�����'���C�1Qn��C�L�2�z���V䈀���Nl�}���[�?f�8#��9NX *#�[=R�&��P̍�k�Md�t��s*�y�l����6�G�'�� +�Zr��i�נ��`mQ8�4_�� c����x6~���Չᨏ�K'��6q�����3"5y�?f�I��`�0�4:�''�^��!�Jsj�p���^�9F��bԋh�����k�U DE
���bԭ4I�A��<|�F�/Xv����Wyl ���DeEf^e� >�S^��$��x0rJ[���f9�.�U7�&8�GY���&-y&���ie���&��x8�7ɤ�I�p�@h�����(M�wQ1�n0��s����M���|���	���͵�?_@<I�o��hN�,��`��Ů�fQ�A�?C�KaK!M����+zl���N�l�wb�SV�x}����U���T~ _~	_B������B�{R���k��"����	�hZ��3���ǉz����G���z��(��.S#�PV�i�b%$�xڹ~�X���@�	,8�}�b�S�f4-�̰�@�5�"�L~��@8�u�	k���^I=!	��J��(">t�O�K�H�.G1jٯJ�w<q�/$[�Sf<�+���Á������4,�QyU6��z�fzR�5-�=*��|������;�hE�	��B'u[��S�����u��Q*�;*��@���A*q�1iOp��$��|�r�	��"|�d�3�K�,�4N����>]�I�(����TmD`eo�E�y��b����$ ���A�P���^?;�-��A��Cc��)��F~��3��e�s� �,�~o��9d��6��!�n¡V�	T���8�wx�b���+�_���(�|��w��[�K{�~Ip�J.1�J��eN���ܻ]����4�sm��!g�y�~[1�>�[�-柔*?�`�aƑ�\e[��]�΁ͳ�����$��¬rL����"'/���j�e��0C5������VW�R�8�h���x�ߴ}V�~�h�5�"�"�/>bB.�!���B���W1�������;����SҎ[Ȑw�K��t&��<��a�������o�\���r�c�ngV$���#��6S�h�_�8�nK�R�kI��r^�p=�>�C=3����#�I�V�U�c�X*���Pd���ƌ�_loN
y5�T�Q���^=G|���
x��/�H�n��cS�������noC@3������>�噖�}�ܿ��w�x�]a��Dp��:��^��%tE)US ����O�:�Q(�c���~:��(t����A��L�uV}Ù���G�s��R~���ژ[�ۼЫ,�OH6K_���n�鸜��4�r6�-�Ĥ���o¹D�
$��Lh\B�!�����P�;y�p���f� L�uJ�Y�M�9�1���s�l,�\��qN,m|U�,��A���~�5��.��표A�k�m����~6`�g,Li��n�{0�mM�\|g1ҩ^6e�Y�,���Dii���J��R]c�g����|�>��)G\A�I"G
$�R�[�P�U����^ݨ�f�e�	K�V��6+	#o	v�s��ؽ��V�pBc�	���p+����N��[ȘH����Z+�D���`����u`�D�#Z��<')Ӏ]���Vf�U�c:Y�~(�a(������%޹�|t>�b��B2�S�F|�i����Q+)�6S�&��Gǜ���:�c�-3��b?ښ�m���Ua��'���y�kZ�	�������[`!�`�,Ұ��3U`����6���}��KM���Ϋ	��w���xKّ�A�Mʫ���JK�C����M��ű��֦NH,Y�1�h/�<���0�ّ��L���6�2c˧ݪa�ׇHi�<s�^�ڇV�H�����0	C�VV���.����3PV�����v���Ron*=�t��G_n�z3_1aNi�s���>�twx5BG�P%���>o��]�v1��4zL�k��%o}̋��Ǧj��J���ڻ �t�A*�?l�q�bv�!%5�1	(6��I)�]H�|�c#Ɲ�U$YnI����f0�����^����LD9�+�|�Ȟc:�$��^��~�K�L���f}�Ag!Yf�p�������X�VW1HM:��R�(�`k�n�^��/o̱���p�ݤ���R�;�GP���;��z��wu*ʭ/��j1�R��q9�K�����/Rϭ���W��p$P}Ԍ����G�l�W惚f3��0��0�7~�W�Ro�r(lvEn���$�8\��9B7���;N�R��w�0������;�S���\�>�� ���Sz�t�� �� ���}��2�7;��Jȓ?���L�M��3Ȳ���z@|�
���z�Q��e����B�X�6rI�-8��q�!ݳ /u#ݰ�J엽�؟ Lnp�-4ؘ�������� 2�,(���
���|�V���y8I��-g1k��^��T�~�� ����b��6�ۡ�$�6������*n�ag$�c����={�%lsߺ❺0V ���F�f@�iu�-D���e�>��ZON���h1:'|Ų5"��]�}�>��[�(�4�-Qm-u��B�;VfZX�� ����Y�Ui��3\�2���J4�5���-�z��5���.��p�^N>O9S����`�ޤrA~���F,�<�k�l�b�{�9ARю]M�Y�Fs�����q��̧�gc��,m��=��c-Fw���� �W��;�� �2%<SG&B���O�b��z�nb\�&L,%����_�Hό��.��WT��ȟ[�;i��c4�G�6��o�l���|ʺ��g?���v7g��.!Ҭ�3��7�$h�Lɐa�{o�*�;��Cxc��Ӵ�W�Xyx�H�݄"��(�y�� i$�~��������Hx3�"��t�r��.b�.��W����#�MVb<x��5/���.���ޢ���|��r�Pw��q�9/XV�Ἥ��)��	���l&�I}J]a�H%���'��;�c� PO�T۲��~6�n*�Z��!'\���?g]���ܺ麖�5���������.���y\A�C@X{�ɉ��b�)x �Ζݮ�<"����w�/Jn%�ǖC�;�?�+��-ӟ_�� ���x�猷6D������ߪǊ�kr����bugwo�#-�sȹ��85�<�s�ɅX{Jʝ���r�e?�"Y��=Km�����Ba�O,�3 8�����.�������{9�^�� ���"�������]��pw1R���ϕꤱ��Nz�Z����Տ�XG`�pnsL	���xb�[d�`�3
d0h��O4�4)h�>E���N��zf���z���o��ٷ0�BnL�-���h�E^�y7^}S��� ��6gċ�P���b���Խ(�P��44"���Tn�5��N��]���%�p����.�f���uq��8���I�_Q�.��x�yp�^x~ِ{ e+
=�/�ŻBu2/�?�D:����%���,D�V�y���R���Fr��Ӈ�-P��X�վ�^��vl��4��tVS���>��8Z��ULAd�V��V��G��Ȝ�������|Oz�\�~���B�1M�!�e���*�&|&7c	?�^�� ����{����I1�b�(�&Bq�;���}mf�%߁���s��n�x�	�x��/W4H��T���	��y��pZ/�K�(������gi@���|�J8��Tƙ��ʝ`sM� ��P��T�T�Xt�Lմ�w)�g���i�O>�Q���v8h� ,��ܩ���!������=̞��2r>-ƌ
.��ح��s�0I�V��)�][�j�����#���� ;�|�4��n��?��F�|�r���Qh��Ds#5�b���T_�<��*����*�6�����+��V�f�P��@K�Nj�pY��[w�һ��mk@O���}��f2��&��(7zxB9?���D���h�6e �~y��)�;b���b5Vӧ��Ze��S�3�_�1��!r/�pO�Ȕ� $��p�N������%FV�W��ǐT���kQt�%�!]1|�u�r���H���k$�]Kی��.Y��h0M�>��	Q��-�����T��֤���B�יx��
U���pRz�.��G���*��s+��g��$��_c��C�I�˰�ex�a{�ka̙C���%�aGi��:���A���.��h��e=ӑ� '@�K73���daPv��TuX���Q�27_J:Ko�"4��I6���;�o�ꗴg�T�1��D�]"E@z��a�6@
��"�w���h����A�2B̯I=���U+\'<��
��^"Q'P�1U�D7�o|�Dm�Me�����9,������Ԃ+E[��ķ��ׅ|�n�i/.�W�}H��)�i.��I�R�1���\�S��5<� -=�Y���G��>��-��Ce�W����GhXU�P�? {-�('��Q�F&���#�I�"��u�Ow
7P���5�'���	��y�w�.籛O� ���� �+��?�\��SF��?�2$�v�6J%�*k!�>\��V�X�% )!UN�(��5��`9̰������x
��?{���])��>Փ��wcU��. <Pϑ�Ԕ�R��v�b�3R��X����C�}�~�P����7���z������ zυ��U�<�+-�����v�q_�_?�L�盔rڥ={��qB��kj�O=�G>��9b�2�-��t�}%#��'b+��_qMr��
5��!� �j.���W��n��w�^E9?E�;B���>&�#��