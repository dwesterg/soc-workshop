��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd`�no8�c�7���'���iy���	�h{9­��礋��eQ`VLq<��E9�<(&�AA�Ͽ��j��A^P(vl�DP����rw����绂^%������ʱ��׫ �J�5#�:k�	�q����Ɩ����D֢��r�(�-�k��B�V+��oy��Oƥ_#���UW��K�Kt�?�Ns��~�$Hvl.�P�s��Q���q�/����~SL��#R�5�-X�^4�^I��u�u��kI�x�(gҖ�4�b��#?����1g�~ǣ\C[��*���FYZ�6	���ƣ!Ԃc��j4�G�Vқyv�����F���fz��r�`LnW7���L���6�)�0f����%���8���f��،99�!v �6��xB/"̗ԨGN�X��a��ŀ����,Iz�կ�V��2%f��s�������ڣ���l&�٠�-Ǭ�9��u8cJ���J.}V�bA�.�f
�;J�[&֓u|j{��]狎�8}�{�[j9��))��q������z]
��6�V��;���du���Y�ez��T�j���Hbn�ʉU|Z��Ll�+?9���ڕ�}����r��ѫ���kӯpN�!Z��f�/"B
&�7?CqF�����Jx,��9hRwq���ּr��{7�ݱ�l;iD �n��0�({@Ye�R�E~�T�޽Z�3c����d0A��#����1�TO�W���~ݟ��ׂ	�;x�O'[�������X2Ѯ��S�6�k����I-���֮l����m�!-��O�
Y����O�UwF|1Eb+�P��ufEEM��l��AΒܸ����[)���s��D	���y���Ă��J8i�@�ұ��ۼ�K� �uBS_l�[$�H~~���ә��s汹�oƞe
�O��x�=�,^я�k����}9*L�����EȮ��c}#ť�-G�k����*��koUxF�h!%w�f�k�]�)����BW�j�>(tT�M�ҳ�\���X|���8 ��2H���>��a��ńFw�9_j���%Ļ8N�x�I�[�|N��&9SQHN� �1�6{�MX�X��%�8;�>awS�E"���nJh]r�a"jY�ǀ �I2��X�f����ń&h�2݂fcNr2̘�0���m��O��Y��Ne�����x}*<q�� ٢��&�Z�Ֆ�t�_�q�Vy�_�Z��|��P;���]��s�q�­^�ɔs�#9\F���-^OR��Ғ�GY�?V��%	����L|Tq��A2���XE?��P�';�<o�d�x,U
+�1��Ϗ���Vٿ�e�	�)W�M4s�,"I[˃L��������ܬ�m�H�_ �`2���*�������Y!LOBFZ��d^�M�o@m
	�p�^BV�3�}���&4ᜅRZY�2J>��.�q4�����}�� -�D��vb��c;�A�pNP�dH��H���>���N�W^�F�W�7	��\�ݽ�@@xf�����~��:Te�vJ��P�eE�:�L����Dm�\�'+�)ra�6B�9�r��>�P��Dz1�<om��P}VG���otl�jC4w�\�uo�k�BD���\Q�b��[�]\��O�}���%�y̫J"�����m�����8\y��mH���NIܥ�
#�43A~֨��ʀ�f�xU��dB�tTg��j>� ����W�r���$���vu%ݤx��:[}�M��z2]od��T po	3��Lz��Jgys�g��Dd4��8�Ўh��S���gO��c,���h+<��g)*Q�.t�{�D u@���"���l�ݭ�OF�ո��oj��{�d��6(�#����B:ۧ��������W ��\���U�K��쏨p�j�nH)�wU�������5+�0��H"O��zjܓ0ý��ɰ��ix����|%�+���\�|w� �T��ՠa?���p��j�K�L�"�f�����ۍP$�1@�*���E��n�g�^x�U���3P��,�hЛ#}6���1>=���bv��5��uKV��a�mHt�{u���^�Z���ެΒ�Ҙ ���_ݴZ��Ǜ6�5���Zb
�F2 �uFY(��,�VX��VR*�\�(��"�1_�D�D��=J:̃�gF���K"pn�5��#r��[JS08�AG���:^�^܋���?��ZJb\�2�oz���L~��ŕ�߃�2���=T&i&e�r���i�MH^G��1����rY4	V	G^��&��7���P���zٷ����n�_)"�3��y�H����l�s<�<�T�ڎ�yH�ȝ}܂�{YF���Mp]�Hɍ��~��aQ��Qch��W��̠�l��t,S��!�=Lj`��.�h�c�B���t�3��uO�������.����^�:"�Ǜ�	D����m�[=�8�`v�k�^iݹ}�u�k:�]��Dg.��%q���O��ѕv]���#wo��ߋ����e~���?mAX���[ec��OM����2��H��z���Q�u��#�!H��0�Z(�nf��$�^g'N>�>��9&��|��NABzr��el�\L�ŗ_��IAy�a�Y
{�M~��гgD���\���4:0/�HQvҚ��bX%r��wn��+�^�Ci����u��*k������thV�����a��T%gjX�~'kj0q� ��}%�Z���ud?#�4��9�5�.iu����J��lO�{Ӵ2�Q/9R��� #ɦ��^��b��>�!Ʀ��*�*�4�{Y:E8�:0Q���+v��q3 �Z���$��tJg���}=�iFg��VA�z'13"G��q=,���/��I|�B��h��)r�ҫ�����Zf�/	�VJ�D��-������&��f�2M`����o��$�gR��㛍��t��0�ն��J ���J�iQ�/�U�]l���`w-]BygO���*�E���(��r,�O��mJ��~A���a�L��d�8O{m��\��: ��M��C�G�zq7]�*�L
�m���ռ3��b�-ٱ��G��x��j/l?hy�Tв���[\U�6��i�����[X6���g�ҷ�댎�0�,]���WZ�C��/�F�hSԌ��Uѯ�Ӻ���Lj,w�ר?$����?sv�[A5��0K�����j���ξ$��4�v���b���m�{A�f! 1kN'�-���g�8�Z�	S��EȽ�F�|&ka\_҆��Jk�-��n�?x�v�{�wյpn\��Fa����2��)H$ /��KT򘻧�{\QX�t�!��.�Y�������٠���z���\l?�q��"]z�ZQfx��Ai	f��2hɇ@�0�5=��?��Lꪟ7��=�!$>��z=����0!e̹KG/Yd����85�t� ʚ�덫e����z
�y��^�(6P4�*rG�-a4����QOV���I����1\U���m��z;�0&D�h�blv��;8j����V@����c��������'�R�"�V�hþ3��S��$c!�F\q��d��z�E'��G�M��c��{h�/z�ΚGHG^�*=Fi�R/S�!�󺹯�v@��$o���9$�����&�7[+{��3Z�ܹ���W2�h���r�p1H��p:��q��C�d���VVyk���w/��&��ǘ`�F|?8Td1�o/�9�:��)�_#[��M0�Q��4S)��(b�i=m'c����޹f:�`������x!�U�?"-P���-h*�U�jd�nɉ���H�`���&��LO�QX2Y�/�Q��O�%��)�`�y��9�Ԓԇ�ʏ6��K+��Fj�f�D����M�[����Lp&�cR�r�'a�p}7-v���G�v�n;eq�o��t�^�X���4e��Z���i\V��kL͞�|�����"�ySZ����{��6������o�A��d���/^}i�u�f�����{��y�]M��M�#{�&�	0���[ F�Js���#��	LJ%=Q�.�^�=ؙ/6�N��	l��d��is���ޮ�
@fW N}e�M�� `�f��n4>`����&猅������K��E%%F�h�l�� �m�s�NS�]rB�`C�/Y�pZ����/�vAC,��QRY������g��&2���
�La� D�h��5�|����P� �-�;��}j���^�>i�"ul,��d�_|P��2af���3�ĖM��hb!G>���V\=��H}+qZ�ѬK�n�B�q�Co�
;I�׫u��0>� ��=)��hݕsþ2��r%'T 5Qo���p�/숟��Ǐ�|HK�V�������Jގm�{NЃ�Ȕ3�Y�\�]W���YW+L���Ɩ��������4���l&�&2��8�w��}��������@&.�����X��0���a�{78g�y�pm�r,�� ��L�D��.�k,�;⬣�R���MZK���=4?��� D0�mʳt�n��n&�"��+��_
v>�*��Rk�S�3&~�o������<�c�\�={�(k�L�ak���|�����(6��b�o�Е��7iӷr��c��--�Z���. f��њ�zR��u^+2�ޑ�1�x+>��t�rg|�"w�)�tkߞYࣃs�����ܼ�Y��Y�(�1Zp����h.���/Y�>,�,i��S�0qq�e$�0p�o����}"��g��F<RPi���}�"������5���=��c�U�z>���j�-�f��w�d���fa6VdF��/T����^�gn�̾��2����k%���@�oG�y�XV*�:� _+�����0��d�S-A��۬�\2��nG��?�����,�&����g��8KX�y�`?FRι�x�����5�<�L/�DJ�g)6��Z�5�G6���z�������a�`��)8��V��#32��DU]
ф�g?.J,�{@�滽Rt�1� �p0�p