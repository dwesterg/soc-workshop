��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd����WD��pBYo�`*xu?�|�xʢM���Tb��G��3#H ��������l�uh�re���&%�ϧ��+e����%6�=u=CJ,�k�v��h�罉8�����2W��X_H�3���<Tq�ﱥz(�8d ��Lr�yt�{���$�^����W���>T�}2ťPog�����ܹ� ���Oȓ��iͷ[Ɍ�����.���s"�į����\#z$@�|!e�jy.�Yj`�,�  u����M��m���7�5o˜��R�s��1�}7��J^�V��.�~a�~�,�u�P�4G_��j�I����ݽ�I5[�K��R���������Q.Х�?·!�O�n��J�"6ӆa�h�گ�T8æ�_C�	DX�Tǐ�iR��5B��ݡ���O}먖�d����a
�wi�E�)fVТ��I���n�]o���P��,�D�k6}1�v��Lj���-���Ǎ"M}�P��
n������5��EK^t���r��}�#��N>���V�a#���l`"���-F����`��uY
�;�=�&;�;��Y�,i*h��/Ϯn�#\ݺÂXy��y�6�৽�����]\MN���+�u=X���
���Ao�d=����B�0L�SuP��w9����l��۫: uI���T �LD�(��K������x�&�ުO�;�8��L�)��<Hd�M'ëw����l���2�{X�0��)Hj��=n�����?}>_��(e��}�e��۔��j�وbj��_Cεܥw
�����i,T�7���(��&�6�*�;̬�[l朰�����Q��K�\�N���*�M�L`o�u�W�dudcO�2.f���������"8�F�Ax�2	n��S9� Y>9?�M���h0=����Cѹ5�C�[��i
NQ��	��ǑҸ����~��,s�x���5���Na���� �Z:�W�H��vPr ^����~fQ�|*Bn_��Gʊ��A�sN}q9>(�t�׼��C�
��bb�[�[%�64�L��h6�]�w��"	1�[��9]���*�������W��a
���dm�G�C]�����ĕ
A;&��pA�1Up>� ��"@t�P|��Y8" ���q�l,CMD�(,��6��b�G��^��o�I��S��ﱃ!�@�8\=M`�����m������yZ�ZL�!���n讘��G��T�T�r��D�ys���6D�1�G9��P<�.U5-�"���|���*H�J��@�w�]kd�_u�+��ܢ���o�&ucְ���h3�-H^dmƝO�������!���C6��P���3#}��B�]����R��^��tT���i�A�f����ĸxW�gOop�#�	�&Y�_��p ��U�����Sl� .���"b�)4�@�i���?v��Y�+�<v��=tl젔�3�'�p
���{�[�����N���MF����������(��7�o�l��u )�Œ�(��T��-��=-�/=���pŕ���e�Q?(�R��䦚�l(�k��M`��Q��U
�Q�� ����u������,jxu}d�
��I�i�����xC{i�q5dYx��5zt���$�_+�(ۭ���x���^���056O�*�'���*r�1,��R�z��I���&�>f�LvD�����ǂ�<�����b+�L｡�f�1m�:��a$jX	c����[�0z�7_�lFR}�mHs4XK OW~(8EL>Se��x������.MA���p���W�u�$����B$�����t��Q��i*�?�b�H-�I�?/��eI����!`����]i"mѩ�R}���
)R�`�*��k�P%�83�H�p�"|v�7�5��olcMV�}��S�P��_#\�^-�㞗v赔�Ȑ	�|V�����u_�+5yzEX���S���s_A�s>��)¢�GZ1NGE�����w�ͦ`�nH��|`=Ɉ~��Y�yo�tJ�[��`���au����U�~����)�&��7�����aE?�:z�c@&9V]��u�c.���/�19OGL�=9��4���8��݈Jйܳ8C}9/RJ��b����������"�>�/3��K�$��݅��"�
�����SL�Mq�˿){�,3�x�Ou?OM�x��j>c���`��p=w!u��I��6�<$����K�u+V_�w�f�������$z �1��*�͋����?���N��=<y/�����_q��E�_=*��0
ޮ��)�U��,'T~)E��g�' I ̜@�a1tqL�6���+��������`Җ�r���*��1˟��æк�M5���=�z�F����c���Kn7��8��C�ɮ����D�E�q!	kM��~m�L�a�Y��ĭሑ�=��0�G�愅5��cY���:�+�k�&eh��a3��|h�v/��sj[�I�����?����&����Y��B���J
!��g��c���}���	�i�N`�Y�Bu� ����&�c�J�ʝq��f2(+�U�,�g�U�%��C��&��Ϝ#���nQ|��v>��O���~��M�����3�A7��8:|���(fP�j��|���=�{�@�a�JD?�3<���	�����u��PĊ�B�T��=�wI�ԙ��Ds��H`�Nח~���(���7�M��[k�3�Z#V;�~|�))�G�D��mf���Y�)�3y����2��[*���vl9�y�1� Wm�RD��0��SfI����{�9��'��>���F�j�@?-�&���/0��p�>^i��e�$\��/����_��arS,��ɭpĉeo��ւ
tըo��cC&��<��|��fv/�>�LH_̣t�����	����RoԣkM��:�d���U��>�� ��>&Z�W�g�0G��3���Д]���Us�y}�]�4����)rc�0�������]38i{e�ðt�̴�Zt��$���Aě3����4�4�V����L#}_�=R��)Z�k����^�	��c��6��^9�jo�ǒ�#�����yQ*b6��o�D����'�<$�`��$ fYڂs.{�[�P5���@~�6<<L���F�e':<Y?�A���w%N}���6]LƧlD�C��(��q6�͏��f�%��|���-�_%(�Ze�����x��*L8R�*%%���~d�%3
b�4*pu����U3�"��4k�2?C|�P|�i�>OR]E�$��>��<�5\n%���i�Lqq���D�����F4��U/�C���>}ZKg ����Q����Q\2����@�!/F�a���i4��P��n��<���C��� c��b8�9�3�����|��]�"4LG߆��qreX�va�7y���T�qvdG�䬦��*1p���L��ZC���W�>�D���cn��vg��ǽas�eD������}���]H�F�\��yZnw�������(�����4+�ĨR�H��@��_�����r<L%�kJO\i�N�k#d�K���.C�1�v7��=OWp�)�O����Q3�ϝt\_Z^껲y�����Hf.?�<����P����i�*iק򸍨:����>Hl���}�V�xf�S�?mf��h�Qb���/��=�*Sjt��2������Sbt��T�_G��ʸ��ͺ�Am�^m��6�q��J��0�U\/R��k�.��/���,��7�EYp&����T1-l��aW�Q\�V�K��G�x�S����O(����F��B�_J�v������,2�74�
Kx�3���	],fY��)�b��[&X�o�%W6�+~�L�͔���!�O���y$��&�Fs�tb�Yy֫�3��T�d�.��N��C�"��
�}уwP���1��C�<ǃʩ?����]�1<{��\���ؿ��a�`pL��x���	�,�s��ۭ��q$�C��mp�Ќ���o��xz���1K�B�m�f�S/�X��<l�	��D�'C���jFsDZV`�F2e�q)���d	���p�6�?�Jď�_«~���Y.�������:�Qh�}����(md�:Q]ę^	������IÅJ`5��
��P����9��M>2�;Y�խ{�q�ڶ
e۵�����˧���x�I)�K|�&�Q�n�DHOZ(.[5#�d:S��3�Du:���.+�� �g8���B�d����\�{Ʒ��1q͢�<�+�:�Q��/��b�����:	��C���c�I�a+q�)�qJ�@�����k۠��8<��T���P#�;����sfm�eX�ؓ��.䞊�S?x�3\Di��Z<lЧ#xB�O6mpH��*�<2��Ey��t�Ph���#�NåG��t���$z�уw��>Jф��_�u����>(�EaN�^�<�g�j	ʶ:����G�/ȼ�HD)���ǰ��pc�-Jp�E/(��@3���f�![�~�J��cl_[��g�Ye��};D	���m��
���L$zE��W=_��@�|��Q��P+{�Z�	��'>I�*_dr]�hG�h̞r"v6��"��b��+�)��	���d� ���DD����S?�-��o܁J�D��+E��_�@P��<q�M8F[��g3� ������ʃ/�ҍ�~��7l]>T�Q`�	\��U,D��fj��XLN���g��*�*2�V���R[l�괚��h+*��vFlOy��v�����H�I�2@�V��qT�YOK��[��ԕ�IɾE-#�([��6�T^�q�H/�Pb�=��:Cm���2��&���J9�m�{��b���e�%�1k�S�#_����7�=��@/['�U�eM?>��s:��'��^���^\���w������5;�i����O�:��5�m9s��%��̞������@�3j;����/��� ۛŰ�Ʉ�D�S�8�d��Wۍ�����9�W�>�tɞ�S��h�Ҷ˩�x������;�\���۶֗�V��c�h�ɩ�X�5���'3�J8`
j�5y�Zۋ��Z�̀\Nv���[􏅜��*��PG*E�����_�����/�r��?M��J��H�(%�G�#��;Ȍ�.S֋j�y��IVsjo� )8�-��z5��$�^#�Ĝ���C�떓R���&�/����6��r1�Q��l�,�9�2T����$-)���K	=��k,����+�/�l[+oxdq �u��x�u`�Y� ?z�}��U8��x3����(>��T��9������xr�LF#o�Ͻ�D+�N�R%�)���[_$y�d�t���ԗ� 5EPQ��ۅ#e��G5�����n�,u�F�$ǂm��S��m����5�
����T;�����W����ت�L!�l�2y={{>U7U��	�}Y�Ƃ�MZ
��-t(7G{�����9��9�0U��_��S����~�*G�]��:2�[��ی���2�_R9��A0����r�`�߬ގ�ۢ��.��`r���my�Q'"�EM����9����-���f�fʐY4�ﶂՇSy��q���A&�x'�Vu�u6k�r:��u�v_�.#����k�]i2m��6X�{\�eM���>�����(WS ��s��m<Bj�<˓�QMe�'Z=�g�0�oQa^��;�U�09F����iw�Ѱ���jPv�5+Z���F���̡���,�߸�&�Vl�!�"~|�?n��dM1ja"8#�k���������9G% �ZӀQ���76�n!o˳���~$bH�5�]Dء��[�?+��N���'��9	�ډ��Oj%ZX͵4=0U_R�c���"�o7K�zC#ڹ���1�E��J��N2�y%{�R'z`tf�$��]�6(�Kn��F.�i��@�y<.�鍩���H�� �O����ͫ�f���R��'^��.\J��	�a	�Ng�c{���A:g���CL'ѥ6��K�q�
�8��AA�ߏ�V��o��L���_���>f*�P\�g=
byD~��]#�����09'vzl��kI���Қ��� �މ�i���Ci_�O�<��'�Z��B�2�7�^��Y���[,���n��y<W�p�s�e.�|c��gD���|Yऴ�L]z�����Qu�`�.ѱ�wb{/��
����$K���/f��e@���S��dv������ي5���lC�b}��NU
��i�}�s���W��\N騑�O>2�Y�aHd��B}K7�>~��3Hskc���o�>\��i�R�'7[���Yh޺��˲��k����
Pl�+��%�ᨈ$a?Ώs��p��������}�j��ؕV�_�aP�Z���?8U���Xy�Q!��h�{��[�De_ԢuKA t�&O#�M1_�lP�l|PS�����I?�uO�3cK練ul�A���ۚ�)�����*G� �3�)��GHlq�7��Wp���㪸��.�r��꯴0)�uշ�����f��E�1n��k�� e�o�]d�٭f:��.�f0 fKt�9����c��Big�y��8�� �����8$@꺬Y ��W����U+��"
���jɞ�ѯ�-O�w���R�n�����-;JW�;[�w*A�E�t,O%�ϔ�s� ���㜉*��g-q�Ɖ$g��zg����K�5�$Y��jz�g���J�	8���txިuymQ�_b�i�U5�n���g��Xю˥��X���^w3�[1��	u�&��{w��Y�{�T%��6?����@t�x��[�k#�e��ՀhI��J�L��n�]j릀��7+l�/v����C��ǁH��<W�)J�*K�l?�w��P�E��K~g��lL�S� ]�K$K�^ba%��OO%z�S��S�c�8��h�)�93}t^�{�d%ts �%��ʲ���=9	9��uR^�b���g��8-W�}���> ̓��{L�i�~�ѓ����Id��}yؙi[0����u"}��w��I��M�]�z��R��:ȿ�&
�{�������� C#D���Xւf?�_خ1���Y�`B���o_�d|�˥�ִH���/Ǵj����_�x�����~E�f��UVd���0U:hV"�@�Il�z��<hs�mkG�	��.|.�L\YP�QMLT�=�-�F,�/M��{>�A4*���ߟQI�?1�l�C��ew�KL�y����6i.D6� ,������ �O ����%���c&{�p4�.2�xW��2��U�2�+3�y�,V��z-a��L�	���x�&+c��;
Fo�g���2Q��a���u!�2۵�{Y:!��]�bE�K��^��W6*�Y�0��ߡ���OF�a��β�:��;�2�C�/��@7�-YZ�uM��f�O�B��cp�F��u���5I�'4$s�^G�����\�"��'��-��-)v����T��g5:Og���g^ۈMdl§�bo^ƅ�bx�J���/K6���u��o���H�>���Hm<Y�xNX��^�O
伯c�rҡ��B�����1���澦�bȀ�C�Vg�D��pXG7�;3���Ap�g���6�#�?S�vJgVgo/ׂ�Z.� 	���gfp�C*9�5�\�Dh��u����Z3������{Cl�����W�\�Q(��� �f/