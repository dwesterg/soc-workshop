��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�#mgv�Z�K���E�ɑ�h���f�̰��o��*����|$�In�	�h
n��[f� B�4�H�b~}aӜ�҃pP�*�]EE/k�������Q����6L���bTb<�R�;����Y'� )=���t��c9d*DB�)��b>D�����)N��0��/\"�)S[h.��j��]{�Sil���	���ś����@ޝ9�I��u�u�m����|$�EJ�ǜ����מ����p���rN�y��T(7�>jR&2���ϯv�!b�<9��)�\�E2#d{�z�l�i��x�F,��J�{�$�#:+��0�-��׽���;�&�n��f���3�c@�r]�3p�7ۛ%�)���G_7�FDZ�|�7��+�a"f���G�WZ_��,Ӯ7�c�On��Q����׼����G�Fn��c{l)N�۰���#���16���A	��z���A#�)�x#X1[E/%&��P��,���ԙ�/�I6���F��b��d�fr����w��}�����8>{F�{�����كw���1���8�~� '�R����t1�p��2�3�5z��Ŕ6�N~���{!����U�̔�j^WC��;c1�1��{���߀�:LZ����7w1RA���:�#~	���r/5	�N�y󍸊g���G��V&z�˧�L�g(&�>X�=��S$j�Y;�̱�{��E�fz�;{�+��7�C	͹��
K�b{#/�=�-;_W��{�I[���$�o
Kn���|o#;�$'�o��kX=i[ͯ�5F�9�B�x��ތ�Ro��}�w8�6ڀ7>���]���1a�����f2r��Io�_�S@U� y���Th�mF=V��Ao��[�Ȃ�*1
,:�^_b�Dv��.)�v��3__"��/Y��o_:m�(|�ĢV^K��f� �8����Wս\���ƣ�CDK&�lE�1��ރ~ �)�K�iv��[g�>�j65��p���D���0���6����Ґ�����q�#�]Y�@!�*��"$��B�7�
�O�&�9/��К�i��B8�=8��Ȥ1dX��� �3e��G9���Z�_�7�&N�_Y19�XO���Ȏ��T��	���A`�H�a>�;<Ǿ���fHk�Hz��/I7#�/j�����D�Pr�2�* 'f�T��T�<,�v\����A6��#�����[Σ�Ѿ�5�����p$-����[�����C�0�	PZ�4:+n���@��M�,k�;$�1N�RlX�^�$�N�&Aх��4xR���3���ͮ��ػ����<X�����	QgnΊ�4�Y�wsb�zw�I��kԵO��㹓��B�	a��� �"Ƕ<�_�w�����G� �Ӡ��A��T�؀5����R���Y�a���b ��������񯼛�`ե}#�(G4=��$���\���
U��9�t��s�OA;A�5]~2�^������(�E�U�`.�� %���q�%��J�̛O)+IP���W.8���l�q�ޅ���c|XQi��
kU_�M�����-L���Oq9�C ��H-yP�ð��QӠNr������L!��.,�wN�.�c�����FK�Q�܏�������{���	�|����#b#�0�%3�X�;24dB��(y������*�R�) ���2ZZ��b�����x�:9����ܔ-Z^��YHu�ܠ�Y/���I�x�Pѓ}WC��d����<YЍ��
�n'skF<�ǦZ�.��1YKO7�2<(毈C�_�R�0q�K�`ύj�-HٞS��7;��7a���W��X��X�9.MV�˯�&#L 0�T�&��o�]��G�����q��}��R�\+	��ZZ�U`d5}vX��� �����{Z�]A�Δ�K���I>^�4��޺�n>y���
Ė���ǈV���3RQȎ
"�Z�"<�����6l�n��׻�m</erS�Z��o�]8��>��X������j�⹟��Ct��3}��<��"|Y�G${H�N�T��CZ%�9H��i��q4��IJ�A��!�K�����b����p隁�.��O5����iS���K�GKF1���A�/�5�&!���X�p8�_��J.��� to%��T��:)P���^��̆&$0��V_��Y�a�0>�)Ԥ3g�u�^dv�����6���Ԯ�탕�k�T�l���<ה]�Fȕ�D7'E�\S��'x�#�� ���F�F��@ycb�f'�i�(�Y_��)�w�������撞�;�X���5K#;	!t��Z���3S�ȁP�����7]2u Va*�J�%� EĹs�@�</M��Jmjtz��J�/�u��v���Uh+�S�1��q�+n�ZC���n��y`�!��4Q��tʙ7°2�`w������Wr���P��g��HY"�q�,�L�-�26�TS��RE0&���IPz�Uۗwf`-yp_�qS��Bv<�l4	��u �A��r*���1��n=6K�E�N��`=rIz?�3���An��;���Q�|��b���a�G���Bz�:�{}牠 ���>H���t�cfɢ��8�c	�L)��hi(�oG����V��ſ��)��N�Ej�o�7g��Ț�Kjb��}a��.w.�[��NA�ց ��
�h{K"ǘ�{���s�m��9��^n� ����A佼�F�6M!��؉:����ln���s~$�I\~�P�V��ج��y�����!v;�1�k���R�I4g5�]�ϵ�[��E��Cx���쵷,�]��?�*�w������)U�
q�$KY'ȼС$=��x�~�����Y��p�++��a������_��Hv�H���_&��M>I���ԩ-��k�@�ܑd��ٸ�s��la~��զL�LcU��������=�ږ�h�Y\�_�������C[I�����A|qR\��@��dLD��*{�5//3��з��KF׈W淖�_��5
-0d�Y������+?N�����ڀFq*��zm�c�D*��/��K�r��HIJ���!���>�cD�}�.)��'B¬�7Nƫ��+�\�����Ԝ��`L��0]��n}����8*�1޸����N��7HJ'b����E�귀�Z`@1� �+]�ٚg��fM�tͿ�iŏ�,�}��x�vbW�nX�Z�h9�I��y���53m�a����VtӾī ��x�K�u���Q3��v�XuZSL��Ď�����.����o��dدj"��7Z|]�G��$�
;V�^�,��:����x��:bWl�X+|8�y�?�)�.8��,�[Q���`���X��͡t�u��hə�y=���yc-���lk�{��k��O����I�O���l�����w���<��Y��l�Iu�D�U��� ��S����ʥrOƮ��U�#�L����ڬĊF~�>�Jth�hLpbha��H�%ـ���u�����e�!,��� 6�/�uʩ���)�۠v�O��c�d����k1j�����1f�����s͚/oZc��u�M#��tܜd��/����Rc��O�@�'r[.�op>�)�Ms3G_E���E�~��'w$��'�ܘ���r����91Oչ�l���Mө%j��D���zi�E���[:��O�h�����/{zƌ���:���>rqm�.�ˢc��C�����Ti�L�嚟%Q���4��Es�3ꝉ��J7�y�dW��KsW����J�F�^(\0Á�ݛ;v@�-�P�z%Ef�����qJ|s]��
�)�I-��B�o�V �
�/�z�B�
���T,�3������>6�3?�|V�;�_�'�[⌐�s��s! ���e� �`�7�^���a�#�Ҟ3u�>p���,��DҨpA:3�Q�8�y�W��cJ�.���)����ݴ1});/�eY�+�m(�-��[�4{>���
�y&"!N~F�e��6Mj+��7��+`�ؔ=ş��L�9�i�ŋ�-6lx\�޵7Xr�޿�����<��[�AC��*�J�*�f[��Ԯ����.����K)f�̇w���������b��&FʫdV��'}��l���
��sA��ygYpJ�wXPF'�\ޣ��6��n��u�����682p
�h�f�cB=@_��w�����$�+�����5A����os���j��#����h	Y��9w���F9���Et���%Qw^�9���MF��|d:�����T��c�Ǔ��Z4:;!+����}-�e�W����A_	U�\�X4�����+/ڇ��T�%�M����!�����cwGF��Z�r�M���7}��Jh��$!���E��>�X,�+�+Z�V3;tHn;����5��jLڐ��D�IW��/Gx:�:���'�̭���
���ۑ�38>
,�4�9���b�T����ōp��{���9��{v
�i:U#G�x*�TGxl�`5���i0�T��K|p�6�XN������s��ʎ����<F�4�^�W�F�)e����]~)�o�$p�NV�!�ȯ�ǜ�׹H� oX=�W���PV"��9O:�l�17h#SVZi�>��;;=@\������}�E?�����-ꈧ1�R;�zL�F7l�2��V&)�'����]9�oȠAuj��4��|D�nk�_鿉��1.���2n�
�)��h,�5u�P7�����
���(03")V�>��d�n���'���eD��Z�K:�����㋵�]�CI����$�Đ�Y�1��E"��m,���z3�9�A�z3ϵ����ۋ'��Gt�,��k5�[< UF��g�۩��3R��f%��kuUG:�����ց�Гg����W�h�ø;��-b��PS<�z�q�Ox]y'hIQ�e���+8�|��\���<�`�I�h�-3��������j��3�kiR�fW�[ɛm:�BT�$t*�,F��I�f�#��`����>��j�5S�D+eVO���H�����2/����[�z������P0&�2��ҍP�3~�H����_+��[��ba2"_zo��s��Z���΃v�S���8�b�Dr,b��H�C���#��f���C�Jb��&���z�Y��.��W�\��3Ee>,��ƹf&������D�_%<��.�	{��I�Jr��PQ��L����X�d0ke/W��lf�::��ڭ�17
�%�#lxQ�/(��z�/J�>+.k�iN�u�N|��A�";��I��!3H�%�����h[��Oت��ǅ�=>��`f����,���"�+�R�<ɋ��G���{
=���v��v`�#�"���n�j��+�\0��ۻ��q ��Om��u��?���MLe�JL^�X;��8�	2n3�H���ȿ��t(k��SGf@��fm��B�_^F?J�F�HLx{��΅�(Uٶ�Č�����:$�bŹ����6���C��y��
��(�(Y mT�lDPx�aiUR1�3^�<����µ�����z@��l`]sK}9�vQj�N�W�K_`P��:]�M�3���*|hn��Ƿ�_]��A�:+n$#� !��L����3 ���I�%F���{�c�#��o�����8���m����̯�"����2F.��OU�L]_����*�����\&B84�ч|�|nʹ����j�7tJ6bnHJ��A_!T��8I>��A_lgZ��*��;j��P�,z�(�s{���N��N �Ϋ�U�;�P�]9ϟc��R!s�e󶷿�z��vS��ޭ.��*�j���"��8oZ������6��h"��LA�U?Y,]V�3�U:�"���0��* f��À��������c�V����.�P��<�%V<���5?��E���%�)��:��w¦R�l���K֙�
�&�d��j��G2$)�3Jv�q�D����Wd�z��lR�-{$��]�;������V�	�:qw@�[H������dQ���s|��wi���/Dr�߫X)���̄��R�w.� ۊ�n�.��|}�SV� S��I7��oK�����O�'�A��.�ndhn��2ۡg]1���p����M/��dh���������=�vx�!�ϣ*t0��X0SpΞ��&������f���� ��.�uK�����$�RX	 lr�_�:V��y�]���&�;fB�����i�p'|�Q��Hj�o ��}_g%�`s��$�"�(fs�.m���|4��RE��M~A��A���r�<g���C��"o>�unO�1<��DFm�`آ�UWE�n��#�����PV�9�m��G���%�Re/5�5�� ���\��(���<΀:ӿ{C�QCi-����lʁ����p�1�4/UTթ*CR��x�� �~����rt����u����]ǘ.h��C�[�6�EMc���±��-6-��N�����J-��gT��Ew���G��x�y���E%��y3�U��D��A}�Q��{E���!ўQt�i��%��R�H�4,<��;Be�By����c�@�ŵ�of_�~��s +�y�Yc��u��vu� ��)"��\�V_-YS sH�߳�e��)N���h��3R몂�Uh��^jn�g�=�3_��1n���ѺÊV�����.�5�	�C��K/��[���2�o0�
 ���I
C�q�Y,h3�>k��	���,����bs��N���(&,�z���|�mt��D�D��Y��q'����<ժ����يy��0G�
��lK�٘w��� ��6��T�8A4���џ�Hf��Z��|��3�Jg)��;�9>xZ��̕��W��������ֽPd�L!8"�
Da���RA.+�֋��BZe�D?�~�a��͖���f�45%�D�$�9JHT����R�<8���TQ�Mv@�(������͒,u����Qc8��Oևү!����ͷ�s`����Ӣ�Dg����ͭ���e��$�R//z�-�(�|��+��$ߓ�'�s:_�J�#ZO&�K���OsE�����i1�/�#m�8U�7^/Ǧ'g&�]���ſQGbK��j�E�as_��e�L�S���kS^m2�y�q�S�9VMW�^��o�#ec.'�hT/Ry����v�-/�֬:B�m$���L��'"M�8��UpR��n��O1]��+��Ba�t���dfN�8Tx;�������Σ���,�M�m==Z�9a/R�:X���\�@7���%4�׈h����0���j��o�x�����$
�O�g㏛g˵Ȩ`9�Qi\��F���)#�oJ�ǧ��;5�����h-����u��������rN��	��_[�_<>�7��\F���L��5h�<�쉺߼�]^��7|2�Ӥu�/���?Dc�z���=z��ݬ���V��،`���h�2Rs��2?>-���?a�s%�����z�I��9Xf�I�}�nJ���g�>&RܑN�b���E��n� �	���v ǳ4�V:0
V�b|���DY؝�����?{Z.|�L7 :�����T�/Մ�O�ԗ�����I1{�F�,ȼ[��_c�)ʱ� ����l�a�� ��Ͽ.������@;�?M��D�b��do�	3�nh:��H��(e��IP|��H�g�"O��"�O�kI%�������Е$��O���Nn����,�n�9#��5�NN�������$1�b�2R4r>�m}��j�*��_�)�ʉ#�%��tw�#�l�٣w���c�t��
�l}D�ڧ<�Ϸ{�
c�6V�5��R�xI8ޢW6Sw���h;ƚ���e+I�8�a'�IP�_��FC��N""a��� U�M���p8�J�i�����gX��*���C<م)n����:���q�4Z4����RYL��:�ﺷ���R�<.�@���\)oV~�T� {�8"���_�Y����V8|����d��u;�2�Qa)�s����l,���G�jus"Ӛ
Y�wcӰ�B�opC������9Ǡ���I�BNa�xͣ9V��������k�70�#o�SQ�?Z�H�� �KH�j��7βt�O�@Ћ���sY��`T����}rb�¨b5�^SǂԶ]
4Bn����qbE�/�wX�^� �F\�ԔQ	�^�Z�c*�	����x���2i6�fK�HaY��k�����S���5:tlٖ����>ô��+�w�xt��Ŷñ����UBAs�
�H,\�#icE� ]�8���a��3�@Z8���0Ю��D�;�H�g����9riD�)tw.�W�ǿ����Z.n$i��I��t$����7�F@&Іb�����G;1�����3�JJӁ{sD��A)�ȉÿ���ڠ/�� 1�n��O=2�2� :!��Ş3���Ӿ�ԗ1�� �A�%�R�|^9�8ߐҏv
����gw>�B�c��&�����ϏR>����q܈�D�����	kfxdܯwS�˚T�,i�)p+��ݿ���������D�I��>���m�
�_	i�{Lb�G_���m#Y�a����]�.)��T!5��[����80'��z�e��#���ޗ�ȥd%spͲ��2�vϠoI�����w�N�Λ�AxJT$�>�ɯ���l��+j�N�s�& sH�X�ϫn�
&��p�bH�F&?5
lP	��riO�g��x�֋�����8|�=�8�Hy�[�m��-��*�<�旣��4�t��H�U��6�\��;��;�/<��c���[��Q�(�Ps�%�\��zQ�	�� �us��USg�$�]�1�~h:yY��>�t�)��th~�T��-k������){�/ۖP�Wi�i�賥�B�Upmja��uߖ��WYz*k�>3.M<F6�����5p���+H)3�EW�#��:]��">޽���u�����D�Tm5;cd��;=�T�Ef��5T:�~�
�"�
�@1R9#���k*8T���m-F��ܱpU�/&�V��إR����y����#�㡌��F�8��E��T\�
u�i��b�;��`���R�x��h�s�ͳa��KJISa,xjsgI:xS��he�UG#'9I��Lh�� ���}�Q�eׇ�f���XE\t�f�:�����FDF���� #tĆ$���!���LT'_�(#��<�x�b��qh�ȴ> �ED�qq
z"��D�����E~<������P)l� VO�rU+����6�h���(0?q|���Ll�
�)h���g�޺�Hm>f>���:���3���I����%[��(z+�rM��w+nS�@����9��r�!ވ}B�R��@�<"��YUk%�k����2aE�m3�}���ZA&�>�!FbĆh�5Ok=�}�KU{it�~3����-�C�H����V}�w����˛�����
w�m�8t�̷%�32ǩ|��?e��W�(��sO\�5Ĕ��{�I���}(`�;)k��k�T�c�J��콨h0t���ö%�:p�1�"��AD5��L��` 0��.u"�� l��`��o�b(N�pgmqWeh ��=H(=2_��)�
�Pq�&ef	����H]ci4�f�`�v��QCv�O%�۞�`��Sg7�*���QNҹe3M��C�93�y��j�B�n����w��,���*���uI�wО���P����������:s�����fEK�;���D0�h��6�Z�cKD���3w���IN"UD�},[H�im�}�(Z�a�$��DT��q�՜m���<��ϳ"2��6�7a �O���� u��T��6kb�� �v��A9�X�/����8UZ�\��&�	�I�˄SMҜOP8���cX��]�JL@T<���ڤ�2�)׹^V/��v�Q(`0�j����o��QH>���,W�%�*����$�u�\����K4�$0g8�^�\�[��_�!����d@���=��2	��!��8L�&�3TH�[�D��t��yf/�2w���T�n��;5�;�YŝPD�	���y5�z�j����a�����"��\�!I%'��AG�N�0���*�V����!�+!��B�s/dei�Ӫ�d���%��;��6�8ZTf���]�C�v�J��$�z!�̤���Z7�����\lC<߬�_�FCX�*��j�[z��V[���]�ϝ����N�ŽT�a�a1�w.s�U�E�{��n��
��R���Љ�qf7ɣYrʝ�����&�t�no<��1ZÁ�j�*�<\�ۍ�u�\s PYD����/M4��`=�Aw[�W���
�L��":��o�@f�2���A1Ntb����Z	�Hܞ�E���;���Wm��b�<E�lh���	��6U��	��ݔ\L���e��0H��xď�2�������
���U�(�6+W�M����D����6��-�G��(�Y��;��I���e��J�����Ӈ��@��ĳ��*�V���/�����*��L����4�6�{2&3���X$�Pl[���]ﯛ���yc(3�$Ӂ�@�ҔoL8�HP��m�J���b�+R.S@ �����Ut�uO_5����씠�Gg�0����<��e�b>�����0�m�т�%J��=
3��q|Ҋ��8\"��v2v�<њ�K4=^`�6߿	�q���o�N_z e
�}��9w�y��D"�@��u�9x�����̖Xy���v2`-I�Z�d����c�.�sn�����C~�����ֿ�J�c�)s�\j�@���y׮�H�߳�^�<�����CqÌ�?�,�� C,9	.E>�{f�ݓ���AzjM�����/ 8��S�Mve!s��T���)��6�x5�A	.�MN��K�HQ)��	����W������:����H�8Ž���줋�J�Fw�#8&^�1�)��$��?���I� >(�i���_�s/Nm2�7�a�\+�����=�zZ��ET�M�?�����0\�K�^	Я;l�}v��"��є}G7�]:dBȵ4�_�!7)�#��������l�#m��\�X�l==�!L	�E�ٰ����W�17XT���N�Q(��Ms�U��(�`�v�CZ��HRX�M�ƾ��EFo�ϩh8���6���P�c��0hZ#��8��s�i��S��1u�+v����@���
�&�DA�q�j7�_"�t��顎���KZ�G�x��-�:���NŜ����UN2l]*�ʆuV9nM�>8,0b�¹Ύ0��ȦG�	���c�P�<�g�|�T�8W�xH�L�g$n�c�Tם2��%�