��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8¢�}E0�Ķ��V@�~y�x�1M.�=���}�g�.(���T�h+x��Y�O�i��(�RZֆ����M�7��c���W����Z�iOn�Yב�����Y�#�kT%�.Q�AD�"q�	��������"���QA��A�k�m��Ԣ����4o0Ҹ�%�I � f/�٨����,%&}}�i5 ܹ��
Έ��n�p�1������;f��|mNQ*��̩`�֎τ�2�F�,���X�^���ڇ��q`���pҤ�F�y��TߕʧԴ�����tz����9��������17�E�&��87���Ҏ�r����@�=�	{���~hßcZ3�n��Cs���eWCn�^���=��R<n�����������o�FY�<�ɕ�`�ԝ��b�I?o�j�Ǫ.<7ɋE���س���xn�Q`YѬR�h6��s�>�������>�s!�Z�F�a�
��D��MV�ƃ�2"cwa��ң-��7��	�P��vp�r����$��I}X�i� ���Y�~������+m���F����Ԏ��z|��/�����{�cSM����v�8������?�J/�\x�(
�0�]h�~�3�g���g$�������ے���|#�Ax����TK��ȿ�RE��*uơ�A��WO:�-��@N�w�V�務�}&�T�ҫM��&�ލ�dw:#E��-$2���>�m6Ct�,o��ظϗ�6�PW��p�H�5��o;����jX
�pS���? ������7���0������<�w�~Gb\r�;㊕�rW���ޭ��r��4�41ͦ8"Q��$1�.�lF���H�Ű)����F`ő�ZBJo�������5K��VlC����q�"rl>z�}��?rU��Dt����)P��\��i`�4�<�<�9�$(����!�}�<����I��]=��纩LaGޓb8�!hZ�&dph���,JѢ�A�7Y^�\�<5����S��+��b�$��ٴ������k-��|�SP[�1!fЧ�4&��ci�h�?�Sv��{N��i��ډ���d�ԩ��J��>�	#�w�,H�*VJ�Ƀ'��V&W�٤��d���n���[��GzۗCF+�j[�x�r����%íuJ�����*�Zo��.T����.��p�B>�b���|H����8�Ws�Y��1J���V33���vu4~}�W�8��\�����O��A+� $1�ڟ0�
��>V7_k�ɼ��m�))��I�����[q	�Wh ��jgv��m�~�k�EM�@%�F��e][�����;�l�3�p�g�q2�;��������{��'k}	1tkd̴.�ƕX���bh$����yD�~@�9����݇��< �%���d�Ak���l6J����5G��S�ڨ�PW���X��3";�M�dN3��bi�sY����J%����O��EQ(�_[��dT+P���C��J��`n�EC����+&��iD 5'��
>/��f��oD��t�'?Q�� \�ڢjS�Kzw�ݸ��8��5{P_�@F�RyW��f��v[�䠫�����g��ќ�,�BzX��`�T�3���`�1�x���ӄ�0�:����l��'���
����_n�p�I���9�f,�k�_� M-\0Ϊ��M}	�g$'�3��@hb!>��&�F����RaI��yj<oQ����#�3�����!��h�rm+Z71�8�g|�tuCiP�/�Oz��[���~�}��L�1�c��\:�����U����5���g_���A�Iq�y�i�č�;e��Qx]e�������\h�Tk��ߡ��`5Nq?� ��
=���FV��~�����W��m��S�R�B�b�An���'�+���[w�)��|�ר�=/م��T�~��iè]��Ld�R7�R1(��4�7a"��l]8S��Q�kq�U	�ߒ
9�WJ�_ y�ۑ�?*��
<Pl:IVoަ#�D>��Ek�)c�ӥu��&�5�'��������t���	�ʘ�xQ䐈?��#Ag���W���*�=*؏�q+<�YD�t��E@1�o
2˟)�r��z� ���O�\�	s`{	e�dܴ����K�3a����+
dས���*�Wȸ�S)ҳ.�/�!�c�mi��ɯK�OR���W�l�"\��1Y��Y:�<2��EQ}�X�ͪβ����� i{+��֏&�t䔲Ҩď�	����2�/��Ŭ����W�v��3&��k	]�##h�[x���L�������:������H�e�9B)Q���"2���o���%��K���ʋ$�͜l>�:6��K7f�(d��5�hd����G�h���T��� D�1D�OF�����os�/`& �ӻ
Y��~�����e��^��LT�w����=�:�BZ��c��LD����<���o��
3����J�#r�����=i�Sg�8�Ю��/�Q#p#��� �8YlT*ץ�����6sw��Z��E���mm��@���;Oa�w���=A��VRR�JH-68�!&����(V,H���@���8CLE�j�|0tnң�H���C��k�����K.�(�W!Vn)�:�����(��h0�f���>��a6�^IW*$��n|��C�T6юy�N�J���:��䣪!�[ ��Y'aI͍�/��~j��}p@�U�/:�ĿЍYH֫�:Y#@E�	���la ���2��[2�"\{����)
�+��+~��S�Θ�-�Ѓ9����@�u���kgO��B�pqNW�sƺ�1��+0�~m�����ƂDL5���Y�{ϲ��p���GDM5l�(����ȕ��1�G�{h�&h� G��:�v�z����=,|Y�L�: *;���^�����^�z��J&~H�Xd�w��$�C	x�6 �7��xMؓ?H�&H>9�	p�T�v�>GY�i3H�Cg-���d�iگ��^n��4�	{���I	�S�TI}�6�L-^�I+�:/xS��q}/I9xڿ�����E�7��?���t�j.?$�&�p�W��e��f��Y�=�ɮ������3FWV�^��c��]c�@�&���َ����,\V�\1:�����h��d��-JXFs�+�;Ϡ�G����Ly�3G��i;���@�cqΆ��Z��JȴP���u������.�ai��&�+�z���$���<�Ăj8�Xc�a�/����05:�F-i%s*����C��rϺ����$7P?l���/a��0�N�Y���ླྀ��*YoV�^����W��	��\�1[�����n�u+��"[Ŏ,�AVH�F��	C���Y��+�5�
�C�K�-9,]��R�؎Ի ->�.CN�p���p�߻p-8"��kpv���1]�7�� �����ӥ�HR	{�y(j�[�ֺs�̊����K�͉̒O۫�%���q,�NC^�H�_l3�X����P>_������P֍�0�Bx��~X�|蝅ZT����;vAh��_�ڜar#{� ��ϑ�Z�II$V��3��RZG��yQRa<����Wr��;�[�+h�"N�=��
��P�~�T ���9t[�%� >��H�J��B���S�gKd�>oא�jO5�e/ѣ*Nh|$3^�l��cR�-.�`�Za	�(=�8t��F�蓥�B��!� s�6�� HTSՈY����l���!�4
;o��4"�vQ(Ș�n�?2{�;�b�hD).����^3�8˵F�m��ؕY�1�36r�ݧi!�1�p �M1� R����Z��yP��	�\�3�2M��0����GA��UN��d٫5�z�*9��-�R�HR��Y�����a�UW1V�ō�����j8�R��ݮV�b�G�oM��6�;�ew�E&X���,`
D�=��1�0���Yu�T�`��Ty���u� �.����Ct{U��m\'<�ɵ�eO�mm!��IY��Sh,ҌҸ�a�ao�^R�u���Ӻ��ޱ���mA_�~E�"����By9��S��ho���(�#rI�������^a�S�%&)��w��Z��^�4�>8�,Fo��(߃O��}MQ�4�a�-��NJ�=hn����5W�E�� w�c{�9��A�4W�l+a�ͺ"��|�����:�B您����8YHz������x��v\�ݞ_J��4|���+��Uz��PQ^���Z��E�O�ׇ��Ӭw\�nwg/|X�bf�$���`3�y=�7�a.�B�م��H�)�RLurQ	b�.��Ԛd@�1m�a���(m��>�m�n7M�É�~����|V9��&��� �r]L8tm��JAs0�a����9sy�3�￫�/�r]����Hn{�ݜ�0��KD��ţ�-.M��,9���bD0h[��i�!&ы�Yd�Z�!>ňF	_����V��ʚ{�Hu��z5:�I�P�â�ÄU8y�M��]|͒KfZ�<�����rGRP�m��[��g#�s�1��yǃq�n`\!��f��� �g۬�_��G@����B~��{EZ����H����<��pkh��ӡ�W��$�����P�WqV�w4K�_��Y��6�T!(��t�n�"���ӓ5b��T�e�}M4����fp%��)��g��-p��7�cdr��Q�xϚ��e�fL��B��(�����C�My��KIi���'s�O��Yv����p�c�n��6&JW��dN$�&�V\�A���4/ZI���{��|Tz�,���j���4U�ט·VOó�<Ӕe����V�>��.!?�#lHyŃ������$0ѵQ��4O`p��5E�����&Wƃ�rp��y��Tb����!����4^2ұH��i���|^|A<F�m���;i�Ee� �)��y����qS���nr�����f�����\ں,9�qS��\�z�ӛ��OVl͞�$�h��
��<��=�<��|�5<$�&�/b�;Z�2��zM~ud�m�K��P{Uo��)T5 ���y�ǥ��CY����>���� N]B${"�2���Mђ���Ԟ@���B?�X�y@���=��AmZN0bwD�����<��~�L�`�?j�3	C�=��Μ)����fhG�V����_u���-L4WT���>���o����Y}i�#S�4���r_��cߢ�~=G���^[��;�Eߧ�����X�/R�iv�~��	�4��@�2)�~�L��(�����{��ڼ�g�l���ԭ=Ny�!`p��;�ҙ�R�%�*��xC�+�Οa1�*���K��
��~�0�;�&�i��l�Vl�"��k���"���7��b	)���@�I���fE��1y����s���\l;�<54+��C�t���r$�.$�/�8�ZNhh��s�[���]��P7 O�8�s�$P���t㚈t��[_c�E]Jd���}״�$������S_�/�RI��6����Aoפ�&W�Ԅ"�D�yA�Ue7�:�>�W��	�����NCbo�L�I���Ѥ޾թ=������08���¨�����O��H@\H����~.����`h���,i���q�.��0���M hc2|�R�$Qu�KXG �܀󾛸2��!h���T�B:�j�>h�Y��:�8��m9i#3��\����1�c��$�tH�"��;��SsZ�ި�'?����An$��(����	��`��t��\09#eE��Dn���š�FX"0�k�ڞI:&S��:P�_�~�X��?�a��̭�|�F��2�ͣ52_Ol��:ˍ�Ruz|u�闦d����`�&�Ф��S��Ŭ��`��@ƽ<(}���x)n[��go�i:��Om0{.�v�@���>ANe�)Ⱦ��<]j�Z8����N���N)E|o����6�Ŋ?:i���,d84h��6��jg��`@��z����5K���;`]��-;٫6����Ul��7���Ѡ�c��Yha��.T�g��Z�>6���th��|���_l��g��!ؚ,k�^f��hǟ���0�rӋ~_�e�l5d�R�	̔��T����q*r����q0�ŮqR����$���N���ix^F�URq4�r��]/�����h�4�Hu
�H- �5�y	��������������Y��G�z2��s}}�;)�$��d%�Y�B
�{8��w�5��25�Â�ۘ����»�eD�aN�Q`�[�$�~\�I�s���`*sZ�i��?I�Ő��7⽏��{����-?	5�uA� Lϓ�c�~b��j�
QE���~��
6�8v�E��XYe���zr�
��5����F;�}EB܉��܊�#�j������P��'�T���>0�>rZG&6S})�M�/��1Zɠ>a9)As <l�#�5��$�*z>#���v�D�����as�O�(�(�h����,��Ҥ��
*�����[�%E7�x��u(�m�%� +�LL�gҁ���U%�e�-�-��5y�+y=8n@Ld��D��j���-�F��=��� �	�� m&�q-k�W|�`��+`����F"K	�c]>0	�bz؄B��Ho���\�5��"E�hB��#��+��s҆~|W��B�+s�}�P��=-���ϲs'��^4��.f�}��4vo]����?�-h�k���La�������uGi������wu0���~�|S�1CM�hV�����p�Ҫl)�t.S�a���J.�F�r>'�G���;�ƧCA�HBW�E �gޜ<�.@w�$r��\���/����j����q'ٲDܮ����*9k.	��^���jy~C(hLGg��*���A���#!o~PV���/=���\��|�!i����gu賂@���Ay����ч�@��?�Ea1 �����Y����KB�M���ہb1�5�Gn����ޞݝ>��PNj�H��lp /*�)�q�A�&�h$U(��=�n.%z���(H�R?���Z�Q��H�C@Jg��<K���jl��1��7�Çۢ�<(s�Y'���3΍����G"�J�3JS�=��^V�����y�8�bD6�[\ߕS*��Q����+O���"����Pt�`�����Tʏkz��qmo�;��<]F1�B<td �l�/WJ^)� �����螅�	�]m��GQ���u"ƾHql�8N{�b�Y/�J{)�TR��4������RǪ��I�o��ot_�.� ��Qr�����ߍ}�~��'- i'�k36����J�1���,Ȭ�%ǿ��&��<����J�i�����*�XcKj�b l���!,Ra�ѓ�g�*y�ŷ��[t��c��W������P%_�)�'z�����٣���7�Y��jK2_�oJ�V�M�^e�6�t#�:g�?T���X� �(��J�z�ɀ�w�jld���Bj6sv?1�^�E;��Ujy͂cl���=����5�� ���a�6�8�0��$�{񨓥�*��ä��0�d�q�kE�a� )��l���xkn�@X�:��k��!  {�nK����KH�ne�	sT٥��u|sj�xˮ������=�iR
�Y�"M�'>���ǹ�<��\)��� p?:�F$�3G�d�}���}ſ_���1��[vJ��i)vpx����eu���QjD�͗pD�:��JTxxU�P=�}�S��~/�b�/�ɏE#&�y�i�Nd�<+*Ů�eߤ�\�^��Ƶ�ĥ�v|�7 bFDq�3��zEV��{D>��B<!,�>y3F��1/������#��L�I��а��+�/7�۴&{���J�X���J�&�qMȌ��|��m�.�Js����~�~g�F�;�'�z�h�)����p�:dZL~M�=z�X�؃Lga������q5�{�����f�|n6%�i����K>�G!J����벦��B���15�]�S�(R[aɔ�T\3�S���(tő�i��3#��ߘ���}���.��Zz��B�"�C�\fW�A��}XAaa�
�Sz��[� �5�aq�*h��9GG��/�\�#��Y̦'	�<e��1+�T��"�6S�Sq��+Ѥ��ڭ�ӲF��??�0�Iͭ�=Ho'����2.E���&C�`�{�k��sDY�L%K��Jų��	�^�d/'���doܖ���hyV,_����X'�5�u�w!������Cù�H��F�D�@H�ՏL�+U��WІ��ExL(�]�w��M��w �c�5O�kf�~H~	I�@�]I����@r��<�i�˲siϚ�!4hP�\�Ԣ�NY����i�] ��l�yf�Qe���G*�Y��e0��ׁ��W�Tbe)���g��{[�R�"�{z+��܆�`�qNR�P�ok���e>�����bHWQ�P,�b�fѠF�_��ܜ����Ɔ�v��e��UD�yOߘ��4�ND�qq	/��u{�*;K^n��N`@�h��$3���'���m��݅/w{xl^DƖ`
�$V{a5�������H��&g1�^_d��idU�;��sګƛ��J<9SK{�J:'_�Q��ͽA�!2�垑+����4��Y��+2:Uk�~�fY]�L;��ko���e7i��1�S�� � ��҅�?�Wv��i����N��b�ې!�����d\$i�s�I�����xYޑ�����E��/�D�nK��ڟ���-p-�Wm�p-�*n��Ro�ܱ},Z���<��\j��L��x�U J�5[��d����Y�&ڎy7���
���
���y�`�gM.��Ү�h*�AV���I������� �[A�ĩ�u��?*	�A�z�[�\�Q��B0��������:═���TdJ���q����GoZ5��I�ծ��ä��������4~��IF����Ix ΔaA�*6�9�:mշ�M���'X�n�jXp��S���uQY�;�ɠa��cC��cI����r���S6���qə��;4�&��^u��L��R�
+g����&�@`��<l�z :�w7�B�o���E�4�* YELᰗ�ϖ�m�^ц��s��V���n-AS)ڍ2�i]����	߶�(Wҡ�
x�.���*�.J2���K磱�p,�"�Y�T-	�6'�c��iޫ���]ئ4a�'�G��옑?�ʸ���z�|��|sx-�'����*^�02� H�]6Q {�kTV�����<���R\��D�g�,��^5��I �������4���P�Ϳ)���#��.��4*Y�w�B��������jyZ1�%�����%y�ڐP��������~V�a�$�I#���
����ݔ�<Ze7�z�9���*��4s�2K!���D��5T*'I��iRl��J���_����!��jI�f��6aɦd,-o�YE����4��ǚ�n��s��yz���lm�*!b����q�sz{� ПP��eY�A���roѫ�����ñ�����?U:4��8��� 1��u(�Hk��ub��@���fr�|I�Hs���O��0���y�3����F�xkXs�����
�jm�~[h�7��{8�i_��;-�s�=�І���,�)MH�����<p�����cWXn9,3��($�_�#~<jRȬ$��J���/�y���-��<ڑ������@���d������Iqj-���e�a��&�D�$�߂|��9�]�ج`�D;�_2�\����!/� Y��m���|u�C���okO4�������4F#�CD��Atc<�����EK�p�q$�J%i���,�W	9킣@]�9�TQι�@�GL��c��Q@�\\��^��¥g�r,�$C�L'�W��ɇ���7z&�Q��?�@Ҹ�'4ٺ���0��3F~��8�L�����Cq���q�� L�6���2�ڬ[޸�߃'^o�������H�>��*�/����ynr�tE�]���-==9~�wS��E~Z#��O�ζ��/�[�梳�Y͵�Q7�8����:Q�VDC�uWI>"XG�� ʊ��Z�N��Q�M�į2��9�mJ�+�!�0#����$w��$������YU�NO����*��H>x!t�&C^��B��&�s�خ1�NÝL��)�/c���018�3y���X-0���?7���]���hM�E2�r���	�
�^��$��FLi����p
��f
�����쩼\��xoB(������`ރ ��t}c*�_������$.8`}�O�9�>�ہbW4%�l�k�=`a��ˮ)��:�~+�UU��!?��Z7d��ݗ�,x�"9��*D�&;��N�u���]���D��'^�	����b׸ؑ�+ͮV�k�R���(f-�SѬхq�SA��AWd�y7>�ʟŔ?_��6�����v�������%Z���'�+=��>A�%j2�y���� �*�ܽ�	m3*Zu�T𦒦j���f�E�{fm��)Ϛ��Z�v��"�3mSҺ�GJT�H��U�i��475�dzxw��L7�*�iΊ(��Wۃ��z���es2uoJ���P�����Ωw����b ;A ��J�Wl`����]����F�.�-(��ߢa����A����.e?i����l�J�`�m�ַh�']\�%Q�wf*�ղ�) �;�ݝ�����J��6�te�W+9��w��Ճ���C��P�J&���Af�OMu�0���|�0=d�`0f�I�xV�ϊ�ߝ�XS���Ԫ����a���ߖ�GQ�cb�	����|ZW��Qд�5��ݳG�������ly���3���U��L��BZ�I��kK�$<��w���t�+H�|�K��J3�9�{���o���ǀo�ۺ*a���o�^�	��Lj���[�8&vS�_����?A��d�ĸ�8��y$S�ӷs�9�꫇eB%}Z�>��-\*B3�kN�qITI�j����e�>�G�(P<&	��E��������;�v�]��w��SЪv�ٴ�~A�F�{N��a�����v_����n�N,�/B�1��.t\"���aX�)Nd�>s�b] ���t��'j:��������%�B�>�.�AG~��CP���c!������$�A�kw(FjK e�2�n�o��BP�wΎѵ�܏9���y��XCr�ð�.��Y0LiW�>��|^g=ρ"Mȩ`���'��P������k�?!���C?E�6v7��Jn��u��`jX9��Y�?Ę�q%$�@�V�[UT���\\Uk����ޟ�CI���Kj�a����kW�⨽��'y��JN���E�k��`�wй
m��P�v�>�;_��E��h��L�=C�����ҽ���O�<c.��4[�ȹ�)X�;f�x�읖YRtׁ;�OC�R�O��!� �2T(�t�ס���e P������*�?��c�ܗ�ܫh����0���V���6�)�kB�d��S8�kzɼ���\M��C��-Y�U�*��|���G���=��m����M��'	&���4�u��� X��������l�W?n.P�Ñs�>�Y����8ϛlF��¨�=T�m�R8z��f>�;�4=a���(��<^
��Iط�0��~��]2�����0����m�����U*�ζL����-�������S'q�AG���Z.�[��I	���͍*R�����lk�sOu��["�t���h��9.�@����DM�G��������HfZ�м�>/��6+�	 5 H�T�����8,���|_Č�O�A�r��s�=�|���Q�d��O7P�+�ת�ѡT`��M�)R&؀ �om}';�GH��xn5+o�v�|��z�sa�A�k��+��5�"\��6����H)�<ZO� /K�`z��������fB6�
t�i�I�h�WGj����f&|��Su�� ��c�'�e��%��ͯ��q��k-�OV���k�þ��q����>IĤ�?Nm�Y���?�)�����D,r����v�i�
��
�@���Q���ez`z[._&	B�@(�-xrD]�nm˛�E�@�$<���lذ'�KCQ��ϣg<�g�j������Z�x�s����4�=���������>����x�WW(wPu�(�.��{�*r<�_�~;>��;�p���My�F�7�r~EI�	��&|�����"�)���T��%�'���c�%(��?5X��p��cR��u����I+���?r��l"��T��A��#��=�@�%�>:C�o�۸\�S�G	����
���Ʀ	��m��&My�|[�K������jv�P�{�?���!�Y��a�� ��ϊ��ic���ks�;0��!�Ϩa����~p��_@�+~*�#S�^��iU�Wˉaɖ��y�d���5�ď��8+���*��in#����u<Z%�9�56�hx�G� <^��%!Ӽ:^��!��r[�/��h�N��~C=~h!b �_���-F�lv���(;�yH�Q�~ �E�|�Z�hj����@�{7�-V�Ҭ����v�92R�z��4m�����f�y�b<#�&�����,�5�^�"i���"��N�T幸�^�֞�`�l;t���0w:=��4��:m�D3����b�����8y[���i�t�:����ly��a�Nh�#��@flpK���v���a�\��f�ya����h;F��B1y�.^�wZ�[��Rk ��٪�8<&Of�3�l�l8f�+ޖ[��c)��/�G�+��iXn�?�ݫ�)�C���K�41��a�m_`�����:�dHѩ^%�B,�_�R/ �V�.�Vz��X�`����@6��ʚ��!�^����[�q���/�Ŀό-	��Z�P0UE7,��H��k��u3������CD�V} xU�P�V�Cku�3о~;5���+���� �BŢ?vr�Zi��4��1 *���m��y�`���"��R}��;�bi�����$8��d�z镆)(�>e��]~Rv��'��b���$k�k�qHw`�3�$8�Yt���h9�q�Nx�ɕ����p��ت�Ύs�`%�V`n���]���/}a���X)&NFւl�y��:����G���i�l/*c_�f� M%���y3��}xݿ�6���SSL.�&Ix���F[�-5㫅q窭�m�"��óWe�5�o�ς(�^"��E���☎�`Ͽ�5���H$��RD�2E�!��b/)��4ȚUr0�n��uە�bZZ�{fw��[���"����n���Ti���=��q�8Nd#6%3�x��H����\(�7�r��Z,�X�b<+C��_\NG�8<��K�KSdD>ߚ��?✧��J��u��bط J�Dbbje:�i%o�x�%�{� �����E톒x�^'�,x���p�g9[��_J�t4��~���kGJ����>u�l!��h���v$��_��.�
��� ];�&�T�}ar��}�B��DU�*�f�H����'Y�^�W�J�X���ZX���iq��rW�+�ց�x)��1��i��bJ�R���g��S6͸Z��W���u�Ӷ����zs��#	�@j.f_4�Ԉ�Y�4����Ri�}�&N;����c��sV�w �F �X� �]�]��f��Ezu�L�D�YL�ճ�?��<NDe¿�`���VM(�SM���0���HS�����$�5�4�v�>�+I�R�ݹ{L;M�z�6��O�ޡ��^5��!�ѬL1H`��V���e纏�j@ܒjXzIϜ�ғ���B�@�'��+�~�1 F�[R�rF���x��Z��Y�F$���B�T�B�j;���"�����@���)�ae�i
VNư�z#����Q_=yg�W��?�f�*0�l�z��A�����9q���а<�A����>��7�n����-�|n�:�։��<#�'��zX���v2�����(��L��.	���b��''6���!�¬b|�q�j�:y������6s/��qCzT��a��6(��7�ͯI��4wCz����|�&�U^�tu֬�����aTvC�5��_)��	��I�F@L����sճ�K�����N�����U��$�bF�-�y����
���Ώ�\�崠��E����(DuW��G��Ioɗ�o��OJ(+;K�Đoӎ,R
U�H�ng�CTFe\��`
��5Vm���g*���i	��b�������!�RQ`ZrɀF�@�(
];o��Z@̠9�YI�_�2��_k�ڦ.�k��>m��M��l�g�0��J���eh͂69�����%�N�f7@���'�믯���Ω�%�>Y�f���6*zN,p�'|�r�>2v�/�v��t>IXy���
�,(����Z�C@��:)~5�1*�ۘa�u[��m��b�蚐�"�_���L����zT&�<��p尙�����v�*��c���7ކWX]}_� ��h���~o�6�E��	ZN)w;>\�C��Os���Z�t�#��-�~�GZYG-��n�(�9��p�Xh���zVB��k֭3@P,�=����E�U���Ir���m#�S te&-��!MY�|�o�f�������������c�^ep��ZvY^���o#o�")~yh��{vT}{�2ߜ��}WK��[�P�Il�dA0��(!������EP�W"�1ێ��X�5�M悿���x��mi�m`R�mgU��\0�c��C�1b�+�l ;�h��kI.+Y�h�����C�L��D9}��C֩æ'uN̣�`�y��G#�?uRIaU����OA�Dy�O4�F�r[���4��Z�@�	g5Xi�w^��&/z�khT�h@aݭY��Q/�Fn�Ά����K���ѴB�v0޼xХ�ӈ�q�����J}Lk?#ONJ��s#@;*���p'�Rd+�d���k�2���
7�.�GP���ձ��Q�ǅ��E�٬7e翇_�J��Q�0l�*�<T���IR�J��.���Y��
�+V�A�+G0zs
e�(�)W�&F�UE4�rc�n�Xb��F��@n2��(iI��U�9)�[Bօ/����Etd$N�e��ܡA�)ȭ�Fk�Ï^���w0C>D�E~"�H��<�d������H 2%,ƿq����.�$��iS�� m�]�v�ʽ�
�%"Y.gi�w������[���5f��PG�����M�&p��'�Gnс�G�.֟��z~�=cL���e��1vk�����b�fŖ��'"�W� g�#�z�BP`��������-���� �'��,�!:U�m�'��
�u3��wf��'`ߋip.��� �b9�1��@Q0�b���:��ʄ�Co��k�j3��t�a��tz��9j:I�����ۺ��ׂN7�w�Q�1&��@i���K�����;�]��CSKM�!�G�YI�-�Z���i���lx��jsq�q��(#�a�J��r���|nLw}O�Cy��D�����l���h!oA�<�S~~.a����,@B���!#�!�I�(s>��Ԟ��W�? ���A'�lP��.I�WX�)(f���xf�ց�:_�k���WR>o��<�W]s�`��s�ari?���f���&&�1}����`j,�(�) ��3tʶ$���@姸LsAl!���O*�2��A����x��YM�$��|p�q[�ӽ�
�Ts�	�b	�d�b�ވ\�e����=���m�d�L��iq�����������w����J��ϓLGZ����?��-��8�M2��{w��_��F���t����D���f+!�I��q�Mt��&I�ɦ|aCǻh��BL�4�2�3���C�7/�|�������B݆
U�=-TU �� ������6w�}�=?���n�H�{Ji1�� �?���!a��p�,[C�C��=4 �S۰N@��E0��!���l�/���@ z?S].��}�G�ſ+��1$��iYZl�jU�=	h�����`�@��į���|�k-#�s[�Ǫ���eY���
�%���*��G�@��yGkI�
f���1�R	G&1��e�n��c(�V �w����-x�vqgaʶ�I�5�)qhv
N\���-��ׅ�z�!����Ե䭰�����}4��\����=Y�Q[����PшJ������Z�|c`cM��#��H2�t`�k�f;�jߤ�Js�g₠~J�+���W��V��@�]=D�ToU"^�c�D<L�?���؋�.\M�KǊ>�qOC03�P�8H���3�?����D(�h�>�y�a9mUf��%2�.�
�㓲��T����I��(�;`�`&4��8_[ �;���Ě^*�I��9p9���HW��i[����X�0Uٰ[~�8^�)Ħ3�
��(�<��.Lj��w�o�}���.��4+����r��E�09U�T7C��#���C�� w!�߂����!�e�&`$^���l��0~( 9q?ۨ�$F��D��o�_����l��6��z��ثQ�<�\�t$�:c*������Ȗ��2�$`c��;a����w�6S5����3��e�&���$r���h��eу]�}��q��a�� (0Ӕc�x�qRS��ɘM��N�c+� ��߬�X��Z��.�z�Aa���������?�s�c�u��W0쫐�-�G��pX�r�+��)��01���K~?N;-@4�o��� oT�7�̌L�	��~����=����S9�� �X�i��C�x&���b^��s7=���P�#�	۫�B�l���(�w�<�����L�1��^�Q%�d��2�I ^�i�-]��85� N@�E��$��b,j��"�>D�*�͙AQ�y�E�	�|�	�g���n+�:�d�M*�×^���=H����A]��"�*���]fG�,��^v��Q:���m�H7�S90�i'@���e�����<��U��_/��R.�`<G?D�^�o��?�� ��.�)�B,�n���ΩM�6k�s�'lk�|��VRC�3�ʉ{ȴ�dfPY>*�������Y�~_aDެz�����%��"��~HĞ%T�s4���+INf��:RAM�q�7��$���TD/I������އ�j��h�Li���/�D�(I/�����Cv�+G�@��/�O�J�J;�� >*����͏ϕ�̅��*n���x-Xo��.�4~�0$�+����Jro�^�K�p������#���8\w��3�[B�V����걋4���{���7�����]$�yP&c���W��>���35��/h��h𧹫H�X��EHNm�M5�	�Y\�����4�ﻺ��mN�):G3�w�k�����~�Q�a���G`�-(�H�U���!�zc��'ŗ 8��a���έO����+U�ZI/�Ty���/sE�8
q����0�j��Q4J���uMB�����\JQ�����ԓDh{�"���+&�N"ŗ���T�,��v2�muu�f��Y�%�-��R��J���.�;��gF,���_�Ӊ�e�~;�k���,'_����I���-�K�SQӗ�4�v@jMؚCʤ\�\6,ӎ���G�X�ߓ�3otfa�����ͅ]��\ ������
v@1G�/����݌7?N�P�t*��J�U���#S!"�	v\ոep��LI�
ܘW����W!���hl�6�c��2�>Ɋ-4^�aZ��[�v�	�|*���q�y#w�*0�B����x�&��5���bB�d�q��z0>L�٨����ȷ�
:p)��	���H���5�*��6��Ǫ4)��)�Tg0"��|�Q�WoVA1'�U�A���#���ڝ�9!���M��=iLRZ8D��p�D����FP����_�U/?ռ�9�����vDo~��ݶ(�ķ�?T��5s�!@�ז���g��(J��,K�B���Q=,�yo��?���}y1"��s��̲�7j�1�q]F)䍲E�U����;��T�@-��V�gИ�.����[*���DI��K�9�1-U林����l ��:��xf�|}s���MUR��gJ�ۆ��N|�8�u-��GG(��?v3�,�͖�g��\i��9���|� ���ѕ�5�mC9S��߉%I��b$4�es�j�c�F`+m�U]8�a~!�0��>��Mrn�χ��s��Z1I���N}Ѝg|�u�%��TF����ǜ"a��֡�����8���k��؎H�n4��+�_�[ź�>�~�{\ς����>�y �e���iX_~�z퓫�	�:G�|f�T�>~����{]*��u�u$
�7͵妱98���]�7�i��J����up�eb�&UP��fz�l3��g*5�b\��p��T5C#(|�l��p݇���8p��L�Y�	0[F.x�p1z͠ڳ�&'L�ꕃ/���-1o�t	˾�`[%�ձ$ �L���@�2���U�]o���$�;��S�����C4��7L����2�.����5�@���Z��#7�D�k��>��R��nv�SE�����YȀ;W'V��|*���J��:ty����{��59X>�
��$n��>&�?��J6Z����<܏��Q���wf�d���#�q:���uͽ��-3��"���쒼i1�-�9�����F�S��]aE$�Pȫ4��|[\�-;���]|a����Y��y^^��h�Wܱ�-�g�2���ft���ج�i��-,[]�]�Zf�.��<'�EI��Vp�ׅgi��S��E�;	�M�ԋf�M��@�lM7�{�qRF��Zj��רQ�&��+����s�^j��t"�EڎL�]�nx�?���y'�zb��&�S���n'�	�u{��5�'=y( .��ݷ3�
�Q*��	�{�L�"���em����e�Ѵ.���D�VwF#�0��� �'�<����٥�2.�����Wf���l���~띁����~�?��{�<��&��?�}���,��N��DnYʌ����cqC�6���z���_�H�DE��[�rXd��7X��g+=�cD�IN԰����435���2�' ��|��
�w@�=�� +9�%�*K˃��X�ћ��J9��ƻ�(�R��F��2fM�7蜕$�>�����].v�� ����/��t�F�|�	h�9��Դi��0���k�J�O�ۂ	�%�z��HAR�[�H��+���2�F�1���G��c^ү%k p�A��i��_�w�M2��մ)zp�W�F�x�"'��0(���gq�/ �vs�Z�#��Ɩ�ܭ锇{NW¢��n��+���Yq��������-�"n<ޢ�Q�+�"��_�Y�Bz?o�q|*�qZ�S#[��ޏ��#� 2:AAQ�؆��@q�ߘ,�{ޑ16�'LC��mx������\��#p�o�p
��uF��|%x$QU��>B��3�O5\���ӫI~����n�����^��6�p�F����V�:uP�;<��k����2�AV�̭�$�]���4�Bs^D�L�t�:�3VJ\I���L��(����r٣��0�`ۖ5�	�+���J�PD@��pPM�4�V��+���B�):����`ʟ�;���\ށָ�;'x}n��q���]$$8cLzBd���ݒ�85����O�#���6�T�ro;�Ԑ�]k��2��|B<θ��h�9��V�[Ğ�*�7v�o�L�]�x1�����O��@?����w�w�v�����r�F(����E_�T���	�|#X���0�
��Y㗅6��D[��%��V�-Ja���������
��L�'a����Dy�$k?��o���S%�q���XF�e��(�N�dXW�lT#��7��7�@�S>��1{A"4�$Kz���&	F0Rs|��F5ܶ-�3���_lB�@���X��[kɅ����˔B��n���S�>[v�Vo�9P����b	�TZ�!�b~��sܷ���48�8o�HC�����+\س?3\�P!��奒*�Y�g����)�%¼�x8\Ѣ3T�7�!����_V�Cd�q��\8�a��5�){��g�4F7��R��Y<�7��4̪ѩ�9RQ��q|�[�(�;N�Z��lI�}�)\��Mi*�V�F�����ni�u��/� �tΏ�3 s!U�v~�^̍ĳd�	�������\��ErG���S1Mo�f%;��(��ޤF�(n��a`u������G,��D�
���J�#������NqH3d�gH���}.�����~��mGy��?߀��m�sn�_��w��R�2q�^�/��c����*��^�J����C))Nðq3�
O ���3X�`�#o7�����}VѾ�$(.XJ�8zD��VQ3�@Z�|��;��k�ځ�m��o/5d��}e4�Z����Dee6��KG	î��5���-1�Q{c����:9�tT�u�ai��>4B�*�ӎ ⣗<@8cZ�qEgTq�g���S�Ve\�-quX��s�}��?�I�}�Й�=Y���E���^hCM�40�bk �R4!��QH�S,w��� �\��
���� NB<w��yW�����=�X�ڵp7TU�i��M���Y�ܫ:&։?�lxd�^�^�o9U�\���Ʋ3��ie������>�I���;�6�kI��QH��Oh�,����ۥ3�Hsuk ���q��՛?Z
�ăCu��T��7T_7W���`lV��Y�[�x�vn���K��{��D�<g��A�m$�-i%~�<��D2Gb��@DI�~�a O!z��U2Eh�g,��s���C����u�w`!��
��"� h�u��y�>�jʿ3��)5�+$��b}%�����0|vZʅ�M�sWv����SKýYx���ʲ�gaw�����{�p�4S}�l�K�N �s��n���0V�#���l�J�k�f&!C���`��Z.V~O�x���M&�`l��7����}��΢YH�>�A>���
v1\�H��S/���M�}�8F��9Q��і���лa�ߚ�W��%��?J/TF����o�!��}v��DYr���yԧ�T	�`�2�I�#]�;�LA%�m��(��F�Oǻ��p"ffp���^����7G�>Fd�%���KE��x�,���g�����u�"���>}*�o�����;r��ϗ��z�z#]D�(麠D���!R<�볤4�V�i��7>nF�C��?t�S=�
��cg�\��UУ!��!e��m4����G�[�[�����F_�
!.YcZ%m�vxt!*OE�<�����e�)���9yzM]a��+�9mű��Y�����R�s�0#��pld�H Fx����U�p�ۛ��Eր�XrSn�z[ U�5�g7hFi������1���-
`5�ٰ��\t"e�5՛N\��i�JY�?��SD��7Y��87t� ����~av|���_�W^5�.�%z�&�J�H^T\%��I��~�<����Qs1��G�G(�@&���|%��
���7W�eTje�V��`<�����qg��d�S�-�9�ͽ�Mu����xW��7��ɫ��g
-�vElj� �����ǁ�m�(��0t ����X�X!�l����:b�+�;��?N���	�|���ΨL'�]k[�� @�o���I�����#,��p���j�p٘h�"�Ma�d�ϙE��w*%)��=o EI�Y˼�H�ǌ/��3 ���@�כԸ�F01� �go-i5|4���ݪ("��7����_:ЙI4�h�t�����y�II�&��G�\�\��gF�æDя����F<%x�t�5H8D�@����=��.bv�L���S��g*�I!�ק�+➴�O��c�m��^!nsJ��^!�;��Br?-��
J�>K�����_H�����V��pfriv�1������U����"*
z|\3w���f���Z�o�v�W°������R���DY�>u��zdC�P��7�94�]�g9q�;N -4�}��#B6vM�XO��C��N�\L?N
w���]};3�c��;��H�ڃ��*J��ՙ�4�9��sg�BˤZ�|