��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���e���-�O�����x����:��ރ45�[�:��ܕ��'�9^%F[�'-�U{��^xoYc�_�_��]9�]a[�,j�&�O�S���H��Ǣ�o�L�)���POě�#I�b���8��M�Ԛ����P�Jp�pݎ'��ޢ���"?�p����p��9y�=�h_kw)�弰z[ν����'�x����d�<hK�[};O��mv�Gb���Ќ�:�T��$&ؒA�͈69M�^�C�FA�8굱Rt��⬗׮�a50�z�=��yp���*�&�- �4����H(M��j��� 6#���۷�<7K� cDS�.	��C��n�����^ ����J ~�kpi������D�:vi�˯p��8X�Н ����IKd��Z�����W�H���V��T��u���ق�\�h��S/����P�������|h-��DL�����eˇ���۬weO����� |\baB��7$���wx��X�c��m��V
�q:���V��[/�e�i���X�4�F�,dxV}�J�K.r���5B�í������F\El�Ջ�i�	�UZ�ȵC�$	��1]��������c�0K9d|t��JbDZ7�����j��%��y��8�����%�W�E3ׇE�����W�ry���E�EHz��k��2^���3�|�Ӻ�����Mp����}/�����7k�`
���۰��ez�����-�(��W�P���¢��ϭL4�ʥ�Qީ�d�!�d��Z�`_
?@X�۫V_zw2P��E
�<G͕��Ӄ���V �^7O�k�bx	����\/���a������uVg�8'h�(�k��{4n������$V�*/&@�>���\ �u5�2�Q�CN�	8e&�=��GJX2D��==�#�=%�f�?���p 	��5jG�P�[71բ,מ����t99g��tgfH!��k"�Ӹ>[2�G�q{1b�unV>NP`f�W�45�y�/�e���4��Z�?gԮ�X���j��4Ї�Z_`!���]j2�,���m����hB�ȡ����8D�F
��O?��0�(_bX<H��|���A�����)�X젤o�p�0 �=V�u%�k�v ��`�a�ǥ�g�E���NV14q�h����zob Θ��D\�)�e��%'�4�4�Y+Fd����cw�:��,Og+��(�ğx��h=m2���M�o�՟ʆ��<U�.����� �d��UG�/2)���6|;������HQ��"K�ХHI	^�����P��R��K�����?'-*<�S>������VW����[��������9f��,��oq�{aH��@���26�tuy��f� ɡ���2�d�	�l���:)�'&�5��s��$�%����D2��eO��A,���|���V+���DY��aI\�J3\�L'D;�7 l�0�%�`'%�)T�k3$��懪G�5�db1Nu����u?��|�-3�