��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��*�+��A�R$�D�i'��6qG�-}P�j�l�.�,i~yvVw���ck��I�0m���<�?�
��o$�Z��Y�?���W��G�<���( ��$����0��Q,0��T49)B��rل��f�n]�̮��5�`�$��y��S�H���9��Z�.�)1�N��e�a/��d7�qĢ5���\� �i����xl��vaڤ-gHO_���8Zi�0���ZܠkX�θ��|]A�(��h�RfG�����_H}A�N������p���oZ!�S)'�@�m� �	�)9K��:�@S�[��cY�Yߍ��%\�������|�bD�"�1�C�/���K:4��y�K4o1�Ī>B,=��tsk��~�K�>\��*M�`f�M�J��̙ƣ3Z���l����1̬� ���׆��gd&N��&At!����_겗L�F(��(Eů����Z�A�,������:(�	p�i:�d�։���B]�FoR��f��u�|)j�<jO���Ƀ
3Oh���K�=�BD0'�A)\�^U�)N����Q�;
}���,"o�������'<�_ C�m$��1P�;� ~�E��-g�N �B��J+�>g�_�d(U��?~�� ���K����9��6���`���Ugh��]���z@��Aq;R\�t�`���M?�Ğ��$@>������vuk�;������p�QJ�Ϗ3X�c.~o�0d}��]�>��{X+�.OI��fƸ�&���	1��3����J���F�(ݏ�WN�A"!>h�d�T�������Å� ��*�#z�lS�ٶ���ЭU�̨�a�ŹY���1��O4�ݫ�l���SG�Mb�ǳ /W+�_��`���A��Pr��_��(�ƒ�w�Pv'���<t>]��l�v��HͦG��k�q]�!�N��7:���p&�"���^�f@�S"��u���G����\��V�t7�QGR'+��q��Fwe��ݽ��+@��'��*���JM�����n�$a�������wN�!�z}Y9�$�N��a�� ������t����� �1<�皋{-=�� ���O�=��9��y}� 2N��SIc���Zеg����'"�xnVף����ழ�� �2�1���|�찏�,��b��S*c����"P��ʨA�=�é�!�j߇�G�%v O�_P�9��������<=��#����M��&92���)��֤��m�a_0!� fYl6�)��^3Y�G��֜bl���A��f� �BQ]�z����l<plb�;�o�
"|��Î�hF2Qh6���mE@�+ï.@�/]�|� ��w���W�R���8�Q35T�Ko8�ل�R�\Z囹���ދ��|�J�
����Òc)+�d�\C���y<'=��wA�ie�!5��%���H[BMK� ���؂�+�P��Γ��f�v4؆��_d��7�~_q&��t��iJeo����;�!'�(9B�X��~Ü#���a��v�k5��#�3�����@��1|!��	,g�w,�}��j��l�4������"h�m�4E/�?(KP�O���tIY�Q������sq���L�;z<� 41�i$(1�ax,)]ڊ��W��1�Zԥ�e�}��T��d���=zGG�s���C����Ϗ�%�UFG���-���=�~�A���P�_���8�w��Ay@�g+Y�6a�B�GE#P�g]iq���VZ�02�5*�ű����&���Xo gy��]̿�.ޕ����*��n2���}ڮ���!��l��F�B�q�HBq	|��ׇd��8��K�H ��oR;���O�bٲˁ_V�Bua55/J�KA�Ҏ��t�J�a����c�>V#��M�j6��y���&�����̗c���앞<��;��9!b���l��oq	4@�6q\�����U�)A	���:��q�=��V}RUq�F��)S�>D���0W�$��(V����@�d9��E�#�o�o�^��/mv
��S\Y_B�M���K��O��󉢾��(���&�e�f�pWt<J�P� �&���� :�0h��$�\}��]�΀�.{���a1t}߃jT��?%�V�#쐀Q�=`��'��z�B��fn�H�>у7�<.{ b��^_�v��9W/�z�0QZ�"{����J�Gtn�/:ݖ��V|gb?ۄ1��"zX(W�}�~n����V?�"�g�]w����ji��&��`s�FGC6)�WU}r���Y(�O�b�)�s��Ȃ�1�Pp�}S�$:�UHD+��K7н}�Q����l<n����iN6W����6�]��(�mn�~&1z�p8�N[o��V��0K)����F�ӐܦG�ND�}`مi���F1��l�x�n�n��i��ꙛI��e+~�.��eQ�I�;�t��Eg1̮S�b���c���}2|��/�ׂZc�Df�C��P־�s�A���v�L=^�}��'5E��9�|�H�l�`p�������`@<%a �mG�A�('Y�*����u�eҀ�)�øa���d^��x��@�^����s�?XW�ɾ^PQ�Iݶ���c"�&�j]�lu$�BE����|�wwPfe�� ��)~��Z����F=C���~���<ݖ�����7�ށIU�RXk�&�ݎM1�V O�p Ҙ���2G�n=��R�3u;O]�s��o������񅌀5pgg�~�X&S���~�N"��2!YIlo27�$�Ha�H1�M��]�[�5�Ac���A;@�y�xy�KC�H�)6Nz�D
p��ō�M��v���i����ETt�ҡ��#¦{�i���O֚ߑ��+k��@P�]��
G#D�f�e��XhDrç� �~hPV!lA��;�EF�ȁ�7������
�fT�M֥��Y���<A�M"+�j$�������&!���<�H?���l*R(T��v�[ݬ�(�7�OTo��7����w&���u}���$WD��oA3����M�q�ފ6�І�Z����M_}7��yF��";޿���ֻ�X6	�4��.�S����T}�o&~�����TLUS~����SLI�׽������3!
<��)SJ?���}n��\���3�ƻ!m�ʺ�$���Ox+����]��O��
N%�X��<L������$���0=��l1dr&P�Ռ�mL}9��])���˿���v%bٔz7�N6��[rb������ϔ ���ɍ{��F�����>�����#>�U��+E��Rބl���z/f
],�U̓��A�bY�o����+W�d�="J�`@��5Vߥ����0�=9��3I ̱�o7�琐����\�kG&N_��v���g�|﯁@\�'#�٣��i�flzI��۵9nw��⌁y}:�Hް�ET\��g�6���m��E��j��{�n���dc��n �2,���
D7�jW_D�r0p0Q�LQ�����ic#�3�,9��c�F0����א��=�~1�S/�p�7]�`�h�^Yd�����,C�$`MA�J(�Q%����>`ك��ǻ��j-�i���D���j��� �([X���$_��C�ؔl���2���ip�D)��n�-J��c-��P������� �vv�Ne�`��Ӱ�y�B���S�8�"/��qM��釻�|��8Ǟ�)��k,�K���ޙr��Uİ�
�+�޼f�K�`�0�)�L(椼�Y��0RNʦ@��N1���{���=�}�Y��>Yz�@t��]����|��M���C���GV�g7�,z�њL]�n�.�p�)CqU>����x��n�"���_b8�����Ws��
�@#�s��x>����}�|�{�'�q��Ba3| "�4B����U�]L�Zh�%���ne}��Tz�_�E���Q7�7 �'�V�[Ca9�m�I������r(w:�v.?'���O��D�:0� ���ڵQ���!���2����w�,�1c�Ԛ!4����}�)P�i���I����HS�`�ʍ^�at�0���饡����I�iv����;��=2G䔼��$j����O����2r&�&�zZb=̬{�^Ah��!S9&�u���*�D�E�Vv�.��[t�S|�<+@��h�<��q�as��jR�V�N���7��X{�'5���C�H�[c�=J���v���Dg���N��&|�M�����ص��.�$#}m2��Fj�&�@���ٱ�=Ua-Dm�W��D��2�����4ִhzƮ':�1[.�+d4[tGu��������2�����-�D�v��{���+K>��+��7~����F@HoÊ��l�,r� 6���\��e��t@�S~������?���vZS�
������WZ�@�#���(�x.�|W��ګ(���dg�.��0[^�:!��v��/���ªL��$���K"�!����pe�|���������`�ß��E+7V�D�PG/Փ���ld8h��Hq�re����?�f�J����������4$Kit���L�э�y*����
����27�5[�|z��r�҈f�x s��Q����o�I��	��f3m"�fo�k�\(&��8�B�G��v���8on ����In!r֧Y[L�t�*Y����;Ǭ-ӛ?��H���ß��(C���"ȋ�]�^p}p�� �s0��!QYy��1�/ӓe���lp�a����]������֟�: �
�vQHL@]�bN:8�_P�������,����X>�u��짳8��)�:������w9��x=&���K�GV�1���@z�m�v��4�3&}�jtW���Z�5<3t9C�XI{1�/ܦϺP_���������f��}%@M$�P��,ǖ����k4O(�'F����ݒ�;r� L��!�9����]^�!��1�$}'��;�]�'�I�O��mu��p0t�o_�!��������"�XS���ɓ����v���I�TVX|s�(#�译�}�!�vݜ���_�:
���1>�TjC4d�����=��E��?�5��~#c�� �����~�ӽP�\���Ȭ���B=�e��`���Ѐ�ۇ�;�)gH���6��T��X�U	AJ������u9Ǌo�;�U͸�3�9FB������NW:>�Gr(Μ�A&W�s��AUvy2iE�S7�Y� �Og�g��,���-1��-,qy�Ǩe��  i6:0q2�����������������^���],���Ӛ�`ݓ�&}��u�ch�Q���� A�nPzW��nQ+��ʗv�}f���h��}���E�L��ا��_�L�.ѝ�Y;UH�;���&C~t������j2�b��i��r�d�2��.Y�'��b�bƉ�"Z��Gz����>@	V�Y�6�K��iq?HXm�{�eK�' ��i,E{|�]<��� ��Fe�0pх�GH%!�&8��u�N��oc'�̕����ޒ��0��
��� $�j
{*w��d��T��(��(c�k4�|�d��e�R����v4M�@)m�0��~=L����\�	b�C�\�{gK���e�[��.�RGD�ȄֆB�������̞���ZGi8���)���M���������ki��B���(G�(h1Ԓ�cJÐzW�-���G��F�/~�b�U�`d|�x�pa���4�^�O߻�c�	mv�{L SՏ������z��h�t,7��:?b��|���xe�p��n�_-�x�J���R�=WqC��I:(խ�]����u�����4ݒ�5cb'�dj��� f���{{_����Z�c��R��B�L�bb�oj<l�J�!�u�YQ�f��\lR��Ծ�0�s�r^4e��7��c���G�p_.����߀�BQ�	�Y%��B�f�Ұ��Px���ݮ��з�?,������8>���bBZ���m�Yt�!K�P�����[X��\�j�.f�s���ww�@���1ٶn��ނ�֥��D�,n؈��H�O4�Wu>2�0l�u�ԙ|i�4~i��ȕ��^��n��=�6?��xD�!�Ñ9Q��?X�f��i�J|�Υ�A�OM�U-h������_��xM�C$�Wyw\ԥ�n�����k:B}��d��IZ�����%̴*�w��?�W屗M��}CEP�iJ��Bt�t,|�!�?ۀ#;T���W$�OEg��P����q�ܢ1ȷ�ޙ=,�O���m:)*}ATnIZ@���{ԟ�J��)CB�u�&�X�H}��ϗ�����2'��y3������9�n����-_v� �������c����Hۣ�k�[�d�A�?��_X�e�"�������	�E�?�����}��"��v5WK	�l�A!����m�I���>r�Q��@qb�{�Z�]骮�"<|��2>�D�G8#�Pt���Z`�|�hǧإ���n,���BEi,�������?h��|�d�Ӌ�'���#"�sOH(/[,��"���X~�.m���ެ��e�K����\T���K����v��+ťɏ���K��gz�G6kޔ��z!/��~��C��Ǉ\��-��XP���������Z(�Ds��DX��x��>mkP������j�Q95��"ٚu���G*��a>4�I.d�<Պ��ޓ)�����^��u�+oiI�������,*�8�K�,��m�Z�d������]�4�i�;1=�L�/]I�Ec����Lr�R������AwF�T�Q�-�e�'� o��B��+,�9l��ߴ;���G� ��v\�yCUY�-���������4Y���FV���n��FQ���X��S�3�h$��rmI
><��B��\&3{�c��.n��w��"jX�l� f�D Q��� Y$�kT�w;S������(Ps��@W���'P6�:6oқ=������	z`(,�X�����aDj���o]�s���jN��Į��vt>6��!O8����^�rb�P(5`nȃa��:6*%�I�z�>b#!q��|>AB��E/x����g�`k�q%1A�?���j+�#��A<>�>,���x�P��r`�9]�����j�2����9ɵdy��᝙6મ ��+9*�r�����
=[��}CQ�]|���S
��1b����N������@�O��^��ѝ-�M|����$ـ�7g8B�`��D8L�D~�VڼM��%��fm�M�l##�=��yj#݁N�ql�,X������0_1 �ֈ����I�d��[���֍��Wl�3�>f��
;q��Q�V:�x��8����\k��v�]���:-,��m��9{4@�Lw������t-�<r�	�i�J9�Aj��{ф*O�!V���5a�g׊>��}?x�/��#)�~���~����[����b^x���v�ŖM���2=~
��&FE�p)^;�ý�c�QV��lU����ms_hl0a ��B�|�*��ă�*T�|����y�û��YψG�S��><+��(�E?�����o�8�X����c �$l45M~^R�5/3�,A�w��	�������%ZKq�v�78dZ�l�	u}dk���f���ǵJlw�DN#s��)���`T@����w�����O��G�' ��t�&��5�,Cc��gkE��� ��U#L�G�`����ԧij)�n��D�R;�Gz�	^�m! K��|��'�?Oc���ŌX��nVj���Y�W%.6}���� b=��b�c�d�;vG��P�7���Q2�m�5�p���h��K��p������jn�%u�u��j�:�6L��݄�l�3߭��9�o�����dٸR/7'�&��[��.	���#���@,��$����|;�\�Z��n]�����Hzݽs�j��X�AE7A��e�	-΃5Y�"�7l�b̮�y`�S�;�N|9�3���J�]m]ؕS�������hC�Fe�������0fs���ť��#H̔��*�x1/����떜�ɝ_�\,�I�x%p��J���״Hw�!��I�A�Eϐ��[�LO��G���P�>I]^ޯ�$���bN�a5��~�_��cVF�:��lA��A��OR�u�F��ŀje��9��H�/0	S�{��ۮ�����E�����{)���R�S��C_�D3����Ϝ7CIX�r�Ms�������ah������S�ti�T1��^�å�� �]0���g��~��;�� �L.�����a�N��E1�3!')@�Uh�8��i"��4v��������D��1�|�où��w6U�"\*��D���o�C,'$g���ދ��6O���I��'�����L�Yת�i��7��aMV�:0z-��koV$�yy�I��� �e�#�'��m�V{���
�h�������l�rF t���j���gl�7�ZK����O�T^��uș�� �s�3��ZeJD�BP)q	3z��,2ր���_�F]�@�"��@��lVE��H��s����c��Q;
�!ͭ�/Z��0N�B J|�{�	Q�z�����7�yU����������{��#�����@p�#�en�Emv
}au]2�Ÿ9��eZ&�
��W��kQdY��csH�Bᶀ���u;㏧���/� @d/�1f>k��(̄��˂�*,�gX�Im�B�ُ�y���2�1�ZPTWȓ���9E�X�*�q���d�J�h���qV;��.s��8Qձp���()���.�e�E��l�_�T���?佨���FI��M�$�
������x�Q� �;,x�m���.|�Ur1<ׄ��h$q���B�t��b�tٟ�M�p�%����ÍEP-�zʀ�nH��SK:�ٍiaRܓ�X}��8���ު��uf#��gc�׾��,� ,��,i��x$���
fc#薛C���~>z`�9�6�`~^}J��0-����c�����(�Ϟd`��;ڔn��2X<;���
�����!b��#�r:y����V���^�r��D@_����V�B%��rZ����I'��_MQ'�E<�=KY�Ѯ�%:��fz��J��]���b.G���:Y&��+)5���^��X|Oy6%T��>�8��C����ӣ�r ���ynOG�� b@P���^*8����
�c[�A�E��6�j`�]��^_T;�٧h�]�ddX���a:�R�~�������t�۶/��R{r�d��ő�5��}7L�C �1P�	��7g?����e���C������4�Mh���wUx��9���b4次���3�,�i�y��C@��y��0i.�yg��Fj�%�����;�0-�h��0�J3Y��u��8[H�ԅ���\CT<�܈}x��gI��g�m����۟�������H�h�T�G��孃ǒ r�������Ҹb<��+Ј�o�s�9ڠ���T�a��2�hI��M����� ����*����>B�>���7:����w�D�j��*(��=D�,��=y�R�>�C�D�%{��c'd��)�/&T���̾���3TDG�����RQ�Zu/�RQE�Z��Q�wk�;�z�o\ k)|X�y��É����82�����tKY��/�����%l�^7���ҍ>^2VWΟz���8�6VJ��M8�)���p�VsI�O�(>�D@O7��n�奘p̒�׼�yK���g����+�PEU0�;��5�_`���M�%������;Ì�ޯK��6?�r���ɋH�u��t��s�����z#�p�h�fH&�$ȵ'/�A�ښN�``}?,!.��޻�z�.1�_cּ�;H3�hh��3��VE-�w�&d=�f(6y��ŏƿ���{�υMþ�t!�Pgc8kW�E��[�M���,a˹�\P@������`�UyenQ��m5z� u���qh�-O�D�KE����S��v/C��O�^�꧑8˹9��q$L,"c���O��fx�	���=���~5#�7,X83LX��ܟKZXf�=�N��|D,8^��ܵ8����j�&3�������)4�$�/E�bO����C�>eX��-�����;��z�a�D�W�����+�e�)�[�J-c�����
��]l�[^��il�z��B�\�e؏��%_�k��S�M�o�w�?��geMP��mA��~��&+���a������w�$�l<�c|�3|48|�A�/��|�Wmw�}Y���d�n�X��&�0L��7����3���I{�,c���{���9	�k�Fz[��p�.�U��n��L7�lZ��E���9�}�Z��Ǔ��]'���%���;T� |��NE��5�nZ z�)�Z�Փ~� a�[#q! ���X�ט�kc=�#apT�,�<DI�!��cG����7��
�����E�����+�x���b���i$7>WSs?��_N�|�w �6ƅ1ʂ*;���B��aH+N3V��Dzl��z�g�s�O<��_=��O�A�M���P�G�_H�̔Y�$��S����  ����M��JOb���aܐG]�Io.�ρD�1�EVSU�_����.uآ%4-�t���A+a��&��:�Dn������6��]#j��K�#ȂB�&��8(�.�W��m��
G�+�q�# '�07J"5X��'/ٹ�J�U���1�\� ���Q/����Ŧ�^�$ʐ�Ķ.6l�_ԁ��|��j�AO_��T�l'����f�|�:�����r-oY&!h�L��0W��F>̞Il�#s�D�4�z�G��2����߹X �3{nJ��k`V�p��m]>a��q�H�	�x$v^���k�8��߶w*&���k�5X3�gy�f��[�-�`�X�^/ǩ_YW����%g�?[!���w̲�<(�V�q���z�O���c������Q�it�!����,�Ӏ��p�#�e�/������@6f��R	��gq�«���K�tM����@VzW��ub]45d���_:83��X0��/X*j;(�� ^�=������8����{U��4�i�T��-�8^Bn��E�'�	��, �>t��\� ���R�۪�s��B0���ſ�gxLcZh���YOQ5�i^�[�4<�,����Z�D״�O�}��Gz^�yu��ϳ`@��_uH�������͠ذD�~�;.�z0�)�e���ק�nAU~���EC�;`�W�ת~�I�-�f�	����p�8M�ٷ.��R����h��k���Pمo��7�zm<����~ �a+�a�a?~�W�2P�k�jq����^�:�"�_f�s��p�/���~�i��ךN�=�@r�p��n 
[Y��i�0	dI���)�����
%L�&r�����W.�ͯ%���IuT�Y�P��
�P]F�b�cwk-ۼ�s�ϑѮ�����U�AOEנ��*2��!R�96�h
�ռ��c����O��ĔP���G�%
\�"x�V��]�g֧���=B'��\:�*�C1Pi�4K��>����&N,*�k��^��Ǒ���\�	�Up��V&S��}W���+̈���m��D��an�?���;K�%Y����)��AW{C�0v�f���FQ|�Z�͂����fct���e���2	4��n�I��?	7j��8��0*�����O����R薦���������|�(�_��J��= ��pPj+�)���:`��#�Q}q7��oj�ۨ���s�Ep�Ï�7��3�q�ݰ���Ѕ���H�n݉��,�EG���c���&Z`�
���~�%}�n�P����8��GGCl	��K��?`>~��q��,ǟ���jF��{إ�����"Be��C�������5n1���l�W-y^Ϣ5���7�����=��x@�Qd>(�)�['o85\6��2�,S����|���x�C��s4���.��n�/�T,'�,+�G�0G��!�3̓�x��D�"�;��{��)`��0��\o�9�k����g�!��8��
҇K9,>�[s~L�����pl_�)������t���U�d�j��pa#�Wwo�ƍ��X�=] 3I�.��Y��K�O��WT�d�Z�N,�|�Q4%ġ��?B6r<n�ڝJ笞����6I����j����W<�>�h&&
�3���?���U.�%�w7A�Qn�O�+����sͺ~�a~2zI|7�$L�ETR�N��a��@ڈӰe�WNކ��.�:R�}5q�
s|����؈�{�S�)����H�@�	lVL��ehN���)���q�/�>���o��q��2�G�j��Y��lJ��ж�p�jG�%��_@�ɺi�
0{����{�S���Y�����	+[c�7�H$�w�Бe�aj�#Q�����;�q ,Ro�[�w�Ob����;�A�����g#$�
z�W�^��Z�	��X��ߏH ��Jpa�V:�^
�x	��db�XA��L(��ͩc�:�2�:������完�|~�M�5a9�Q.�	4��u�`��E�m'�Ez�e�z�Z����Q0���J���_uzP�G��~w�ϒ�-9m�yr�Y�ΰ�/�;�HmS.�N|9#ϗJh�)�xڥc_xr�5����7<��
J6�Y��x��zZ��T���P�C������$q�'k��`|p����(�S=(����j�EK��!����F�k�(�[)�'��z�$����������>�x��R6��;_����+���k��<&1W��;!��]���J�aIB6����^��P�py4�Kz�6͌���uV�덵8&���=ĩ|�}��T��h�Rfih��h��|�c�$3T�;Sֈ��"i��_����V4e�-Q*4�OL�K��	.�]��VvF
?t7�R�wMb�=H@�U�V�p�RI���Ս	�.�qrI��"ф��/$KtВZ��7�Kjf���We�w9By���z�{��Ɖ;L�D��}K\�7�Z�M����� �/|�����z�i�!b\�w2��1Ң�\�k\v�n+t���h'����>�]�WM�Ꙓ�u �l;=Y�9��<\3�l·��j_�~������k'*쒮�R�hO����p!T'��@�C�����޷͒�g&��`A��	فk�9��jS5OG���*%���͸����ή*K�9f/�&��Y�I�F-`l���a�$������A2sWSZ�����	`�%�>�Nq�cs�^���@�[�刟��/�]�ĵ��fܬ��?�zr^���ݻW�r:��
S�1����kmʀ'�ޡ�՜  2�k����E��D:�CZ
-�N Ґ���3�Y�I+�=&�h����~�)�ɞM�Hi>��H-D�n�E	��ϴKR��I�^�)��^q�b�~'�<��DzU�.��TIy�|�e���Z�m���Y���h��*��ty���kЌ<�1H�u�����"�!�2��9�U `�x�nA�_�ہ
�v_/�[����aȍ�R<�$���ވ��:�
X�����T��䑹CSm��C���w�W��]��s�(��z5������,k��EO�E%������Kh�*��#T�?ě��e���58J39k�90��(q�(��"�Yڴ�B�w��5_�8�~�D�Px�O�AeN) ��(y�HfeH#1W�oǇ|fs�8��*#�kŷ���_�c���#-��!�o�_�>�@X����sƠ�g�/����-A�>~�ǒɨs�鿇�:ss�/�F����X��K�ZK��K
'������.x1�2!�������y��nl{F�`+��(e�mh1��0\����t�t�	{2-��{���A���c�`��C4���,7r����E�|i�.[`��.^V���H�Z^���Rg��9�C`��0���L��L4V������GW"Mc���5��׹�)�7R>�0����5o�i����,p\(����V�E��\���.8j�
Px}~
*�h���iW֐��]�K�=~�/���pA9Q9�LT��n9~����d'(f���Xr��e;R��d[�H�+�HKO临$y�23���>�������`� �rd���<�:d��}G��� ��)��	
mxU�VC����s�����ܻ�õ�t����dn
�nO��Ä�5���}~��$Ӌ���H�E��F;۱3͓?Ŕ6;n�G��@�5r%	�oՍ����p�DP�����MU��͉�Wm1��,ny�l͏='��k}�Z퇊N�r�#�J��C@�VϜxQ�]��"X�y�ΖS!�0�0��N�T�`5Zz�I2�mރ�&�0�������pe�#�Y"�KwT��ۤ3�zɦ�G���>MH���I�'�!@\<�F���_ꒈ�B#o��v��_�L�*x`�r�7��#�Qu0�����A�	e��q�p��\��U����:���`�S��m��:���b��.����5ɩ�t_s���?�m/��`y	�>Ï&<h0:� f8��(�;��[��>k�iƢ�yd��O�ƅ�G���V_�8i9A�*��"Ѕy�,�݈ŪHAC��9x��(��>�������Y�=kCx���y��B;�Wg��:��)��Z�Vϕ�(
�����XhZ,d.����d�b4Cb�W�%�bf�Y��x�s��4)��rCĨ&�͢ݿl�d_p<.K���P��m���oP�n�ܱ9wqPUZrt��w�+d��2|��f\L��z:�e���*v ?$�*���ƹ9*�cD49#۫�c�ČK�S/8������LZ�$�H���e�A��S������ V�d��b{=,1��G�����ǚ�D�̕.!�5��� DS.:ʛ�·9^B-�.��%H���4g�>O��{W�-f�s�1���AY�z�/�nVUp
��e��n[��d���D��U�#S U��C���U�p� XiwJ��`��j�t�q��Rxc��A���Q�<���Y@K/�b���{8������(���*Z�GN[�,�c�{��w�ty��ҍ|WWT�s�o6��2������t �_Fcs��Z�a�\��-���aW3�Y��|������[� ��Xl~��p��W�po��ls��&:�[N��lbݨ�+���-���Z������B�dC�n�J}g)m���! ��%��.]c�Ci~�eLJ�(fu����5�5:��jZ������3U�A;,�a�1��pG޵)�����y�}6�ɲ�H���%D�2���r�k�?�-r/ks:��O�#�p�!D���t���='��&1�O���1�5MW���|6�a �n�����
l��x�=8�*x������
_�/׬ ��g>e݊����������l�2��Kg��<D�enz�Qp�mo���^ y�gs�N�ڟKH�S"Y��ڃ�lU�h,���}�'j�8�́ H i^T�?�� �5���NY5��T?x�9C�: *�'��󠓑����}I��lV�v]ڭ>���)K��'�|�L�z��<��U�[��m���%$�-��?���H�>+�f=�P�v;�h��3��XdI�w�]X ���*HW�q�s�o�$�c����
�}ɔlF��.1�=��S�"{�!��4 �%8Z�7~9�=��Tz���u$	��;�N
Ǟ79Z8Y���K�)M?/�����vhO�P�t���</d*-7hR��ܯ��h&̄7�"� fD|�	�G�N5E�r�k�/9��0�S��V2��B���T
@��>��)H��8*1b�c�3�õ��pQo@��o��a��h�yQ�Gq��<�J����9�bo�sԙ��L�����}D�$Y�C7���.v^�d � �j��޶�\_�Xr��1�#��U %u:7Ҙ?�C�.X���qڄ�c��Y�j4�e�K���r�صL�H�3	%�J���&Wj�ã>jH��\���;��>��������X�J��ts���u��L��-��O����/�HD+�O�>�7H�cM���rN
4B-����N�x�IJGG�}��-������k��r:�����Ɖ�爥�C0��R-Yd���/�^r��\� �	K����(7@r�*1'��==y�Q��u(
0(��\�/�������^P8�k9@����)�cUe(;;Ch�U�%���H'���N�E��X��\6�Y5�Ĩ]�]8���Yɟu\f����zY7�;�����I��X!�o;�XT���,�_�6�^_�T�#�H���c�(�ro������STp���#���~����B�BB�t��X���%/h���{k!��Mq�ھ������졜�7����,l���Y_]L��v�A�e�s�ڦ�*9d�����������3�[��1���5�����tV|���{��G�C?-'~VQ����-^�SGD�>B�f6A]��lR/�v-�	#�ۘl6~]��y�z�8��Mf�Ý��� �� GQ���=]\������
��GM���HA9M	`:�a�a��e�*X=��X�ꛆ}HQ�v�R���n*�TK,A�u��������,����u�x��N;E���q���q���m��!�T@f��w<	����/�eF6F�}Յ�ԯ�,ο
�"���R�_ґr����CF�	l��Gg���]�;���O����ΡȎ����!��fg�Jh3� %W�qX{�^؎q�F�f���u&�7����+h�lHVK����zh��ug�)8A9�FB��a�tގGi�4�F�	��R�&$�Kj�Ⱦ5��KsJ�P[�`5C:)U呺�I�/��731��T^"��YmT~��T��9X7\Y��+��U.����l⢢$K0>���e��>K\F6�\/����{-x��9cx�G��Y>�\~�Ě�IB�L�7]5�'��Bi<A��f�d!�y�� ��+,kc�l�N_�ý҉�l"�Nt�ۢ���w�h��(�Sq����Oה�w�o�/�Ka�Ҕ��/~�Т�e��%��(0u�����EA)_��}��t@��8>�|ysI��%Y�:8����91(��}��������\+�{=�#�Qk�V�����mW��?����jK>�9�V����{��k*o=/�M���ş��ca�]�:�.s�.��p�V��I�ƿ<��HR=n������+��P�������m�HJ쮭w�{h�']�Yz�����6�I��{��`ŗ���*��,6�&۬��!�_Z�7�:�\�; ��J\�X��f]�:JF�A���s��0��� �POtW|�	_��}� y��xb�=~�+T�NI�g��p��X��])$h�ǆ�޳��CE{ڛ�K�q�{s�n��}�P�B2��8�r�f�5%�m^�!�C�����1C��$��/���b�*TS�滱�nɔ��u��5�O'{�9��*w�uF�/cR��2W	�i��d�V�@r�%}B�G�yO 
�h5�t�Zp@0!e
E���B���*,C�(`3ЩE��˦��,67s3}4�p��Q� ��]��;.{'�?�w��g�����|F������*_'ق�����-kV��ڥ[� �<Cg�^�{��ȉ9%VN|�G�Q�D��j~>?Ŕ]����;�>�fz����S.�Ō�0�r�$������~�N��#$������}q��؁,��~%S�5���|�>!e<��K�m�$��MN�L)����?���j�-��1+P+%�zC]̛�ּ������\��KM@�0&��0���Wy5��=.4!ˠ����exש�R�|ȵR���ɘR�a��'���ݡ@��}
�X$/��x�.}��r`.�����9b�R�Ϝ�;�8=r~G�b�+�L�2��,a��F�[�;�]q�C��+�D�~���`RE�=���x+��[�<*:=xWJ��be�ͨ�+Zjڹ ����4ˠ6H$��[3���=A���<�Lz�G�D�9Ժ�N�����ϟ�Q�^�ӝ;��H����f�kcRɣ���2�CYy�[�W%�i��=;k>�/<��c&�}� ;�o�V��2������!J��[t�c[�����P`�7=����oH�e�@�*,���|���Ԙ��;tr����o�iǃ���A���'�#�� q��S�g�cr�ƶ�EA��3�R�PO��M�R��������i>�HG�E���ݗɆ ���q�H�S�>�0�)�����@M�V֙I��|i���숇����-cǖ��%�l��=�dv�Zw�g��M�o��u���?��P�M�gD2���unxe�>�[�險t���0�����߯(H�R��8���QK���9�݈�.j��u��AY����L5o���,����<�񯸴�h�
�#���!�4�k���}��D���{��z��ủ�#$�R�!��s;
��iS��p],=��O6 C��|	�	��iE�@�X�K��~m� ��"7Zy�KH��#M�V����4�@"Ն�ǂ̹���?����QUGq���+Q�4�KM�L���P���V�!o.ڍլ �ڑ�*����G��o�fr��o�%b�F�v��R�Is���iE��Yσ-�i/.�^d[��ϼ���v�XBYD�8�7ݿ��Ъ�-��`����LSZ�I���(��Pf����Ff0i���D�pǥ\ȷǈv����؂��0.�/k����3qcB���>��ڟ���!X|���QЂ�O��_�&�ɺF�hEz���A�k�I�k/i����~`���J>��O2�їp�o���͊泪�N���|Ӗ��SP$#O�֢�5%� ��Zx 	��[B�\G� ��*�9�^��A�>�����rx7S������i��D�!��<J�&-����?>rl�n֔���� ���a��¶yj�/� ��U[kz:���sJ�"ګ$]�{Ш,"�4D�sd[X�7[U L���m�fW��l�Rm�S�߮�@;'JR�-u;��X�o"��)�{jՓ �i�*�n�S58/��@�r�G"�d���d��������E�N�v YӜoO�z��?��������Qj��k�%)<'���j4'א�!�6L�g��-�m^�].Q���	Z�,�ly�*K!KTo�T	MQx}[�����4��ԛ-%�F��|ʬ-*�k��� $l�ʢpԄ���[n�~
�f��{D�Q~x��˸�$,W�|}}���As�VNWW�|���S�R�LUTN�?��[�
�f.�>RŲ�u-��Ȍ�e#�i7x�$��0�Ù��s���.���2��f��UO�.[���!�E���qT�;�p�}��&�����sM|k���m���~���f��4��aӠ���y�`���͠�O�YQv�O�O^I������l��v��1�J��4�ϯ��[zw#G����GX?��������\5�#�j���j���S�%d]�S���^f�e��dT]�=�v�2��:~Æm;�T�TC����������˄$�)�[����y5Մgqgܹ��L"�[���L��p���"�l���
��e���s[�IF������H��儉�EP�&#���$�k相8NŰ�y)s&Y4�6����(R��t�h{_���q��M�<!�S�d/<�CcA���ׇ
9 ��:����Ҧ@��oɘ��|��aq����_5F�������pӎL���m�p>ff� ��_��<sr�[n��x\(�
���I��z��`����3A��y.��-ۇm�h>�����/q"y�?�4��|ﱊG��-VD��\jT�}��ju��|J����^� ��6����g*u���u���������/#}�������a�/�P��HT���(���207K�,2On����A����8�Q;���Vl'�d�Jҧ;�i!�
�KC�O�z���W��r� 3$���!��� d���0�P�`�┞L�{^����q�@��̃V���M�^@T̺������˳�Q��E�� ���T��ǃ�̳ʅ�7#�Φ�����i5���t"k�ЙgtO�1�'=ms١E������h��sJ�K{��*�|P4ڏ����u�robGI��=�����V��F"��G�b�&��g�S��a=�RGBx>�j��/�4UdCx����$��t��d��G;Ԕu,�'�kA���� �ϻ�8�ŗ���!a�v�|��O��X�\&l\ܾt�l���q�YD�}�Fl���u����+A]5��xn�1�m;?�q��Q�r��Q�0�le�δ�	�T��a�g�r83�x����i��u6��	�
B��ݫj�����5B�]f�h;�2gû��i%gbr����&W�
�)�z�&>�J ��G���&<e���1a94F�77��Z=r'��C�u�B*T�P/�bK ��s�]���O��Mw��� c_�-��߫(��!h��f������OZ~��԰N��r���# �����o���<�}d_����`�E���9f?��@�b1�{A�%6(�g� $�]�U�%��{G��@SԞf�������[uA�
6~��ſ��qG��a���6�3	)oL�ki�:Q�m�l�'&�[���z�/�����+�#���-Cd�z�S��@�nE���$'��QYp�*�ὅ"*.��U$�=��;ABB��851: ��ˮ�h���iLkeu��g���XWM8�1��]��^��D���a��)����27�J�L��{^ԫ��ո�Cݭ���,��}�-�WEo�|�A�ܶ>l����*1�V��^�~�M�%�:f��
��k�u�����Kt���rW�;���~�j� 	I�?�a�n\"���a�Ds�7/A�\'˸����/拾ğ�F�����{<l/���m藐��	>&����ed?a�S���/���!G%a��Ԁ��hļUzox�DBt߭8&�xB�)��WB���B���F���j.^}�Y�y���C��m�Ƽ�`��@yr�ˠ�+:��VL[�2e��vgo����1� m�ہ��g[�R�S���`�F'�|���ۅ���]�4��wʍE�wa�=E�V0�a'��k�JV*��c(�!�K~�3w�H�qt�&&)=Y���i��g�\ܿ��$qu�:�e ҊD����rl��V ��s�0ߧ��lx�"����|t�┦H��D'�~�VZ�����i4b�����IR�)P9�eWa�3� 7o�V��D�L��{�Bax��ߐ}Qh).�ع���,"{�+���D�eR�#�t ����yϵ�2�cH���ɰ�sO���;�w(��x�KBR�C�`8�ߓݼ��7�rN�Q(����0�A��a9A7�[��C��0���K7AX�ek^�"�F�V�PKz��@��]�ȕ�����1jZ����3�3�⼨^'���.��}Z���Q|rHU5Ǭ5A�R�t��)��\!:*�u����������k�
��E|�I�ٞ"�_��|{O�*�a�Ž�R{��$��"�6Oj!����
!�n׮�dY���C��zqs�Kۮ�m�4����?#�>w��s+�5"�7��Q�u���@g\���qE��U�sB�I����h`�X B	�f�|��_�=V�'�_ݦ��o}�X���`�ŕ�ҽYI���}C�L� ��1�k�{�����2���N�XoL�W�T%X���VeL߫غM=�5�p{@��3���\��X��>x����FG+c�竤,gW�>2�{�6��0"`[�Xu��d�� �A���Hrs}pOx ��=|^y��Z1�W֪%#� E�P��������2wE��SO�R����IyAc�Xۡ,h�m��ѵ��5g�6����?��0c�R�����%|�Eq{�Ö�A��,(�*�j��ѫ�7U-3\5�4̡Z#ǟ�Ժz�$��%u`��������)�
�{kϟ�wl���fL�,o͖խ�=/�1JA�]��/|܏D AM�uX����+\�b��
�w�H�*��SJ�U,]��rVe��{�����JUX2���"�*��Kf�w�.���W��+�SK��<	Cq"C�'�t0%7�b��s��@$w� C���Ji���M�߅Q��� �m7�#�:���6k�:��V�z��>�)����Y�[�/�5��Á3��2WF�[�I���<=��*�e^��/�������nO8�j^�?8��	N��i}4U�ʦ!j�"CM���]�t;�Sݯ�v�y�v'p��B��h擿X�+\�n�y>����g�:C�;8k����ET}�	�߶���|����#l0_Vw� �f�����>�e�������,�*����6���[X�k�fpKF�3���D�JwQ�z;��m��	�\z_�t�}�zꠄQ���bb5OZ�,f�*�M�H{}t�:�i�w=�{'��$��]7���ʝ�"M\�ŉ6#�d'�~��Z#5.�Ma�];-0]� ,AEe,�~�P�����'�/	�/�7Y��O�`��>�G�xCb��ȑ��[���֍��� ���a���h�'��	�7�8�Մ�|B�8���o�C���.�s�S��ypi��ĥ����\��}����пU�m���&��'�:��XNDB��eѽ��C���<����f�AfxIO����V3� ��nQ������n�Ò�ל�1� U��q�}�Q�l+�u��Q:�����S�%����j�a���d�jxo7]���v`g`�������t��r�@"���^o��1�i���%_�]��.1ğW��4�ڱPZ"|b$B�J�u��JJ�����sݦ�H�Ψ��hͫZ��Dy!h��6իDVK�}����Q��5�`RC;o�����:j�(L\�/a�}ߧ��P��6KD,!LO[�������2�9 "��a��(�Ԯ���ǅ��=����v�Y��Ъd�[WM@�b�>���d�2uF��D���7�0�.�Q��3 ��#%�L�.��Ŭ��N��D`ѳ��1ѕ���$�YS�u���$��˦����7�+;�➨V��,�^����.��.�1QE��U��w�;���6��Q�ק��kt_9-�k�M/,�^A
~I��aܳ�N�0sЖw�k
�5�+�_RO�ra �mwp�0���F�3�>�e�[�X�fT���Ky*��{�Fi�W��I����z�ͅ?M�����ڄK�?ŭw�bcXU+���]���@��c�67ae�1�d&sOA���):T���C�V��#�Ā��m��I�j��X4�yfN��D��5b}&���gd��dg�1��e���K
��ۊ�v�nb*c!�J�-�5j�nSŚrQ�?�PF��F�d�Ƃ9}�>~����kc������đA��U�a�>2g4�R�YQ>$���w]Ƨ�u�@c3��U�2Fss2�r�B�rӮ����6��N���.�
k�FLAQ[�<�݂:TF�?�Lٶ�v�����7�ę�Ũ���j�-�\�>�w�?��\{���u��d`�[<.������]��4��x������J:���g�5�k4 ��o����%E}��s��bA�ozW����On���bM<�.�:��$�4�B��Gfݟ^:ZCg�A�T�#��|w>-��H�������:�i���ϟ��S��裗,޾���Żj����9�
(��_v�5�nm�GM��CBP#�H5��` ��z��3�Vc�%Z�R�i�:�N�wS�y�R]7/�"ʵwa��y=�D���y�h �Iq��<J�x0<KPw �Y��V3���k�V<-��Q�/L��B�3\����f�=-����f�A�
g��Xmc�j�����[W����d=^���
��`Vዣ�$=�#SsF�*����:� a�)ʛWw�|��9o�'�U��zx��r��U�#:0�~/'�5Vl,��czT׮���"q0�k����z����W7އ(;%b���x���")��^�v"�Tԏ�2����ȸ�����k��"��ad�O�O3Ԡ6a�MG��U ]����a'�f�OT;g�۝��c�*@��y����<NzF󈁃�6��H��f�o�@"��@c
�Y�)�Nq����7D���3Է��n�N��7�%�n����g�P�(��X�WFX�3�7�w��z�Z�M���.0T���
�SGA�d�Q��M+H9� xF���[T��b�ΐ~�؆:1�f�>��1l�m:����N��#Q���.��%����Bgj�,2eC��8}֥�Q���� �+�y���Au�H�5T��@�<2�j5�(败Y�|�|�R�g̹L$.EKKP��a���
��	��0��a�AۅE�t�!;|�2�3�V���:�89�٨$�a�D;m-} ]4ŲW�v�MÛ�ڍ?�q����D��눧D����S%Jq���:g�ƻ{S/'d�X�;-Wf������`�r:���#�PQB��;?���wZ��-��� 'aC��N�o	o����#�n�C6qE��,��P)���6�jj5-rA=�v*� ]�"��)���'�M�}GD.�(�⛲�Ȫ@��f�'~b}T7�/_��c��$Z�O]�B&���ebL�'g�' �*��ĭ��W�E+�������aD �1��}��J|O.#��_����'T��[�P�����\Uc��'�Rk���=aҐqJA���Y��fh�H~�����m��ޜ�S9�
`�Z���RJ�h=�?QC�N�"S���:g�*��*;R9 �	�LT*��~�"g'��p/���|�9�uz
����negTw`��F����,��&93Xu �1� u9��e����\X��Lj�o���A�e�w��a��f1uh�Տ�'����8�N�������"��N&^���?�zN��P�s��������wt�k���D�"|�Y d�9�2����ʠH��<�2����`���[l ��J���Y� ����W��n�z��G��B�@�o�����I�y�́^��a�G���G
S��T&2�:d�P4۫$�\��㱰u�!az�:�J�ϱЙGh�J����.��4�0-�'/B�.EnJV�	Za�̑j���S�hp���:����j�+�~�a�Q�����ACg��t��|�d:�5 �$��k5��jНd/;I";<�D���X�#��D�B~�}��A���G���,�X̥dKBP��j�76&G#�ӛh����"�ל��r*������pڀ�����<퇐L��Q���j_�J�����ݺj���8�:X�ٻ�U�������35� ��?��@Fzu�fFK0���Z���qd��7�����\��Z[ �i7pK@2!M��e���k��Ԅ$k��^
�� ���g��v6���sg�L��R��;*\z-ж�^�˺gΕ�j-�S���E�X'�u����%r�<"�<��S�Ȅ�����}�޷�� ���HF*NVqV[g���#���EhfB�G�_c=���3w���C��w�yQ0�d��&�X���!rn�	3��D_���ƺsD3]s����v`Z��>�@��Pn�g�Q�j6U�^����[�(���3#��@ןSΧV�N��gg��_#-D��!��.�em�cB��IcBڢ�<m�@�w�S^d������Y��p-G�� �a�������J�Dѐ�w�F�ӵJ�D$�p���}��)wy����XA��@D�ɚ�IjlH��JF��y���7`ϟQ�ɧ�~�[�i��Q�������ʸ�IT�~��l{
��M�<p:L��З��_'�UU����":��2�yNҶTG��1��ti	B]��t�ktC��:�a;M���h���Zp���cT^�bj�'!�I5�w�3����=J�,�F}$}�wd����ǘ�G/�\�^�6x���8�Q�W��uB��BḢ%�p�	��~�]��c� ��u1�#�!�v�Ḽ]���]m#�gd1^����m�| >Ȑ����Sz��	�`�P�7�0ɖ)�^�i��e�jC\`@\dNN������	$a�0��З�ſy��VH�?��ۘ���N$���n����wX¡Ȼ;ŧ	�݋�%I�%j����aucqA��WW�-�;or�QrN��^_�,v�2Z8�b�C���T�b5�e%;�a)�٬V�;�P�(����Ҫ����lӭL~�:�aIW����?�0P�M�2�Hf}2��z("OB��D�&���ne�$��S����
��c&�������C���ܩ�*�s�~�5Q�x�������}#;^n���%=�*5�#�{:!+�ȼ�V:@ �<(`v����_nwY�=nC���SJgj�}�F���~46X�b�UP���<Pq�1».�*N#�#�?�:-�=?�&�_��DÏ��&��'�vQ���f�U,��ܵ@هz�bF?/[���d�w����c�!;[��#��
���e�r��^vX$����L	1�Z��b���B�R]�6Pf��r�{�� ��S�Oϫe8��[�g������'� ���m`���]Ѷ�0�w�����p+r�������a˿<��g8786������[���l�tk��< �%�ـ	�e� ̖U	�����J��h\ ՞�c{R�p/���OA�bgꭊ�������&���n�{,�Ӿ�-yn��zҗ fD�m�l���7b80��X��9���Bd�g�_�q��g�����/�b(�;�9���Bʙ>���E$q�
�S����5O��q]�	�7�GI�A�|�:A8i�蟚���5��[�+�9��6v�_���M8#��p(z���*U��s-o�)�\��F9�Ņ3���"ڱ��ገ Iq����$k��
�~hֈ���4�"�.�?��ɨ��,E<��ux�?�<a���+�w:�ܳ�by+���@*r�fjA�ɑ�{��V!ɧ��4�a�HkRAE��A�V��;�����X��x�� �&%���*�9��E���[��ŴxC�����#��E�n?P=n%_\����VèU�Z=&�W�8�QoR�{M���=��� [�!����N#dON�?w��ẁ��^�X0�����D�f"^��f�?E���X����4��W�RA_�b�=/�j��L�p���L���(4�}�㦪��#_���Z[��Z�����o��y;���5,6�Z�$�g4�"ur�$jZ��\�X�d�i,n�`
�(ݸ"6�>�;ZJؐb	�����|���<�.ұ/�Л�a[��*\�J.|0BԚ����U5>���� ��X?�]'��aP�*��(O��r�tq��?� ++��1�m�	F�`��?jgPk|^`hem��?u��LB5�����|�لN�<ʓF�ˠ�Їe�,�Gp+Ģÿ��c��_�P�pU�a�q�-�P~�vy�	��h�T]~�
��b$.s��sx�[ⰨŁ��	��$٨Hq1�s&oZ�3�=�GY���趢"ǫaI���l�6���c�m��Ҽ�߂�T/�A���C�W�[et�=�>�/9]��Fم����62�K�*��o駽㼤��`�/1mH�"���Gɠ�r�l�$�̄�^��~<:2�4h�\�m�g�zī����0X(�w�`��-�T�jR�'i4]���/��2��8���ΌE�5v��R��Up���fdiD�k�,A���?�$E<�/Y�Zj+'�Y��.Wwn�%W��/�C69r,$����*�����-	�� �J��XxVr�MM��b�i>-�XY<�,g}x 7ژc�"K���_dGf\�[���H�ݻɹ�q�Y:�P�p�<c� )�6V�a~��/FC��Q=�;��Gu�F�I,c��6P�Q�����	���H��s�g��NRe�A c9K��dd���p��b��?��� �E�i�O����m�U0���s��I"o}|%��V���J0!��{1��WC��=�*H1�\�Ҳ-׹�*�q��86��t%5�<vM0�*�2��<)�8&�nn�W~��]��r㹑<-�^"�}imV�ڔc%��������G�76Ӑ���Θ,C�������_�v�>�C�#�7��ƙ�QvO2��
�jP���'�=G�J��y�!���-��.����@�6�t�>)6*�i'��;I��l ���7\��`�lRzxyә���B�R�,T���Q&���|=�U�jF�W�k��
�������m�^�L���6�_�s�P>i��˘U+�X1�qn@���x;�u�b_ly �-�M`�t����|ݖ�}y�g��CrZ�wVhU߅�C^�������%�	��3&�X2��O_[J�^8<Q֬�^���@|?�4��U4H�[�vg]����
 /ou@����kp~+��s�C%���බ� EY�[�l$�}S�2�<��,jF�ԟ��F��7��w4|��wq��1������6~� ve�M���n&Y9zD����:|�zQ=#7l�����<N���{���3�i��RF�+ �f�$�nfN}���a��-�[�YQ�5Z�5 y�$�I?j�Z�.�n��WZ�X�i�h�)�H]�u���^	z�����������\�|��*���C�l�D()��̨N�_�|�Z 7�n��Ӕ]����nhv�����h���_ǃ�A�$�U� e����l�������۬Q�Vի��h��F�?���HT� JZ��6TL��
k	��j�[�/� �*�=an�45�K�j<��%}���m��A�����Z}=�.0H�u~��i"U8!���
ڜ�K��s����h����3F���`�3v��%���31v �_���nc\dS����
�����e�|v�3m��j�UD.ґ$���|2>�o�s�HF2�� T��/qV�A��o�:��Xw�Sd��j�P����na='��
Wju�Y��l���賦�LMh�n��2����iv삉+�D�iTz�|$z����|�a���x�,L]�'#�u��`�.��XsMǚ�ځ9i2^��I�����p��b�N�Z�>�jZ�ܘ�����f2i���Po�Ӧp�#!C���Oe_�/��KQ+Rm
�P��ͷoDL��ʆHM�c�U�[�+�Œ���m���p�x��� �]����-�ހ�r�d�-��K7?�w~/�#��ʐ�Ѽ�ř�D�`��e��|O�8��^��b�Im~�5@&����Y
�WkI�_5�ٞ��l}�#�Jw!�C�-��i�"�D��ؾ�./w]Y���iN��<}�#o$����@ w7�s>����-���O��(pO	�>����qOys8��]��FiS�C�X����L�>Hh�	�q��Tu�*�R�E=�����c��������`��pb_[�GZ��y�o1s�����r:�ɛ��t&��N� ����ހۧ1��IZ�^�&mwzrs������r	�{3
0��x�̈2�
x���fj����w�~ϼt��?��X��`���&e#@L�"�9�A��f����,�}�O�`d_RN�٨w�\�>��Ŕ%�B6wWqĸn΂�Y_�8Ӧ)���pg�G�SK㬪��J���,VҧMI�$jVp�8��U�d�� ���,�Z��=�r����J��V~9�|�xvU��s�D�0��aTਸ਼��a
;����\/��?p���jM�R��X����N�I�2^���J��U���;x�>+��Kc A-��{a'-xEA���)C&J��*�E�\��04������0h��M�#)s\N�F�f�0K#>e����A��}��A� ۄҩH� ���$�=�����V�~�����'��Y�Ek��Pc�ƪ�v� ̿1��
�K���P�$~?ܨ�ʙ���h�%W�F���@�?Cd�HT� SRY��P	YBk�a��4�aެ��Ir���b�/�c�Ȁ�+��aiXB���VD�i�a�N��C��+6�~|��"�R�ȴs��$��&^�9���~[�Fܞp�%X�0���Ќ�D���x2�}N2U���Xp�1@�e�i
%G�D6\��I+G��������|��j�a+Et��b�ʖ\��Mg}$q���/3H(SQ�zA.��T��-TSJ[��Vs�Aj��sS�0 ���V��"�4*�Y��+V:p��9=�D;��&�3��T�(FY�d$>�����ˆ�F�Os�4$���gXY���2&���SM~A�Tj��a��H�<����OS*���G��S-&��U�٦`�.\�:�$g���W��i�^Q�g�A���T`#`,���'�K(/����
59'-�@�f[�-~8ڦ�n��h2?�*b��X���n�!�6�>��\8�:��ب� �b��"��H���C�EA�C	B(��aW��*$ô�5��HQ%����i��X���%!�]����/��7�rޭ/�~��gc�p*�rF�>����ڒ�#����g!^��
(aѤ7T(��`�)�vQ���n�Jk��W��dpؕv>L/�_a�1��@p�g|J�W�"�A�4ɗ�,�aY
s1,R�A��J?$�laC�@綨q�@�Z^�Kk��2�eY����9Լ?pܮhDJy;xCTH�h"� ����*:)�h�7m�M��I2&�T�B������)/e
{9U[�K��\B�o�#����O 9I�)��&esj���e)���U���$ٳ��*��)F�t�=̈6G���^xw%WU��C0������7��R5�1��?�"q��^\p��A��;,V�������cy�!?�U���i6��Y��ݑ�j2��q�WTw^@J8p1h��>��-J�^=�;��v�Y�ں��qRӀ�{ q��T��K�s|��� jȧ/GfY/��#��b|�k�W�Մ�P��9,��ʪ�.��ᇬ�������Ez_�������f�1xZ��iZ�k����3�۬:Qy��x�F��!�����9z:!ǕŦ���KR%_W�n(陖�^ �Yכr� �V�F��%[s�-@�d}����EU���Pq;$�m��}��っ��4@�dQ�`��ӻr�J�Pc�x�����)�W�v����XLT�̎��O1F0T��U.��1q���#��I�@�n��>����l�ش5����9F>Η޹��N��Tm��'uօ�s?<��-g���5C*�K����I �Mx����o��L.=��,[LC|\�:�/֐w�"B��(4�öK6R���붗�+���7��x���֨w��̀s�T�	j5HV���)����$�_��&%�4.%D�-'��v�!Q�cE�,����}²�<*%��z`�%�*K�2���:���L*��%�].����I:���0�|��|��^�+$�i��O�q���ϣ��A���0%�������oF��/x{*�ֱ�A�(:Ɩ��Z/w���@�;Lw�̝�QM��`��<��:��L+�n�cmN��8�K�����-/�������S:(�Y%�&�略{�ׁ�mV ��Z���C��2��"[�Φ1�@V�G����0�A�,��_��]~��<%91�5�X9�mX�n`�Fv���a;��N��C�⑵m��6#f����ۮc��������̙?��+{i�'j��yױਣx�UK;
[��:W����9��h�$�r�(n�9*و�ME+�x>d�(������%�X�@j`n�<�C�~8���3���[",k[*��d��)wκ�����v#,�ܔ*\d��$'�2v���-G�L�Ϊ���&~��U�L,�L��#�f 9��}HAo_	='o,�~�f�<�2�D�u*A#�*x��E|��y�}j�O���/,�e���T0�F���?��?'" �߷�0��4�{��߻����09AF2@�Zi�Ir�K�ͼ)�,5�6�t<�	������_Ļ+q�u���(���[U�y$7���A�m�P���$���X�2��`��g�����`����cVb��7o���Go1_���`�N��i�JB�
"!I��mv^�K��@�V�ÆR�C�c�ml1`ׇ��Y�CK0؉9��-`�l��>���=v������^ ߵ�!{�̓���
�3�0�C�b�[��S�@\�٦�]��t�H���t�|�x:wv8@��bED�����CRҩ�b����B���>�I���_�2�sw	[�\��E�$�����|&���I���̴/�a�6��뎱{�HOM'$��� e��S��0�8q̭R�A=pNXײڝ�bR�z���ӱhY��<��T
�=�eZ���¸�\O����x$��ofn_m�I���mG����	;P�p.s*v6�x��֭0"<}����Y��>��F�
���Ȟ��cO�F~�D 3�>'럙o�$L�סR=�ޯ'6:g	nد��t�$���� �ӹ����0�]�$<��%�Z��� W�74(^�ᴷ�cIQo�Ɗ�Ϣb}~5p�L�J3?�U�Z:�2��m~��Հ�&/�G�KO~�E`HUJJ��BiY���ѣ�d������,�,�¢B� g���p����SnI:��G��K������(v����C	���<��X/̳�AN��P�����.�{X����7���D4�����b�!p��5T�|� =}���+��.����F�Ci�%�C20Hi��ލZ���N����wsH��u�*l�B�����)��IX3�+̀�[�ʫ�$S��1S�%��x�����5�ݧ4�o}&o8�"�H�KDB��a�?�n$Iײ.��S̾\>	�	Q����Jt�5�c��ul�|�(TN�
�wl�S��#���`�2B��l������O¡X@�ˠ�c��N����|XFQdE�M6eCaWӪYD+~g��P���k�U�gl��]��fa"���)r\�	Fm;�Pm����a�Rn#���)���UU��.$�����!=�����)��̉�ULr�<s�P����~S���U�m�L��-�����|���{�`q���`]%�k�� �4��ץ���Z���%0?&?{��0���u��WE+t���'��)Ńvw���%�/�R�����M�&ޠ����ύQk��g�tJ��ū7}�ҹ�9v��������M{��{�@��'�XE�,��jK	Ә�h.iqp:����V!Y��Ŭ�KA��%)��"�cLh�SD��AsLT�߇�Ρ�(�I$��z���:��*�Hh��_�i��Z��q��6�v�E:�K�n??��NP� �
���`P�E�uZ�x��2��
��0j@h���	���KE��=�F��.q�l����鉝-�c���8�DS
�􏗥����[��؛��l[�I@�'�D��p��~��A5A����~	����8z�@M��VQ�t�i���<�":�:���Q��:��%���LJN��B�߾&����:���V5�"��p1 M�1]zj�.��B\�!�n��S"B�u�i
�&��3/6_)P� ��0aV�����(۱�t��g�-��3�=PI.V'S/6�Rĥ��N�o�͹J��ƒI?xpb
_���`�[`n�Tw��:�07�:��#(�����	�M^ Q��V�.�Ig�*���\������i�ޫ-�ا��W<N�����IN�A��R�ٵC\}�&�D���#2�\���!7�%��x�8�fRm�/�8���kJxؽ��Oi��B�(�)s���i�s1���6���VQ��o�%��cy���Щ=GAf�qIƜ�OR"�6�h��q*�}�m8��j������͔(Q�h��ĤX�3f�֌�)X�r��$��5:s�;+���7��S���&�,m񪚀^' �n��DyA�˲��Ĥ�)��Ѭ3lt���b⻘�,%=_0s�$�Y�s�-\w��%Uc8c+C���%L��E��$#p�W��2�7�jU�E�O����QT ��|~*$D}�U]���vv �f�*���ݰ�Eɞ�wo'�|{��t�4%��\R�q��4Q��^\��u�mFed>��$d)�:C���8��uZD8���6I�F�5����]�&0����.� �����&�����bᡄ6�
}�` \J��Q���>%������sS<4��H&3��Av��<QՎ��Q��{���)M���,���+]R���k^���T�*�o�&��WW��v�R []�=�����|c�	�/�^�̩am����6�1��0� �sc��RS\l��7;^���}�@��[B�[���]�\m�����s>�1���r̀�'�ݶl�P� 7�u��ˤZk7�G�o��{���crn��V{��ײ�T��x�2��	\\���6Я"�`�&P��&o�V5i<�  F!�e�WJ1̀�����<J��CWA��5Z��Xe��/���]s��$9�-�L%��!L�ye�av�!�ǹ:^E@4%�X�>�������Պ
�8r�PKx���qp��Tm�:j�]���uԻ't0GM�+���<e��a�����{����S5���@�B�p���.0����{�X� c���"A��-Iw����c�*��k�mpۂ�WL�2@R;3
wtQ������K�'-��\0�O�VXg�*����i�Y�D� �U���<o�Iqk`kAw
��q��q�>G"�YіM>JXZy�B�ѵ]	R�� o�@��ϯu��=m��q��������e)�g`�����;H�\��Ӡ� �ڗ��EЋ�#'mB*����'"����� .e�"}��Y��8>�<]��#�����CP�#&�8^�_�G�d	�yβ������A.�c�!�����q���������~i��8����Q8��l��<=��p��^}g�-=�Z��ٵ�R�r�Wai�f�NR�ʍ%�˻k�ƃ��
֛3�#:3mB&}�!��knZxܵ��S��%p ���e�J�El8ޜU�Qev�1�%�N�]t���[��D�?�	;1}�h`+s'7�v����R�K�$��NP^��00g����?!�{�����4�����!�#�.[�Ϯ���$�a<�t��x9o
1DU��/�F����M����LH��~P?��UwX��2��� ��nN�����#�h�ñ����0�a�	���(�D~�`�$��⒆�%!)4ĎV�t��&b��}�Ra��}0,W�����3�Dg qL'7N�6�<�C��Q}��o��l�*�x�	s� �Ew�8X}s�<}���o�wf�(�*�A�H�,�1Cd���q�Ax����}ڍ/��j�< 9��$����6�9�oـ]���'�2���_����.t�*�c?��E�2#xM��0��3�i�l$�\^AӀsT��9�����	[q1�ڃ�����&�t�i]�4�I�,���6�2Q}��lj���j֚U����Wݰ���4Z�
�;I��}rv����`�ebM�&<�?3�;����L��tvӅH���:�D|m������p�A*S��~����OU2Z�@��;���>�lBz�����X��PM�B��#�"�N�?� $��.��Z���S^�5�tݨ����-��=o��F�)sf��WX�X��G݆n���~i�Qz�qd� ��l�ƝD�M)�Ӯ��НXf��Ƈ���l��a
ܑ3�A�l�ao>&�a�=�5'��E�3\��i��*h]r)����˕Dt���`擡�禥0<�@"�:���6�s@�	�x���T*#����@"��t����`���%1�ƘI�5N���Ru$%J�1�*���m��o4�5��A�නU[�|����dMⳝ�L��ov��u��w��2U�1�x�)}������Wu�	6��=������ �����/�*��������0W���b�0͈�^\"
����l�e'��5��P���<�����0.��#�`��`aϢ]]8�ɣ"����D�m��뿏�-9�Ñ{�x�?�����S㜸чǿOV�J~� _\����y��.m�=�!�2z9G6~vS��9}*�se@��3y]�m�"�݃!���e�F�Tl��6�����Y��vPx"�h�Տ�d��mc�h�
�B��ة��0��ѧ*�2��[gJ#�gD
#���8����c���@��$�"�7]U��C�*�1�1"X��OBV�+3�@�"��$[��V��X5:d�����cFҦpō�
އ\ uQ Bry��{w�<��G���۷"�P6��B���3�0Ӥ�Dǻ��W��lf�']eal��<���,������aV��)��+�3n��<�kC�q錚��ŨgO��ū�6i%pr6�8���;�^���F��.�L�	��aL�ް�Aʧ ���� �t+c՚נ�3�E0�튨��q$>�����(34��Jo����TY��J�9��11�n�D~�Pgp�ur��q���ڑD#q{��º�x%�?��|H�hJ�2ն��4��M�G9���$d�L~�!`�i���m&���rFd�����&2���bk�A.65
l���K;�[c_�f��`ľt��j��ȑ𱗐�j$����]/𶳘��Ew���G�����1��T�^�'�) ���s\�������,�w�d�� ��7�<���w ���I�YD�07��NQ5g�W���7�6D��1����Gl�\���]k5%�i�癃��q*^����4D������E��OJ�T9����q_4��6���w�-�*~영U4���ҠZ-_�v����+|M,�V�<�$�ňTA�h�VD�T@��X���Xb�MT	�ׇB@�U�kF���w��p��Y>�,�t1�j4N���̟j�{]�E�U�k�� ���ib
�V�a��em���H��V���(���Z���&�Ԛ���C�� 3_���Ɗ���a�,p<���*,�ep|ɐy5u*���9!�}�{-�e��1h�����9n �EV-4�6A����s}׈�&��/Ⱦ��\�C��Vi��A<V�u�y�WrO��(s^��_�9���y5Ӣ�&����� ͖_�E7�C�fm�����2ooԂ�*�g�с���(�8mHX,p�	Lx�C�)�Q�y�&���۸͢噐��l�"��M&���DTXf����M��(�"$_�^���5+���\�7t-��:�p�xأ�v������2ю���l�����Ye�R�����<���	�l�->�LT���}�(}�m۬09� Y����`ۏJ�Edu�o���1G�����XKIf`����:�p�8�a��k��HgSJ�ⶐ�)��Iߏ=���%\2Mѐ�RN���^����˶��V+�����C��IZ�_��j7x2�}w�����jט~L���+r����cնc�����n��H�!b]/%0��+ȝ{���	����kK��R�+^�����T��U�~m���:Rx�Hͣ7I?�.�"�Z��`�-_���ԏ>�����������?����0~ľx�+%�s���>&�ï���P��0�M�O4'ϝ�J�^Z{krL�:����l�Ap�T.3��&��8v�>QĶ�@E6��V�
���ZK�QL4{����˜�m��Õ�&�rm>�E;�x�3b���#��h���q`巧o\4YjρZVv��g�v���!�=H�*?򛚢d
;�.����!��!�V)�+�v���H�tӺ���\ٛ|��`��5"���LЍJ�����6������^�x���X�Z:�YZG�����q�'����6�����Jd�t��+.�r���M&�9f�ʾGJ�;������ɋ�|�P��r^]�t��t�D��hiė9���_G8<&��WQ#c���V�18c,,����T\��3�2�z�C
o��Lf���,p� m�;�0��-�.ș�j�uk���_��$�e��T��o���@�ۍu)��$�AF1"ڤ�Eg�}TRx��?�P�3�Ѻ�o}��*6�[�b�@ƕ+��2}�i8i��G ��aD]8�IkGU�o@t���O�!��72b�+n8���/�T:�D�:upW!&�%M��T섄#�5i�_O��T��@�I$dw�dlj�|����L����Ђ�����6 ���UĠK�`+��X��L��V���[�չ��T�*��G��1I��O�u0����7*�nT�$"�t�yD}����S���̟MoǛʸ�S.��6�H���f�����᳗�V�O�"{~Uo�/�s��y%Y���{��6����@CxH�'��7��N�Z%�}���p�S��+{��;���ݧn�����;קalY?�4�$	Jv�N�ً&��L�l7}]CJí��ч����0|ݳ����4(G�0A7��ق,vp�z�0�΅�J7W��O�f� ��I@4%��4���	��S��2d�n����&�b#�(���7Su3Wi�\�@�/-�C���=��tL�h��C�d�o?KN��.;s~�7�\3�˳�c`#��㼴m�+���ʙ�k\��Frj	���U��]����ƚ4��dޜ�=H�N��D��vnz����"��s�T�ޢ���l���-Ę� ���t��ʩ_�Gn6�H��cC;Ŧ6�:~U#�r�'� [f�m5��q�AE��]�|uʺ�b�\߻����fX��6+??�T?W�z�֦��;5a�T�U��a�^za
�'���wO��}�q�KԖ��Q#�=�|��
��bQ�4IH���3cW����7�'�I�t�ե�ޜ�V黳oʖ��q [wr?�� �^k���>w����v�ʫR� "i�"8�u��o*@��ͱ�\�b��zF�Կ24AD�,b]�><��K,<�O:j���R��CO�r,�ݘ�	��侊&6k~H�${T)�N���;^���m��;���LY5�l�6Y�F.��-�xc�K.�ޞ��O��m�Ӷ���C���RJ���4FgO��[��:y�ҕ�ÃD��A�a<����a=7A�₩=e���S��������+� [C���刜R��mR3�W��Ca��hM�)�Q��L9��ϋ�Jm}Az5%�e���-u�'d��y7g9�Sq�$�Xo%�J���N%gҜj#��g0�^��|vڡG.Z;0e�Q���7�ݑ�e��W���'����1~��G�ppS�-��·i��	�d�'$5���������ᙥ�z�$�*2륩�|���9���C�uD��C�x˓�
5��i9dI�����c�0�W���B[��Gny�\(0q�/���H[�F-J�K�xƱ7�R$��K�$��ď8�N�6 �q���Ո(M�]{\������pY�v�@������m������C�(��xR�Mh�����"�'����p<��r8��j���g;>��Gf�����J/�e�4��)UJ���{���S�G�v�LSDeͨ\��;�Cq�b����n'@cjNN��?�]B�>��L�t�'��;��}�VD��P��(��c���{�iK�=*���.]��Y��2���I�H5�Y�D�w |=�%�D࠳�'��K$��x�8��RyLN��hz*d��LB�e=�_T�$Ȼ�T��Z���21����ʔG��["?��]H����HL�ؙ��B���p*Y�Q���N�I�б���GT�������$�K��o���(hw5�6ZBO�W�=�U|sn�(��RR�u|��Rd�[!ϡ�����Z���m�K�>�+ZwU��?� Y�&�³��(����]���X�{Axt|����<����T��R w�釰��*)@�jp�2c�$���դ���a&uD>�u ��X��!���E{Z4�Qj�,ZPB\��<�u®�4� �˪У��_a_��8�
�������e�`��� 
Oa`����e��w�d�]�RbI��Z�F���_g����h<?0�?���O�O���tT����է��]��j'z��>���[ȏ]
n�乐0�8Am(/]�).t�Y�(��@���
Z��l<��zMi�ο�|�_@+�M���0�-2�y^[F�Ͻ�G%��g	Bb�BJ�HQ.�dG[��x�QDm�)+х�n�s���,�o��2�Fo���X��[f}e��~���z���J:�K[�Z���5��b���xYA�$����zmxd�qǶ��s������ZD�Uwn��w�HI�mB`V|,��ݫqlՁ:�x8#
p�-2bL���y LD�����!1B�/tzzCV����a4f�ql�Mk����'d��)8c�4�SkKK�B�I�,�6�c.��P	>Nm�^O�>�
�}%A��<Ť���ί5�A|�j绳�k�W�YҭBܔe/mZ����Vx�p-�I�����:�uc�ev�>�����I����d7`8���K)�����ʣp�� #[ 8y����Ž��B���=P��c���!P�ή�*��.���U�9�޺a�ҊD��W��]��d�����*��҅=k��>a �P��UL_��b�l& 	lR5�W���p/�q���a�����`m7�8A�[iW02����2���B��C��*葱�{��v[������լI'�Ӯn�9K���+�F�6 1O�SiV�h�H/8A�z�䄖��.S�� �?��Hlx��Ou���e�����DC�(�zPѾ�g����]�^e�`�ood\�J周m�kƱ��S9ۏ9Y��ivwrî]��:�q2�Β�RڟO+�>��s�������?5��d ��C&V�g�D�%�8k>y1���]�zl�}���#�D��H���v������v�R�鼺J���~x�]Y�^s
\P�^����Ky#Z��a�n}#��L��i�����F9��(��ؖ�z�p@��'D�v3��uC�7E��17L���\X�u$�K�����~O=��U��͂Sv�I�4�����vg�w�П��1MD����AB�6�u�%0��AD�hgzՏ�������$���0�N}�rO
�L��fMXu�-�O�* �}�|���� �33�j<�:���� �n�{����N-�gg�Z���{9�|Ͻ����6,��k�Ǣir��0���%����p�2t�ܭ���zQ�]r���:;Eu�D�i��M#�Y�M��3Fu��Q��F�L\���>ʘ���h.٦s?�$���Ob��<R#�'�|�/s6J�������f��xAf/�㠤,۪[�Q����Y�*�Hx��"e(�c���B��m��t,+V��{E£���U�O6?N��.\��p<�<æ�G���J�U!˺lB%>u����B�����.�%��-�����R�(�Y�*�h�򚥴a�܈+����p"��a`U���w�zo^ ��8 ��E�P>fn-2�G��a*�l>�	�"o�P4Jr1�r�Y7��B6����'�bGS��x"~�FU��n�rv��d#WB��*�u{�jb�,�5Fx��IP�!��;T[�f	Lf4�?������Z�� �mm��"�|V�4S��Ǔ�9�5�u�.f�l����T��n����������Ki��j��4pM�ͨ��R<W}�Z�K��[j�6�(k�ǘ�~���h�S�ާc��7;�ɢ{�G���>W�/���vۥ���h��:�󠕻 ��x���veE�@���#��Q;��b�v�^XPV�e��V<����e⿹
k7ș�:�Nz����kLX"�h��z(���w#F�E0Ex���M��*.�0��厅lə9e���y���WǕ#č�H}N�G�Ц��v��ew%�+��k��w�P����x
�]��s[|�;�j�sFq^,��r$ 
��͓Έ�9
�궥����1A��g����6��(Wa8Q��|P��ByՠD7�t�](-IB��T�OK��´���TMg_��p�R��L�W%���m��=�.�ͨ%^TS��� ���.m�Gw!�ߢ5 ����W�!z�z��D�{�5>�o���2[�P��q-Tw�V�Bg�Š}Sw �5�rTH�f�BwY�A�/�U�z�����1Un��x�e�|Y�E�]-P�+�����ǀ'�\$u�SX��:d��[�^��3�i�%���A)��H`_��*�܉ G�4��4��w�c��ܱ������!B�OF�umP%��NW�2���W�����}�M���v7\�Q��)�z���d �9ѳ!H0D�I�L�W�4V���Z�kLuܲ����OEB�8j�N�]ꭖ�p�+?����l15.����`��}|��ٶ���r�:'6��敕�!{dXy�)���v�f�w�dXc~~EC݋;㚃JA�7@l4��N��
jl����a n�h#��Y�`R�T�a��c���8���MP^��� C �'�^T/���ӷ�Ox8�
�M*���/Ц�P�,�Z�Rs�Kj^�1<�,��P��K������N2�_�k�����E��9�A�
�ǋ~n6_�y�-�?�&'Pd�UR%��z-�ě@��!I�#Ű�³傱Q�!���Z���7�Y�(��]����۸݉
a���hoMb��h�B�"�>`-Q��������Ǥr
}��:�,Z���^�qD�p��b �? ��(�
"���l�l�Bzx޾6U,��zL��p���ƮF̎ ���z��jKl~=���"�<w���+̛V@�4���\'�Y6@��?��^I��4U��A�q��ukr!e��gCO��a���wy���v2۟ܜ��^�j���C����!@>kuޅ��]Ҹ�%��b��i���\8^����{T=Ύ֒S�zO�}e��o���}��uz�V�|����ֶ���>2�dLx2�ig6�+G�x /�O�D�����Ui:�����<���Yl��Cbq�T��s�ZY��s�p�c�s7�L��WG�_@�aC�hnD���J�JJ�	G��i!����I�����F�[~g��"�U��˪�q�F?
Y�y@h�^b�07@��3�?�9�*������3C�p-�3�}��+�s��������:VD\hA�G�<��֨��w=�}&P8��j��۩���c���������hp�a1@��2!"��f{��~�.5��D�lX� V����Pm,�^Dc.?��tj��89�|�/䛥RJ��*�s\ϛ]���ڋ��Z�@�vXgCW��-��p?3���;yeK���3W����B�+Ns��KY[ >/���$��`��������E�u&U�wm-Apn	O��:��6���}�a�{u��Ф}���F'�0`p����nD��;v:�ծ�Tos�B�,���0�zha��)�(ԏ7G��	�G��K�&q�/�p����</�T�Z��B�<�4�c3�T�7��}���y|gO��G�WBFs>�T�!z�����綹�F���h���1P�a���M<��f�okk�ȭ9:����4��evdz�b��T[����X7�IO�B:W�5��G�U�L�`�A=��X����W3����$�C�A}U�Cwj��/�|�0ة���G����Ff!w�e=�5G7��J�(g���x�3�����7��'Ü�G���u�l)Ը�ɧ	f�2x�2�i�����j�~ŭj�E���9���Hٵz�j8gh�I���5��3�y�Xɖ�*.�髇:�������:.���'��-�ՓFeU�HX�m�D�X�I]�1Ҋ�BF�s\��!�BoN�;���)B�BI�g��jj-,��5o)��ĻCtk��z�`�s�lW|���ذ�/�	:��������eh!��������f�:mT��+��3��Ԩ�
W�h��@_���ò�Gٱ�c��;8w�h�_�R��{͐[�D%+�����f��q�n����˓�/躁獚�;<`��6f�����
������q<�;^4���0G�ɬ��������7U9�n�|_�QL�dI������ &��u��z6e˂�3�^����°��D�c:O��fW8K8Xv��>b+��RnI]Kcd@�4�G� i!s�hT_4�zZխ|��&1`�r��fvNW���,�Ԑ��~Ms�#����T# ��G-R&G�N����ɿ���P�H���4�P�Y1ŷq э�\����֘�� ��F�$}��?-f�{/)7љ���х����"X�N�@+�,,���iP��7��ټK�mp�?��"OZai4������^]"��u��H�X�,�
�$��S���|�^W|���-e0� k�Q��k��Mx�9�Lu�Iz=�00�#���{��H!�ѩ'K�]M~��BTZ�r�Ӵ�v���V�l����P�rpS�{S�j��d[�V������?���>�ɣv|�`�E��I�*o�%R�y��8����\�C�y7�)����HM�+���"�ά�?3bC���;�:K��aܙ#2�ю7�T���=�����*�g����nS���)�֓x}(����X��j��ı��p�����0%��~n<��	�1�Q��C�p�^2Vz/�Hp6�D�l<��S�Թ��6-nu��l�9�
rro�]�o���UlY�`Sk�kL�/�מ�{;·_ѡ�S	���G�`Ҩq�i��|Td��m�\_L�.��m��]��[��Iٖy��M{��ګ���͗`8N/���I�	F�� `�M�O�r�N���� �Y=<���Z=�}#�݅� ��Ii�F-��z�r2�c�
��wM�Zl��2I![F�S$�K,�/�{��S��mr+��_-�BٍT;>�����'�� 4� 1�{ԧ�@��:�2Y�%�x�&n�b��hiD�Jnӣ��+��:�/�60<�iC���Ї&���W�!u�S����$��KDI�6X�F�����LV���VNrj���Uz��n����y�,��望���~Z���y2��61щ	w���L��L�E*'�ц=89�gKE�J"����)�G[���K��5S�6|N�0 c���Q/��}�ta��F�1�8���Q�z�K�`�&?S����?Yh_��G���4ݑI �Gz�n��ȭ>�t,�U��L�.j��sX�\�����+<Jl����r��y�ҝ9����5��g0S`��vϱ�� Z�}&��ϛ*���O!�F��s��t�8��Ot,D%��*j~ٛ~�K�S��2�Β��'J�H���g�6 $��ޭ����������L�uY �L��W�~�8j:���;շ�|�I_���G𪂃@�#�B1,�pu����>����,#�7�F�& kBN~�V,�$��P�W�גf����"v�`�Ч1�j��]k�w+�� ���[�b�fm#�X���ZH��	�*Ia��X��h��h��ٔ�k`
[�܅���t
��UxԲK�����ԓ�3��A�k��Z�Q9pd��܆��ױJ3��ـ�H7�jE�����_�6`�*v�2��9`��7�ݲ�\�_�~vo7g��ӟG��-���5=䀨���.W�G�̆����>����	�'�-�Ƥ|)�hZ|H�!º�G�`1ጔ��(9���/K���:삂N4�&���u������j�)r��\�֎���z�[jU��k�z�x~N�������}�/(��<L��}�-{�}LuRjɞ��2�졅n�����w�2��@YUcʠQ�3�T�ʈ��e�jv���5���V��l����� ����:���L�s-i�\�W%�)����ˮ�y���ȞA��9o�����)�F�Q�SP���;�+'b�{�q�n�-z���Ÿ��ŕ�'69���B~�s��(L�����0��g��Z��I�W;�s�C���,V��:9i,۲H0�m\���Fhء��AR�W;���	� 9
�:b/��e��UI�B 1�<� 7�Pʐ���G���}�����;�X��-��v��$�Kؐ���/��H
a�(M�&O�][ۙ T��-�/Ĭ�p��0��!����\t\R��Cǁ���*��%Լ��NX�������}@�n�h$����9`�o�Y�!�=|��IL9#r���%��N�lSn��c���TX��@Q�a��o� $����7U幩�3ש��l״=��lF����ȡ,�趻����z����*�F s
/L��sc�:a�-I4�,y6��c-����̈6��p�DH�s�*�)dQ�Q&*�6�h��b�a����$0���	_-�8��'h��a6xX�S����>���0�`���]�� ����	��}� ���B�=�������$���j�(��4W�@5����A����Nt��r�k�G{
ZJU������&ҩO�k�/�P�!��+[/�ȭ�Gtd�����ͳ&[�OBc	�H�!��ͻq��q�Zh�G%rY_qM�#}�b����0^����df9�j�)Pg�F.��"nI������,�+���/�4mۜ�.`�ңU�{7�(�á�Ԑ���EW&cR����B��|c"xH�y&�%���v|����r� ��8rL?^t�M��ܘ��Y�:u�������2�k����j�[��g�����m#7���(<�)l�(����m��Iqj>8W������|�n)��r, �'1��$Ҳ	Òq�Se��_
�n��rrNh����td��)��M�)�V�/�3:�s\q�P�?�~��&I>6QQ+dvn���-�$�#e�ث�Y!c+7��?�H{؁�fv�ńߪ&s�K��Gx"|G�T�GI���Ua�=�iƩ+u�9P��ŚM�����0�	E�L�5I w[���pJ֤������0&��6V �Y�d^��{�}�%�����IDq}0L"��qK�u�|b�Y6�,}������������T�84TUo��o��Z'IWz������_q�(�'ma�˔��u˯�(��)Y�f?R��z] G7	�܃$ϐv�w�n.?6��L�2U-��mZ���ֵV��w@B�e�Ճ뾩A��c�+wP�[6���Z�n����a$��<�Z����HݍL������Тv���!$>Z⢹u�'�
��vy׌��[lA�N�B�E�L����ߕg}֖��W���~�bK�vn���4��k(��|��m:G�!O�h��k�4j@Q�� "�q�U��Ւ�D�X�ة�*Vå�k[O�Z�lw���k�x�~�W��>t��H��hC��s�qr��������̜|�(R�_��O��|z������fШ����L^ ��7�h�v[B�l�hR��F���A׉���]��O�m��fۿ�Un���5W�-}nk�G����lh�O��C���F��o޹��H4s���E:�޶=��c*Co0 o����{�}"�0R�4� �RyqA��T��(����m庪��Kz��h��[6d����֏}�^-�� ���P��MXgߚs�L�$D����}o�(C-Z<fg6�Jg�>�����tLq��LMiS[���At'@��5Xz`6��ݰ]�%efl֋�p��r'� �T��;G4_O}�j��xw�����S�x-���sSx�:
^��~�pd-�@t��_;�	ӂ�ƹ�E^�H���az3��z��ِ�LȽ�7����#ȟH�^������G'�#^�cǊPӴ�m���"����C�[k�
��)���'��3�훗���*�I'����ϯ����o7�C=xbHp3O*��?������T���Ԙ�NO��W2/?��y!dH�ؐ���^�~�<Ic���@y�_[m{Z[(�inJ�<:��*X��"���-,}C�vnp�b2����$S�����&Sf�T��\Q�5+�^�	B�(2>�K\��u2���4s���\fT\�	?}��8~��b9��&��L��,h�1��QF�r�s
w�n�}�Z&-}u;p��i�y��$��^���*u!ډ�	<��!�{�p%{r�-� 9�3���������}q�i<�KP,�XY��W�?[��n����(F��Bч��*^?�#��*߄�
���(��~�������m)�R��j��jhZ�.ӂ�m`wm6s5C���(�p�z��R2��(,�gqY�d7�D�g��G��H����>�2�A=��bZ$xF�G4�Qm��mL�CT��f���mq݅���*��Cl�)D1BX�������V�Ia��!�H8��U�$d��Ye����ڑ�Bŀ�mJ�!�%52�;���5�ڋ;��?��F�.m�p�i��Z�IH�Z�Z�@]a̪�]�	�.��C����C���T<_�-n&q�2<���	ޛ�o�g0�r�Ї}:������ ��tX��I .{�����{~E��H\lŐ�l��Q�����c�vZ�
IƱ���16���=�:&걦\���� �Wڽ��7�9�/kp�V��;�&�e&�i��	Kf�5aE	�'1��W�a��!tl�"�\V2�2y�*��� v�q�e���Hن�z��.Aќ���3w�������Ɏ#�S�e�
��s�p' ����ĆB��ԚF�(���V�p��p�23����*/*����M�J�����fx���<`Ht%��ktC�c��H�+�p(���d��B۞~,�{%�9գ�x�!�/<�ߞD莥����I"V0�>�b>҄�Ы��R�����/p��n�N��vL�f@�Y>� �֛"M��lԖ�Q�BD�ֵ$ʬ�<�{����&���]�!�̃��s���u린z#� �	i`���KİR�5�e��s�����W)�E�̏0�n�8�:A�5�/�Y��9~7�n�տ�a��Bŝd��O�P[H��5Pw|��-�6��5wZ��?�cH�]��;��S�R�����_`�Nm黜Y�������F�ة"�5۽I��I7���$<����7]��܍O2�m�<Z�c��S0Fmp�?�wS����&�Ay��7=̎G$x衈J�vu�Ps�R�I����n�b2ZG#-$���Mm�5O_w�tZ��L��}VWg��Ak��̋pS&�fc��&f�yLh@����eEܪF<V}[S\'�$�0:����zGI��~kI~���'x-̯��x��׹�st˲i�%V[VC���[R���_�U(cE(��}x���؇$� ��`��V�?r�'�l
n�YA6�|I!����/h�h��T� �f��}��b>����wu�+���oz.�m�B�z�Sy��Ѭ��e�:�G"X�Q�#�:���S�<f��e6rY�Y$H�4�����	�^��A2`����3PE�G�Q�V{����ř���bX�O
u��.;�)��Y����1�ԭ��W�6�=(li�U�)�^�s'D���� )06%) a��,�����D�ClK4Gɐ	�y`�e�Q/p�����;d�N��!PmE e�}�,&��Q�2�zC��ӊ�-���B'3� 	~���\z���T��R��`��)'ڃ�'����Iz�[o�Q�н3%�������<��^svE��9ן����)~�*���^nZ�_M�/	���a�DM����A�YL��O@s��rp�dg<�m��R�)�X�ה{���HL�%��(:i=� ��{pp���*jS���Ѫ:�4:�ܻ���2���Dr.�)0^��fo��i��u�ʰ��iTԷ��ϗ���K��| �鸉�X�->�TP[���-ـv���=,�ͫ+2�X����O4c�����N���,G)d��I�7��e!�j����%�a�_����Y���&�B���`��gjYZ����V~,.L�u_�G�%��BA��d]�	(�j ��|���Ue�ž%�����@{�ꓘ�!aC�����tX�"4\Hc)�H�Nt}ۅ�cZ}�0�����K��d�|��%�R�%M�
F刟�l�(���)r/E�4��u��+S����#������L��T�@�"�����Q^��Ӂrt$� �w�y$��*Q2u>�2�4�W����ϟ�Bx�B(�7Ҩ2��D91�CJ�]�P믄���ݦ�C��\1��K�Oгvg1ܗ_v�uqT�7���ļ�*zG#�6W�c4~'�_ҹ/u��艄m١�� ~�9�o�S ��P�:�3�h>�9�[=1Aj��"2{F�����xW�t���(�*@F|)=!I)7��f-jS���s�a|�Vq-�Uon%�2V'"���3A�~��@,�	�n������8I��>]Y� t07���F8?��/���DEt�����T��$�l���4'���q�#��.R
�0�+g;���KW8e��u���-���ӏtȒHe,�nh�����r1����� _�l�I���Q���?��#b�
����Tm��/Q�;��:z��}fl}G�{��鯽K���y ���έ��L徖7(� ��h�C�S��H<rLG�[4O��*v%��cGޯ�?�(��	���C�1��q�-&߱�uX�bݼڳm��4c~E�����N��9��q�h0�c�R?��&،�׍�Q�*k�:a�U�$���s��`ÌC�9 �(d�y��j�%hw�3q7ci�HZ��{��E�E-�+ ���;Qq�j���e2�J��!)�Et�$*���^����ɳI�C��P�y�q �W��ȡmDy3QPƕT"76>��A�^�qX�j0ߔ�U��{q&|v�YuRt�		Z��#�t#TV��#BaM��w(�ODֈ��A|�I4g��d;�4�#2��/C\�QT��R���.��5v�b:Y�`�(���K3|�x��N��A�ǯ �$����4�يa� �����h�s!_ލP�Ó�=�F?��TuohL�8���Ʒ�B�\"�c�?1�}��"��}��,��p��9�V�A��<�j�4k���hL{oQ%r�T P?'���s�v:$��\,����]����D�H�i0Ĩ��Z؆�(?- d�!�~�̆<����	�r>4��boNn-�|_�2����郰�.��l ;1)_��*���9A��(�(�-!P��F��w��M��c��z��|�%�yN�,��O	�N�)5��_s���ߴ��H��?����_9��a�br���2MX����2��,'/�%rЗ�-]�J��!W�6��k�)���ON���C�_x���
5��iK͙A��IR�/����9��+�� ��@�_�Sv7ԱS�ɜb�I(���p��u\�[��i'�L��$SJ)�	[�p�@RM)\D}���&/J$�ġ��i�rY�D*BkE·���V���s�-����u�S�G�\�#���{	g���A�1�����ȣ}�u�Ҭ%�*���J��"�yy��� �	�i5���r�*�����c��w��@4#a�N%��#�V��NG������\����vg�^n��i��R���ŗ����q��C���t!�$|�dD�0��2��N׍,Sy���R��V��&/�P&��;N����{�z��ޘ��
z^����%�(�f6�h�򤱳8t�����_�������A����l���܉Ji� �*��U�hwA�֠�_MP���Y ����P	�:g]�4(�� o랏bC�Q҉j4��'md�v����73�����o)\ȩ��d�E�Y�9<�b	��)�&�f�=�c`�JXr�N��s���۝�j!���Ym.@��o'TU s�����{�"b��?t����Qñ���q�r���64�?�(G��U��yU��>�s�NϩH9�-���$��*��Zj�Th��i}�S˄t���"��ͲD#򕨸F)�*�cң�D��������\	���~w�kӅĤ?�4��,4��\Q(��I��t5��=�V6S4�[e =L���@��Ok�+`eH`��y��2�i�Zg61YެY>P�7�>RxK�_id��ya��o�AMa���L,���wF��`���c��|��}Mp�h�
s8�ƙ����w�4�XF�I�73�.Q���͍`7y���ș-q�il��[9F�/Ӂ���'Ee�
7L�x��'L��r�4����l�@ɢ<=���y��Wfy�#�����-��}%~�!+!��;)�I��%�xȵs�����d6����G�^��c��S����z}3�x ��+��g°M��p�9y4����fj�����5��KEx�ⶰ�pw�߬��+e�"1���N�����^`.3?&Bpl����3�����ݖ��)�en��n9M:;� ��:����V�1�Bx��.7�-�ٟ�'��,PC�,���`0���i�`�]�������C%���I�fM���݌y�U{_�a�N��Q|�vMq%}V�=(�T*.�����b�[#ƚ���r����_!!�o��=[�	����v|�m<ђ�������� ��-0x�g�B��0��'�c�Ϣ)�Xخh�"�?M��+�z�:Pl2�~�i�?��~��; �ٜ�ՍQ�oKB�LA�$�1��icZVOd&^�s������͓�9��=JGpb�Z��;�Z#x�ŌX��73�"d�#�U(�d���&���`I��T������9l�ᾑ�\�����(��v�O��"����j
�%/�`m��m�r��P@xl�a�Y'�u�+�����$�LK}]��߳h�@Q���L_��?�ـ�R�4�5��oȯJM���7�|}�:�z������D�L�DI%��i,$*Z��T�#,�Cg20�}�����t�W�9ݞ|�M-����/��(��i�; ��u���l��c{����REH?�/�	9ঔe�Io�L���[��B��D����}����jH��(�9/���p�B|'0^Hl���tZȍ�,�X5�����[��p���Q�- v��B�?�9���˞���+��C��/������+���1{�k��#z�+����	-��4hCmu��g+s`Ǯ��H�}�Nr�׋��E��h��o%8H��xy�|�,�k��wvh��"u�j{(��oi��q���G��xs��l(���Ӫ:�s���JѡӀ��>�hm`�wܺ�W�vw���H�fTX���O7��R!x������͕������ߧ��������X;r�T(�sS���2%�f��b1��\����"t�jDݒ�^��١�}
���]O�+���ǕE�g�+��K*:��^C�EpJ����Fic��&/	.�:�Tj3���;���NVT6YH`��F�f,bi��/��_���W�����c���(�n�+������3M��#B�g;qij�A����*�w��"a��������ps.u<k(aVA
bz�� ��W\�p��;����>�	�q���mH؝ޠ ݕ�!����.U�V�d�}<�.x�Iu�dH�2`)qn�I����P/L�D)=��u-Ye���dY=R�	U�	[Ѓ�0ܰ(�a`���/@�rBN��A�/��Ȉj�|W#)��d�1�"L�Up����-%��/�[*Cd!����b��N��5Ph��p�U[���k�,wzٶ!���$Z&u�p��Z;R�C�{�.�avc���j��*�,K���{c4�Q�y�I�(0��{��]*.�Q#�C��Rٌ[����ʚ��qЧəj��-�TO�l��~aª�r6�98��+��/�����2��_�I���
1���с�F��lfpa��P����ym���m$1b���S�Q	S2�q�϶z��|
1�ާ�>��lf���Sp_��Hy`�b?��l¸U�'R��e?\�?j��m��/��������#U���X�z�J(^��TB��`ɛNp9��S⋩�����/Lk��`l��m�Ϸ��Yu�%��<��ϛ��C|�]�;�]�oE��q��!�ԵJ��t-9��i��������V�����xN��NV��'�L�e�%Z�3d{��0���T�nY�$$����ա�%��{w�1f���Z]]��X�q��Q:U��H���e��N䕭�B�}����n
�Y�9�Y�$c��6�s�l�7$Ւ+�B�H\3�")�I�����Z>,��;Ua��A]t�d�wc���ۅ��0V�8]���Ĥ�v}�]�{7h��Q_B{\����?�N����I`̶Y����P���,�HDG��d�u��u�4��v@K1�����_��i��ʳԁ�r���'}��� �:�K�y��z'����䥲�`�v>��Oɫh�ֵ�o1,��5y��j��ˆ>Ӿ�ۤ���+at���8�s~s�U%gHB'�hBl����=#UP͡��!:g�8���l ���{_�B��vQ���j"�*g����{5��\�
�H���!����� e���e����-9U����m�-ӵ�E�rڙ�3������~�A6m�uԾ�oDغ��1o�a�% Z޹�7�M�i��8�v?n���tE�����w�SE�>n�B����X�iq���6~&UqFR��ׄ��A�KX��Y��h����<L�Xۚ�I�v�j��*m���'������v��WuNZ}��Դ)�j3&�l� ��d���_�_=>g%&U_\~΋���W�]�)@��0��VԦ��{�q� /e/N�QLV!��)J���2���+/F�`2�9a�?���:Ȁ�Kb�i�"v��|�	0�ߐ�׹m:��-H�&����q/�mڰ�� �J:X'�yS�~jm�gqD�f�������3^/�Ӿ������������!� ���LAsc�Ȱ7�s�u��
P9J:5�I_]j���$�w@ڹ ������d90�������>,!@�h�w����svj�j�0�WS�x��x]35+�D���l�"��~�5g;h8� ��o��m�̘%������GL����9{[ ��x���E���D`��{��o�*8�j�/'b�����٤���h�>�MҺ��;&�O��)<^�l[�9��(l��)���� �A��	�o���`R�j��-˟,z�Sݣ�T<�z����t$o;�/���@�g�6C���ۡ7"+���1)hs�AI@�z$�ZD�5Lr�6L_:˗M�����
�;5łiN_�3�e��|�p�~��#E�v{��Eޤ�>ǿ�1��b$�[�U�Ռ!(P�jz��c��Ż��V�U�<0�˚Bm�n�zG8��XS�mda��P?x^��&�q!?PL��P͖[Z���9�es22�'BHڤ�n�Q�������ٮ�ax�F*�v�m���) �<�(mߌ��2��[�fO�	+A�{5�8\%N�H�S%�'��[���T���:һm�S?l��#L�W�x���R�)�&u�σ��ӥ�~�b4����g��s\�3�h�8�pu�Fu����GV]��+x�o��f��Βo�N�����P�i���j9�}1q�K).���&籸��|6���VoU�l(0����g`�� �ѲI�{B�P���a����4�䇩�!��a~�+��]��%����W��]���x���(M���u�@��4�ΓY׍�3�y6>3HJRX�,ɣ����I]��ՕH|�����u��\r�Q|z��҉�G��Z+�¡�����γ�#L'!ث
���~hs��,�ݼB#Iᖧ��i}أ�w2���˽¿S��Qt_�q��D���HY��'ٷ�<Ƥ.��$����}Q����S�o�`f��0M���-ce:����!v9,��/e��5��N��_�6�	� ؈� ��ܢ�!0�}�E7Y�@��@��*Y�=��=^��4��
��E��E�P�@�y�W�F�t�>N�H�ր�_����PJ)u0�mbl,�M%��s�r��tQ��t�5�6�M�ەB�/�ac>$����{��;���b�_��0�E��B�Oי��f��$82,����<���="���[^��;��)�d��{��������<�_�Z���(������VzU���Ss5Ӧ��ru�O��i1�H��hF/���4��YY�HՕ?�>G�hz>`T�2B4?�I��?߁x��.���m6�6�7}�ϧ��޳$ŉ��
�E7�VnؾH��F\Έ�NΘ,ҵ�W�9OZX�얗���(�x3gZ�L��W�43u)����󰺿�+����ӆB��s��s �J.��& �f�3#S�]_� �$|�":v�)��ջ�0l�xl9A�T�C=(,�8*������C���?����ͷ��E'	,��x��y䰗�i֕aa/� �y'V���:��(�M�N��$���1���n&�x�y	����H�<�*?��}�>{�v@�w7�X2��U�M����#
���䎛�Nn�U ��H�C9��������Y�
�gxaڶU�P�T�"����u��>��>�����f�Y"f���d?�������3�]�0�h>$��a�L��p�(����R�-m���%R��m����l � D_
�9܄�܁
��12r֢��B�$Eq��[�2�mgtf�jr�B�WW��w<�t͏��Q��
k�v�\O�;�J�R۫'�a��%sO�)r������	�nh򄋘y��:��"7�r,o�����mcL�@�0n�j��H����e2{��Z0H����[tE�gU�|ܔ���ਜ��|�������M�z�
Ј�eqC1�T��+<�a�b޳���ʡ,^:4��X�j��&=�J)��h#�msp�[*n��@��S�!Q��I�I߯����o��9�`8*-b�ϟ�vX�1}�'�z�#L6P���Nkq5�O�k�������@������\(ٝ0�ZE0|d+="6������+�.R���f�����J6k��ɑT-�9�&�=5V��ڭ]�
�������5�U����L�H���!��c��)��������C���_�x�	�Ijc���9����͇jQ{0���P�ҙ]eA%�!e1�3Uv��@�H j�(}�J�)|�BD��w���K��9IS߁��nv�i�T��1.�h�V�����+Pv����c�I�;+R�������)����L���'(J@3}�!Ő*��J,�{�� ��`S>�ZTb����qSD~�j��x�@�;��\S�����|O�-�&1G.#I�ܡ���/hB�Z��<���$�	�c]߾���|��`�2�1����P]�#a��Q���';�0
+P�Շ0O�zO��E8�������VP�a�B
/$RyBp��J7H�zJ�E�xg�0J���|��l������-�y64�w�=��f8
4�	�u��e���5 �4c�M�vm����5�D�-�۽�IdU�ש	�Y��a�ŝ||Y���d�
��	�t
h�2k.P唺�''!W�PNb[��^�^۳H,=�"{(���`���)i��E��ڣ�*��xc�ֽ�e���~�M,���/�y�SL�+ۉ/G�j//�g�R�k;�6���$�B4�^t���y6:?
9U'��Mu{EVTz��]����4`\6��m?�:X����9�����V�^�Q��^�=���7����9�'��Iطm/Z9���+����-q�v�t�В%�h�w�mD��;wm;Y���Y:�5vzz(�w6D����؎8�$��Y	�w!9Yϭe��W���6a`�����豾�0�Tdr�Z���� r�N��ҩ�*���V�t�s`Z۟����0��_}~���?��hH��/��wi���XúMQ���������QAQ��/��]@D��R�4�Z�7�R����C%Pq�)�#�P�����x����t�����EV�@��p���.X����t�
;2�^!"~�@	���s�OV��~�/�!	�r-��x�`��9@�Z�1Õ��o S��rxPEM��}�?�x�lH�n1c�0U��]��!�0X���\+�����I{7.�E.��V����)m�5���Y-øS���{�#�l�P>Cr�>�+�� �V�֟(3	�g���f���䦅�(V��L�7�4���I�YR�.68��h�3����On�Pŭ�jAp��F�*�u�\�8�p�a��QN�)��{��A⩚t;c]:,��VD��Պ#��VOs����{I3E�p>����Wf�s�~Uܥ�!(��~i@���ly)TN��g_��N}(��2��;-Z�=�5+�n�܇&]B�D�p�W�0f��بn��P�ʯ�R�����D 8��v���8��A�f�{߄ m��y�D��08�{<�Lg"屵%�qp}+���|�'�d�bʷNe.(]�	���SPU9�O)z�cr�<�0f�o ��N�ⷤ�_��7s�LW�>W��n��g)]�U���j�r�����:�4��A	��X����,�����z!js9t�I��Լupzu_��u��i:��1*ME<7��6�t�5~��]uWO�u�
��Ȣ؋4'���6Z�1>�(�bz��q|�	|�kuhC�E�N��3���f�ǓS��).�O��~��(^�J�\����J}\��T.A�����K�z�q=輹�j8�46^{����k�j|i_���Iz"Z0��T�Bº@t���xIs%�1�v�z (��e%�q�3����C���\,���f�(���B�,�<��~v�ң���b�;x.M_w]c{ݓ|a�jiXEע�����h^Р�|R�X����
XV����)�Zj� �렖��ѻ�~{2��m/X�A��N#��E�=�@���!\R�C�u�v ��+����*�`d��E�C�R9~V��=��]t���s�I�V.4vy�/�A�Fapə��P�fzrC�� ^�n;�=��i%��o��#>�С�ԍ����b�nϒ�ׂZo"���S�H}C��1�~����M��Jv�SS��N7����r�ٜ�u5 ߴ�Q0p�b[�РzǾ\���%Q�=�ҏ7��yYq ��?:*v
�w���#�cpkP���gy"��6���T(n�J;~Uv��_���C3������V��JF���o�����4
2�����H���)1i�N�藲���!�vw4\�x;{!�V�{�])�W���6"�s��9�������V'i�b�;s���l����z� y���Z����Xꆝd%>�EA��F�"iѫB�y�j\?���p
��vy��N�1Ћ�jZ�����7-�o ��
�4T5�QY55�w"���̎�g�������D2VW:��@�%%~i��-�)�ǅ/$>14�O�{�;�4����� ��w�&��9�{J�
�&#v#���ل��`�	�q9`����.A$�j)��H[E==�.JץW��&�Ȣ��!�s���)[��%K�B�ǦJ�?|w`�����/v�-[�vM��l�����3��X������'��Q
Grx30��3������T݀R0�I�
�	�P���c;�y�"��͈��$v�2�U�-G0�3U��.^3��~Z��W?

V�p�eG���ο�g��OC ���p�LC�F� �e�,'#/�21]q�Q�-v�L�դ�6����v �7֘�'e_�0�`� c�Av@[~Z��4 �5�i�����!RP:09zR����9�H!��Puj6��'�*�
Mf�Q:5����~9w/�&�}p
����SڑZ3�Ƨ���
Bq��s��:�E�lg�ӱnK�vq�Ђ��ji��x
X`N��e�B���!�\���2��]Zx`���
�/k'�ԍ�C�$6�Ho�*��Yy�Ԑ�u��bf�>�Jv]�W-Y=̧�X+�����50 8'�RB&5,�v[����^�S)�_�<2&�v�A�@���$�j�w���N<�	�j�Zg,  rY$'"[̾'���8���g=�����2��0�W� T�:��yF!��L���W�TA,er�{������> �N#z�@�����Hh_�U�|(� �(�ӝ�$@�3X���Jv&^[���ӽ�jx��:�R����vPIC�JI��Lv�t��j�&�����)K�s������1����5���V�����3?ޞ�=�p��u�4h���ףy�n���m��u��IX�7ONp�������x��a��D6��|�:G'�#�DNuV,��P��Z�
|3����\2q�
[ί���EJ��,C�B��i\m3E ,7��0Ѫ���,�G�Z�%V�@$o�T�uwq�썇*:�`6�X�x������j5�hxP�x�=(�nU�g�)?OU�6	_{�!Au)Ɂz�����8V�qE�Э�M����*c��?�q0y��韥��,���_��gT��#�2�3.ԓ@q}_������i�Jo�`��I��.�T>Ǜi���ژ� |�B��3k%?��˓�{��q���ki���F!dH�w�pl�=z$9=�p�+��u[Ԁ;0ˇAN��h��3a�e@LƏ%��ڀ�_�^t��\=)l�T����6�������IF�6V�x��''���%o
�r 1"�:W�;����bf�Uc'��I���#�=�e��5al��P��� �_E,�͹G�4x&5�`�����իUp5��\.�~�Bs�}�;��Ht��-�sO/����,
�gECօ��	
�^p���X<�&M�읠n�����oy���@�^7�,��>ޝn[�0�]��qNc^��z�O�fR�S�\��YSTdƁ��p�-DYv.��Cd��S~B��/��E�k*�ل?�d!�m��ylr�!W��HP�GÖ�::R�3���bW�H��D>K&�<_ǃj�np^t�� -h[m��^$���2�>���>�Wh���ݱMVQ��ד�ڀ�&�LQ���0ԸY/4s�-
������8	b��l�T�f%����AGE=��lI��d;fqX6��]� �`�<�VTe�n�#ANY�3#��dr���7o:�D�"��c�=T�9��5{J�ҋ��gL{����Bk��n�-k���Z��2P����q�tc�f`N������Ε��q��SW�$�!�N�y6�_R<�����!��aB�'w��(�kH��&�m�=�S~o�z��Q���d�[-%bx(S���\�տ�bQ�qa�`S���ut^�q,shA^���,��o�D��S���he��ΰ5�� ����tu��E����tC��� Ȱ�0�ā�����WG��p���I����$�n�'����M���c)���G�3��{�a��J�$�u��'���T�M�@�����@��S8��.��֋��hP�¨�l�����M���G�Ҙh�wfnܩc1X���z��pٺQF���E�ԉ��vP6��(�ĝ�ܒƵ_3J�H7y;�LP�;b�B4ݽ���F�z��E�
��D�n��:\������Q�O���Pa�̟n�G�zVmp��tBXO��!�䣘_�+��&�ي&�5N��> ��gc����"Q �D����
���ׇ�&�qw)�b�f��K��h��s{���/�/��5�;�\��$oUKY��j��g���Q���}XF��V�G}~�%��iW����
5W6�Ŷ=Oc餓��m��Ig���")5��Mda��@�����bB\P��j�`�%c���*}�%��L�L�����t:\GJu�R�2�ݯ�m�&̇~���RJИ�_����g��F�6V��S�y������C�!��rQs8��=~N�6�9Q�E�d��w��utz��`P�&.�7�yH�����V��d�V%VW�u 
^����ɀ�Z� ����n��KN��&��Q11�o@M��~�F"�F
�D���EHq�H6ɖ�����PGa�-�����&'�+E��P�����ǩ$h��%�\��ڲ\��Зe��U�mh�I ��S�v[���;��zQ+�u��Kt�3�QdL����:�@��E:�r�J�^�Eig7\IX�[O�޿������,���� c�&�׏�jMfפ·�*���^��
���؆q�>�N5�u�m��+���>�ǭ���4q^�V��R�h�r5�^7<��M,MYe[*o��x +_%�҉��:F���e_3��ަ9�rzv��ӂ�j�S�������� Ҽw{�!ɣmyy�V�!���B�#����]~D�6��,��R�Mhg5&�L(�nÎ�Ib�KGYp��7O!EsΨZ�|�J�*S�f�>^5ׁ���u	EF��c��Ǎ^��f�������Pꠒ�$�f��u�*|z�e4i�^��X>-f�=#�e���l��w���-a�l�P����j����)G��&�����>�Ш� ��f^qt�X�"`,:���/S���ۂ���X�ɰ��L��$�v�e��|��]3��f�'��[I��I�#�9=S/2E�L������c�4dS�-.3Q�e����I�Ei��a,��'J�_��u�Ӑ5��)��d��Vu�a�@
��3,|�=��Q7S�6����x������V�e�F''�](���2����*�_rLlt�A�P�y�$��u>����T�}��'��9�0���+�cD�_o)~g�J�=�;�_�N�\5e|�L3�S�}���B�ޮV�D^�	�G�����#�H�doփ�x��`>?N�)o'V�h��S|�eY@��I7�|0��ğ/���Jy��v"�z�R��U��y��e�9�3z4JV�24�Q�I�aA֏C�W��Bk."�����"�maK��A�p9�ou�b3h���hJ�g�A١� 1>4� �C#r�jG�wN@�|�1�!�&�9M\rB�C>��[g�1Z7=�E}J��ch���/lZoί_�iݣ;ἂ�jBK?��y�#�$Q(��Me�ؖ� q�*@j��OA=3x�+����i g�	"ؓu��~n�%����2��zx1a���+/�n0Cf>n;g���Y@r��"Ԍ>#��J@G�]s��i7Kڽ��I�z��	a�>O����3��?<�Y��$��z���
�&!�t�S)�UM��p,�لD�-ǈ�ԕ�[�]RB�������.�%$���6bKB�V�D�2�.eW:�����a���9<+!���i�m��1b�Y�J�Ȋ'>82�C���R��%����DFp��������@��Yax7��3��	{6{�T%�ĉ�T]rg&N@��h�D��L��U�cT�XZ��k|/����p}bXѯ\u'����ڸ��4lE�Z�c���}����V�\0�U@JUʴ����M`��J��"+�Ԓ�%?g�x�~�YEaTEf��p�WD��%^�(�j��݊��o����	�!�i]�<<�zg��Mo&3��������5?2�CbhD,.ضɷ��@Oiz�E�U����q���0����jK]�k)�'Ќ�S�ף�̩k���4\tD��c�FIIss͍�^z��a�-.��d����=ғ��"�y�w���"`f�� i������¨eyz��L�Uxi@]�n�]b<�?��X�vX�,:���s8��l�І�H�E$-t&XU�)�P|C���UC<3��;�Hܨ���MywĖO�x�|i��e{!Ϙ��mŦ�7[f ڍ}�N A��<CuK�b���A�z"�A�J�1Y��+�oLw��K����o��o")�b&K�lW1G�sl�qw !Q����Tv�Q�4
k82��%<{���#&N���>���W�"��zc��w(����r��t^�c��.I���
�(u.;孋��_�>|���dh�f�O�);�n�r�ע7]��<�����F��|sEl&30�㘙�$�17S�����-���s�P|u����=�<W���6BS׾��'��M]̀�WE�3���]�=vv]#?R�]��H�A�AY�K���ů}+W�C���\l������[����?8�=�h�`�&ei�ׂ�4����T���`J� [-�<�NQ%��p1��F(ߦ��8'Sɪ=�CKLx~��Jv8�r�梲���+�b�UG�b�=�TvY� ��"��_RB�\˶��\�#ż�6	�ݖ]��X�b�@����y���Fҭ�輠�C��~ȞC<Z��(��������柁�z�� �G`��3���[5 [3���W��O�}�����0ŠvZ]z!z�{햏�W��q�a���fC*�lV^��ϥo?��1:���ϟ(�F��� �B����/B���,��Y|��g�x�5,_b?�P0�fa���ّ�d�϶��<cV�zt7o��Ȼ��"�����9�hb��-/��&�k�!i�������� �rX�kH6L�~6��۴�o�)���`�_�BT�d�E�'�Vv�/G����r3g���&:�I�о����)'��j�`�K�`(�2=N#yC�U�A��Vm���D�m�~E��>&�?�����٠?���\�*T����l>gٙ����1��,��|1��A�׻�/wX��P�>��A�xd�P��#����c�_J�#�T쟛�t1m�����V�&��B�H�֞�ޠ3��Vb���8�tP��<��I�6|Ⱦ�Vde���9�	Cq�e�ƦT�y�o�L�̝��,�f�;���z_g��K>��-Q�JQED�+%��$�&c�r7`W;X�y�P�j��/y(��m7%�k��Q$�L0�a��v�7�:�آb��P�zl�Y�|a�_�'t2ʮi��~�1��qL�͋\��������=e�L, Ɣ����]���l�q���}p�������J�\�\)���*k9υT����Ky/��S�~=w!�=;;"�' ������h����J3�֭���XM�u��Y�4��ȹ:��V���H��f��B�r���AUN���[�И�?�l���/v����Z�m���RV���x�as�K#Z�3�Z�����j7/���
��V�i (�N��\�`��/���/��*m	�p
���� mJ�̀v˹��}+��#��g�8�hd���qoңVGn�8I,͵�UDE��H��)������ҷ�V*�鴏����Oi)	��q�Ѝ��L׊�:�A�@�����P���L	SEK�i�9�☚�|��o��Îr+���D!�a���c�V�>7=���9������D�SJH�q��`֮Fk����QB;=�ը0.���ak�֥������π��B�����⥆�ێ�}�h�Q,�Pd�'��Q�N%�h���A�����)؅ܳd�\[�fwۭ"���r3���º.�J���3�m�����A0�����	�xy�E��s]�bت�w�8��8��4,�䑡��uց��Y��C/�h���Pj��d8�t�*���Oήk�,����-m羇��7��%�˃^�YA\���?���e��K�lၤ4���X�pך���Q�K�+	��M����>�yR�!��X�"BI7��p�6� ]�1��8�\��}�z�Cgθ��n�q��L�T�Ċ,�=�^�ֵ71��H�^,�m�Q�۳d��-�Ab�{���� �[�X��%�^��#e�_��
��zd"�nO"Y��BC㻍{�x�� �+,0�Ph�vU��h�?��e���$�	,QN&~	�q�J>"����Jڱ$R���Z�����V������u�¥P��ڄ.bw	��}D0W�i(bM�� 6	��J|&�[���W~�;����M:��`9������8�ʕ����!��oi��q���\���"�"?�bi^孎k��!\�Q�e}y�����^Ի���>�|�����"�ak�7�����5l%�U�)��0Ȼĩ�l�؞Y�O��)#)ĺ/�7������ٶ��+���!�Eo�7B4PaLW�(;��\���Wm^7�&�Lu)L�b`Mss��{�A�A�Ixb���v�mxaO��}ڸn,|Z&]N�;�)=�/�v5�IR� ɽ܅m�ѝإ(��"�[�P��V�p����fXq��]��yVd8�RR�{'����!!��Xz�@�aX|������5H��_�Q&��'I��x���â�!��X1=1=�r�X6�k'��=e>*x�8���6��F g�Ϡ4K�[%G�9�ΐvb�-� K*�j�!)�t��^e��Y���Li���t�R�C��,nX�`g�>?���</h�;x�l�E6�bUwe���6��h�����,׼V��A6��%�q�Ԝ�P�q��c#��W.�LIɥC�@G�����%�T�9���������|%���O������*l�l����������(���̭Q��J�e�uy7�w��n���>6�FtR��+^�`>�C�v�.�/��eQHT�w��i�0����H��R[%�m�7�Ŗ�I�5ya�a|�a�p��iI8t�<ݣ�_O:0*��`7��>T��[[vnAF,*�7-k0��ON��EN�dL0�ݨ��H/��A��������'&��P��A(��o~R!��y�:�Swfe���Gl��q��@���B[�FBd��ʱ����z� ���_d���t;c�F	�sM��{�ZQ��(M���䪻�РWP�ɽk��R��U����`\���;`,~�ֺKB�5���QY�F�ꗆ������ä^I$V����x6��`�5C[��}��� (.�Z)���X�zQ�~�!>����mB��.�>�s�g�wŀ#���P�ȹ�������1Iffu~���(��^%B	�O���=�%8[���1p�=�i��tC�N-��d���U��liԔ��������4�~l� ��"ne�.9�fd��h�����D���Z����ߩ��,#^4dw���-o��툲�m���A�v��8����<>s�t��k�M�Cݯ'ů��BN���'��;˰a�H��RC�G³����m�oR�)�����9������Ն�ط}�쵕Eqa�UT/�osu�ff@R�X-� P9��0�E���&�s��b/E!�JOru�tO�=�̈�ǭ���^Z���DN?H&���fU��{Z����{����)pj@��]�:��*`�HWt~e�(+���5놅��je�<�����Ys}�
9��7��y�42� e]<h�{�?T�)wAP� �}�˙�lb����8*�D��E�zۛ� L,6�}y�g��x���h������#��ຆ��N���x�;nQ*��@d�xV��F"fq�#!o�Wi�g�2ie'f1�>OI�Xx���z�F�DX��%���7���&�;��s ?{s�4�k���&����s��z�D�>�n'�RJ`҂/�Ԣ�F�չ�TM`K7�du�T� vPML4k;���0���og<l~�}4�)($�0_Cށ���?A���%;L�4@M�I�%��L+�ErQ�9j�}6N����u��C�i��V�����,�-yْ`@�2��_wV����C2ڂ�Ѯ�T^O�w�)~�;��X�&K}W��z���|�I�j8�fb�9�����1�x���+���J������X�)� ��=C:v�*
�{���&��D6�hQl|�GI�oEr�w�d .y*\S�9z����D��-Z_x�'�biݶ5:��Q\���]x�;��[Qٴo�u���TT�u܆�Qd�̑Y-���9�޼dz�F2j7 �I�m`��Tk���[r��k@�v�jb�vбF��?d����ל٥\�m"�Ob�Z����z�3��'V��^�y�p�4���&�%+⽌�Xt�I���#8J�$%�nh�fl�%� �5��=k����衽Y�ԀY���<�_;Ѽ� ���$ٳ�{`B5y���� 3�#J�ӂ�����y ����We*m���?��ޮ1�݃{-e:��|��x�Xp���T|it�k�M
87�NF��QxB�&�e4Q�L�4�0�y]��6���.�śr����9���x���p6���We3F��#Q�} �i�kg��VGpbA.B:���-�hd*z\�\/�7�L)Ԉ~��c��)�ʉ��Xha����x*t�d���J)�e1�e�S���?�(in-��;�m��D����[�L�K���d�(�l�}h��� �4�	�ڥP��P��1v��ⱚ�M��n�� ��ˁ$��,�j���km���(L�Ó��$��M�)�@�˩�1���QY�`,��)��?��Q�9�*�V����s��V�;�������
�$L4w�ga��;�ºY�_q>3m%ڡ�n�C�sf�(����L"�P���JD+��f�S��B���\0�D�9�HAJΫ9o�L���v�dd.P'�4��ٍ�S�$����`ě^��:D<` h ;��Ə]p���s��)��j"<?���Ͼ���8Τ28RO�ܦKL��w�X"l�1S>v�[�/��q�q0JFk��M���[S�I��5*5߽\��UPH_�WI̼[����0�k�1�>m\��	��o�������"���@��� 9 z�L;��L�V�ͻ��n�e|uF˝J��r�#���"�:q>�b�WYP����j&��/]�.��6�?�M����n�"���t����qR/�)��l�N����f��+����%�*X�����_Oފ¸Q�J�JC����DO�f3M�Wc�<{a'r�K�fvW(=�e�&�\�*Q�����M�l�����h`��2<c���c,�j�5C$ ep�$8��=R��sbɉ�|�.�Kֶ�U�$���A�
��Bk4ܙ<���W[�
ٷ�=���G~3n�8 w.C%><�.|O0��4��6�ߗ/��Fw��u^���G��O鶐�_9�f,�Lu�m�_%%cN���xR��t�u�������{�DCܱ2y�#*���E�!;��jo���q�zZ��S�����~իF��^\�bah��:JFDW;�?�"��9��acK��x�%��{?��<>�m>�GC�s>��'�g&� �jr,��l����eGU3�}%�i��.j�k�Fa>���r����wU�]�Ǐ�EC7n�s�j�i��M�,t{�[ס��=�� F3��L�� )�m���ɋ�J�o6��555�<WA���#�1��͐��L�r�a�+�N!iFE?u�#u�Al�)D�\��7R`��{���N	�i���q��.�X��(������$�|RƩ��@���/>N�Qf��0#���q���v���(8�	-�@B\�B���0Ρ��s����P����?���	�zU�!+��Z0 �سt=�H/���Fc�ŗ
^�7��U�S�p]8�z6=�<A?���.����3;0ɱт��Y��O1 Ӈ� d?�T1߸���C7��O{�ok9�7�qe�����:䵒��P��[�Ҵ���O4��8�Zz��1�dғsH��l���
� ��p<}� �ڎ���xm�����TL�M#p����=e��4�5��v�ۧ��,�o��m��u-ƞ��YȺH8P�1�݋|k���G��ŧx�	��"Ybu��քHޗ�۰�P��>�lI�؟�9,*^TP8��+�_j����@��~lUP����8���6��N���ͷ���S�D���3Rvb���C�Pp�=W���\��NՇ-�J���WӁZՓ�]A���۷�im�!F��Vq�wd��Τ��"!Y���LV��ʮ�v���a���?.���K�b����hoӜ8�+�t�+=O)wMd��
90�ۜj�� ,��x�aJR��Qf&_EѤd)Ujs���B�
(���li��Il2|�[�b�Ƨb25Σ@W�1zF��}��1ln	��"��HZE��5��C�t)(��<i���1�F!�{�e��t�O)&h��5"b�!h,���.�эE�Af���'�^6�֖�(��>��� �+J 2���l^.#K�U"�G�pP*W�\�W6>���j�l8�-�p�*�f�!�Tq���=/+T�+�bM�	�J޽�i'*�(s(�:�?�S+x�����q���m���7�*_T,�C��àL=> ��_�|}��>��m ��@��Ԍ���b�����&^�I>p��w�>+�T��a��[j��0��Gy�\d�0��SE����۽w�6٦'>�9�h!0�$H��ÊX��F9O[I�S���ij�x~z���7�Xe�;�3
��mX���W��RVĒ̈́/)��&<v2���*Hs��W�����2}^H�>���P���т�݉x�ER>�}|�%�N��/�\̼�)���:��8��V�cle���&��� �i�w��0����[;�d-iTd�D]�g�|s�B�xA�~n�r�Cu�ia�����euuVM�].`B	i�jm0?i��m+dXO�+>J�S�s*t��t��򣎑�Q�1X���J	��,��Sw��n�b������H�}�8#X����uUw�3�r�/��kC�N�.H�I�s�����4"�BN�����3��U�ޗQ/.1�Y��m��"�M���ܠ,��eI���o ����NL�`�`.�C�I	TɊ?��~�-C1}�gzP)���	��]3=yHɚ��.8�g#�܅}J���a��(,Q�;���0�����0��g0G�.(�{i
0����O�wP$�3-�
���LcA� �RnhV ��q�<���I�2Y0��5%�$J� ,�����=�
!�?~A��ec܀�Q����,�r�sq��w�[����JxV�f?�@p�?ە��o���pQ���ُ�P��I_8��V��x)~�)Hh�dBin�vPٴ�@/��WK%S֪��4�*70�D��_���4����lt>����\��+����wU^�����&�nP(���<j�X`��x�v���{}J�N��"��c�0�np}D�Y������>�{����B�h�Ji1�s���q��(5ٚ,́�[2�d�yJ)��,���+�hي� U'��S�01�-�ڮ�
��3XE8�&�'L����;#Y���]�|<�qn"�`3:�|ͯL�%�.@͉`V��f�Ag��;p�s���=�#\D)��N?�JLM�lU��]-�'�m��v[���N��c4 �<F�A��[=�`�+�|ه�i�n{���uxN����ی�@��à�?ؖR!�����2�?/҆P���2QS
Z�N�G~F�/2����oGO�.�n�v!���D�1�":?�GwY�N¡��� �����B�4����2Q�;D���$̵|�ߨ�oX�<=���4��uF*Xf���#�1{�3t��GV4��7�C��=���f���y�ѹÐ"� �M�/�A����\����,�:f��V�8�>���*�r*q���4�I/����=�Ð>��R�a3�$��k�('�@���V��(�m�`��~W�~�=�%�.�崢h�����`�-�1IJ�JH\i�׀-��,G��y���w@T��r��g7�jU�U�,\0���OA��A=[�@*��{~Y�>��V��+z�Ø�Z 14���ܢ Kh����@!c�Qo _���9�3�޲ c�Q�4�~\��Ǣ�2�B}�����}No��{UFuk
����*m		�� J�Ơǧ� �$|���������[,L�,�#�j�Fv�ԞQ�!zw��
1�@�:M�#�^�s�`,�����3tM�F���z�;h�3~pk՝����K�69�~=�L�`ςp�d�T��٠��8\���b����Д�LQxD5{�_[��^T�}�|@Ii9f���N�?G��n�e��$�^5D�G}�Y1����`K��A阻�����޲\9"I��Ayz��v��`��_����mQ��\ ̂uH�>F�m���#�'�?���xF�D���J.��>T�Ƞ(�-�C��t���'Cp��-8��V�}�����'mjF4���4O����2X"�Ee4�.j��	���z�e����q��xd��ͱ:�����8PWVrχ�޻I�[�~��E��4�$���r���7�o=�a+�=�*�s�%,�ͮ�]�{ ziBJn�AR�)ax�o���F��c-�rEЫz2*�nF�K ��	�Ą��p:Ș3��D<ڟ����
��Z�������#�<UV�	�5�P�YO��u^E��vC�Mі�2L��#x���"�|g�^0�Xk6*���sKؚ?�@��i^IZL5�ܐځFs��9���{4kd�o�2>��nQs1�l�[ ���Զ|U6i��p�1�!q�������áb�.�O�:~D���n�:[�z�MK*�x*�Uɡ�`�;WG�I��݋י�ű���o����av�S4P+(��!��
�ƺx���<���[�fX]E�l��Y�YS��;�J�����(,g��G�Si��|J���������,�,4���Au��sAM4�h������*�0��E�@@;�x�H5���*`"�L>���ڥ�ܷmi��;���$;����uκ�L,$x�n�p��N��sǐ�qfǁ��Y��Z��0k�!�~��I���-�m�ޓ�\�Be7a����^�M���/SSK1ֲ(s�������v�P��|�H�e2!M��i�Ι��?��5pg~Ǳ�Q��{r�u{���?�)>_���h.�ę�r�m�r1:�����kfW����Ћ�c��W�kTFeB��z���:����$����qSƦ&����`�s��n~��M�mZ؊�:2�u�ʯVR�������������ޤ���Lg���c/�����2_��x�+$�(+�c͍���|���V�y��S�2@���K�}���^���BނT�@��y�kDS�>�'��_~K���A8	V��L�^���3K�(�t�Vǎy]��<v<��`��2�s��Î"Gk��Ї�h�xo=��1���x?�=~M�Y��5E�A��K(__�p|'�q*�|���������/+��+�A뀕<�4��ּϔ��eXX W��ߺ�ԧ7�8J�G�Rz���s�,e_�LY@�G/B��!���MV�!�.��٪�[�5e�q]Y�|���_�hD��ڂV�}4�����q[G�=6Ğ��>��<�B�c��*Yg��*�I뷎��B1���)h�fiL���D��ǜ�H�O��~�8}9U�Z��y癒�o�S9ޑb� ����Y=�N�M5�b�;:HH���[���p��r �V��ԡm�k�qVm����G"��3�ֽ(��ׯ@i R2I|�����_��o�|
����z7٪���7ԑR!76�̹�F���`��Mj�J��]/��k�!��Gc����om"E��&����u~�0A>�4ZX�� =�� r��w��=,�0�}�˘�H)i{���C!�
^���5��}�e]�
�~V��t���j{��Z����w�L�0p]Dלc���gS�l�S�J����T���*�(t��"���9#'U�+fJ$��c��uP��X�F��_��\��� jM�M�4��giC"�5�ժ�}����\�?Ѯ����no�`@:�Y���T��i�Ch�-��4�>|��2�6XB{bр�F��vj�����[N�L2tT�h�U�i����1�Z���	H��w;k�7]�)+r�Zi����ԛeh�hV*�^V��ᅍ}������9�VS)�rOLNљWx��c=���-5�U���%���֏��$kqC�띍��;S"�$OW���x����FM�J�l�Jh���t�1
aw���q��7���-���49B�G����5��O�5H���tHF�%�v�7mb��F�dh���Q\�3���X>�A�Mt��w"6}��H��f��8'�ɡԼ,m���G@�9��<
C�H�z�y^�VcҮ��G7����nS���튮D;cT�4�� �u�=��u��SX�%S���B��~�n��t�з8���(-�*��~
���p���0�4Y4����~���kBwj���@��n�����ϛ��.����2RF�QG�)i7'�<k��+�>�h�O��:�R�,K�a49�G��X��̝m�q@*,��ѝ0$�H���:��:�q��j�>���[��e|{�>)�镁?iA�N���[�C#�~��y�Pӯ~�rWZ ��Q�O0|���_FLin��Έv.�wp�e� ���N�jM�13���>Z�p^F��[Q�K�▖;���	�h9���W���i�mB>���H�&"-�WT�oZ[�4~v����V�.�Wi�j���>,�>&Q($A{}�@bZI��8v٢D����;s�]P����!G�QX�99��>Qh*N(��p�<͊�0����hy��9�[}}��v�ˢx�� ��H��;b<��[������������$L9uݔ�ה$y~V���C�?��qtK'Bm��aƳ�@v�2'o#���x��C�S���%�~��z[�5�������D�� .T� 8��E��Q����g����CҔ���6Ɛ���߯U���H9YpI]�Y���U��s{7���?�:o�ZM�6�z.�C	�@�g<��PP:�T�f��B����-vC�����;�6El�I���ǋ�΀�ʈ<��6���ˤ�Wp�eW\� ~=��+���*���YuB�D.b:L$y	�ڻ{�.ӗ8��R�،#�O}/Qx�Hx�Vq-*bt�mO�I���&�e��H� �Gɻ�����2��l��f{4[��ߤj]�F�B7EG��m̜l��\��qЈ�w=�c���D�:ǴX3ů��M�C�<��*h���ꨊ*'m�$���9�ݔ���nU�6��[t��~�l� ����;<��Ѥ��vj���v��ۘ�qၳ+Ò�>QϦ.�xb����\s!��N)��{ޥ���5J� ��	�1�A�^ ��iG����ap�c�KК�qN�r�>{)�����Ψ�\�+�(�V�Z�.o�Z���ZAM-c�63^�`��|rN�F�ehg?3���_\��,{�g�Z��qd 
#��7}~-�X�cL��@�omp��̌��P���Ŀ0�ΰ�X��@;��p�A�r�B�}�h�"�y�Q�oEf=&���T@�Yf:����{U/��躢7�y(`���q9���2����� ߤ*�R���te��W�-����]�o��S��4w���%l@��Ǯ��w�*�i����F8����c��7�����J���������O���q����l�5�0'n����[��#���� �s�����5C���!D{������j��=9�� | DS'��
e�:��������qY�B���K��3�=R��nip����o�b���FV��k<���
����U.8&oQ�'&�6�K��m!\f<$w��˔W�Z}N�m���wz7v�?.[�����U��Ie�ɵ0e�|�p�2f<�y	Nsk*�7�jg�n�꿓��#S�!�>8�j���z�}�
�4i�|<e�Z�����a�`ݞ���}�k�T��Łm��gP��GKf&z���_�0�2��8.�k &��C��f���PP�����m	�}����k����E��Μ��M-H�^n�V8�51�F�`C�v�y{m�J{`�,jM�*�mҺ4ND	;�G��b�5\T�.-���<�,���R�ݴ]��g���*,A��8���>)s���͊_\�;�H�>�9;j�mP0�6XB1��1�c�E�~A�J�!��20�i	���\�ϵ��7��l���Ѭ�iY�of{)����ĩt���B:B�H�����,fJ����C=li�=I� 5d�|�i&*.$�p�N����c�R��Y
�`�y��8�B���Y��2�Jq,��ֆK�R�ߠF\|q�����>j�T�>}g*�)�'�<�v��ћ=�H�W;%�x,X��n�]�ע⹁�!(h�mH���z���g'��̕�S6j��n�MU�;<P=;� ���}޿v�X�b���^b-p|%�j�0f��U�|�A���ͣL��h��J�8	�E2	N���*���Ij�,*&r�C�c�E2�:_ ���e@OMwג:v���:;̻yh�Oݳs+��U�%�!k�4���$VZH|/� n�^�I�u6��u$x�6��n������܌��Qf�B�<C�E�k!ׂ������w�0��6m{�q��$��n����˳��o
����]���I��*�ĥ(�l!~���^�TM�3ʖ�w��?������5 ��IN���S�
�O��s�/��G����+Cb��{�I5���j��@a��<o�y�p�G%<�͕-��5�
��FG��C���ޣz舗�|.֞�J��x�Gn,�вך����E{r�Lf���@Y�[�����+�������D�S���lU���l���=IdO�>E�9\ՔK���ׯ���'��{���H�Q���;-�Jz�V$�zK����1�f���Ǿ|��C3��N��QE�� d�	��s<��j�c�~r �:$&�N�-/�pR���l��:��M.*}Mb.��wF_%<�φl]2�~!燀�/A0)��r?�]�
�k(8�|�a�b��'*U8���"�?���ck�vd�cOF�bf���>[�[��#�Y+,�Ë"f�q\mw"jT��d��C�C!S�L X�b��d�^w�	kjg%�N���SZ��LM_c�9�X��3��4�DHn�%��0�?L<��y�둌�f�JV��a��v��tE��@��{Z�������L�	�,ԆEhV) �<��Bj��=��.Ă�R��>Km�$+(���uQ0j�N1C9橄{ƒ��*���d��D�w�)�iv3c���w��/��S'���?ԋWN�y�$1˹k��j��t2�w#X$�γ�1�~�x�] �~��f�s@�;�o���^\ni7u�e���\^�'�,���B�^�s���oRO�$O���pA(�Y�/?s�6�
����\�'L죏��d1�)Q�gȈ���āĖ�l�M��aOz+=�J&�f���j�J��o\�o��>*�S���0�� /.L�k��+�)�ǲo<���9���V#=q6�a@.9�豲�&�е�-V3YУU�C�^˞q�k1ϥ��МO��;˂�H�����Q+n�X�3x��w6�����J�ox��ͫ�H�$��)[��xR�,�K���8�׈Wt2�ʼr��}������}�̘��#s�0F*s��n��#�l��l}0�1��K	{��B�X#�N	R�x���'lz��ܧ�,0Ų�=(�8�YM�����K�h:�c�$��5�<S7H]q�J}�0��5���#��Y�9�1t�s�~W�*��"a0��׸���"+:�n,GCZ3���3��#�����Ye����ogWV?t�Gw�pB�E�)�3�-�F��p[�b0��X��l����Kt	�>8�1���V�@nG�x{�A��w�O]H���D��B���:�J&gT,��#���1^�Ώ���FCW�W���Ȝ��k�Nt��m�n�E���oP�'��5)��Z��<��bU�Q���S$�N��(_:�͕�����Ŷm�4��+��k��iX���*>����}u,�:-����7ZkM_��N���!��>5BT,�j��!Gl�Hf�c~ s��6W�@ M��5�҂���1�&.�{,wPI�z�2���P�0���*��l��n����E��^�����i�T�0,�W3v��J6et�����r�?�xצ} +x�ٹB�i�!�-�~�#���_flj+��B�8hI{Fַ����E�ฝ�A�㜓w�%Il`��!*�|x��3���Ԑ�R�P�r�3AA����RYxeˮp�~8vp�zGy!?���m�4�����ž�s?^��E:a�����v\�hC��[�7[V��p�(�]��P
]ݚ���c�mD�}6FLM�Bj|�}��1����xHeU�sm�͜s�8`��1Կ��D����gM�Z%�%��~����c���$ũ0�����
�ٿ0�5y$�~Y�L�쏀��cu�/�*�4��g�\J���Xa���/U;����qF�bL�cn�����g49޷�VwtPp|������E��e
�.�=��^����k�e�(\h����NR�R����Ju����,��Re�kG(Ez��ݎ=� ���S���z�� ��W�!�>��ݧxX#Km�u�$��ب��f�E�8�P����,�^@��s��a�C�'�ͨh )�L�{�g�R�w8-k��U4 �	̉i���l�k���.���u|������V�y��8�0:����Xv�+��K& I��jka��F~�Jx��j^���y�����6��.j���B���"g�y�c'/m0,8lOk���$7~�<�h|���W��i؝o8�v[�jlf��
ƀmL�|�L�?qZ�K�	`��f�N��ܰ��'PWƱ�,�{o�|��lƈ�m��W��]c��b��c����X�{���V)Xڭ}R�ʙ&�E�LEcB8��*�%����C�$t�,Z��S���{���PI�K��J�����.�s���茻I�
�v$��p&đ��^�e�,_]�hSȉ��~���b��|�oڨjmж���͡|�߮��W�0n����?eZ���=Y�~����]7_2�k5�]�Z�����=+c��{���I���*�.��qA�{7cR����;\�6�2\!,��o����8W�	uL���S���]���h!��y�TJ9S��Ձ��`�z�pE��$�p�'*>n�sN��+�:�@o�EeX�K�h�g�،��	��>M�պ��<ϯnЇ������X�f�P^�ڶ���-�o�f�e��?(u�`u�k\�K>wέF.�\����s5M��T1��'�6~�Y2D���3 ���E�;<:�4T�`���/��� @���`�n�Ȉ�:�9��1�hL�z-��i���X�>>$A�̊yA�A���\!:|w1ǯ��6�F�&�{��ҝ�zo�c�:c����EWWsآ�k�`�V�K�߳�q�5Iޤ1s0\f�W��k����u�s�p�Q�Si#D7v����26M5q��?��i�� ���:u���.oj�"d�<|�yQP��%\�?͢����/����J��J=��,-��C�$���@�]�u����d����ֿ�K%�2�~M�@>�ݽX��#��"F3uzrPF(�j�-Ɛ��d��a���/��F�'8��Ĕ��z���M��d�v9��]�BȺ�C��q��H\��W�5�,&��e�y���=\��2b=��b�l#���}�/]��Y��nG6%!.��B��ha��r�|y_iv�����
������_~�F�]Q��}J��w]¤��W3L���&�>�|o�S/�6�D��N��!r��~~�+P��1Yae �mD����0���J�U �(�I'�U�_]�N"�ɞ��ٹ�ND��	5�^�4N��p�:����&������WSű�� 0��خJx1{a�K,��]f��(�3��������1�����
y���k߮!w�a�6�]{�ݪ+��<��uJۃ���@�Vcm%H�y���4i�]���WR�YY��RϪ���7,���i�7Tk,�["��*?���_����R�T���̔y������H���/�q�u}�	�g��601� F7j��v��U4�y�\�� T���u�Ι���T���~��{Z]^�bξAh�J�|����|�%o-}�/��Tq�w=���M��f������K��(�4NNXۮ��Vǳ�*���˯,�+�L���]���N���^��t��v�%67�
 ���i�d�P����� �8�P�m� �����T�k���,��[�w����5��w�?HZY�2I=+�;�O�`y���2ؐH�tƌ�"�.v��NKA!����t��*�Ԣղ���B�-�����p�։�<L,`�E�98�%�A�xs�"y�@��t�g��vXܒ�JZ?��6�������CYbQ������M�$b���(����l4IH��:��)��$� �����t���k8,�}��炳�+� Z�_N5��]���W�V�u�]�h:�W�!k�����lk/�X�C�z���%{�ݻBt�U�D�ʶC͈���B6��`���Y��tNKD�90\��0�rx<�ϹI�r�58�܆۸��zpWf�����i߆�|�e�;���� %.��w��jok�ܰuwD�R�|�S�����\��%�d9[t�96�^�?�6l�+��Kķ�?�ϯR��7^��q������������������}ު4�o��=�3�3�bK�}��9��P�� +N 5�4J\�J� `�PF�/}P�a��~ZdS��r��/�-�!���f�u���,kF+���V��û��P�����oU�
�2�؍+�dV����$UX8s:����zღ_!̝���Iɂ��h<[����0ѯ���9�c%�88ԟ����B�R�U5�M�wOOPk�k�Ɖ`~T5��.&���d����üqs�#Y�c=a��p��-��,�=w�F����֚���(�A�_9�ޜ��,H>�d��5F�EU�$N.*�A�O���/��r������|z6��Mf��g��8��Ţ�;u���QS}Ik�+����1MU!ѝ�}��`�Z6�U�r��yB�$���9}(�Dq��;��/�¿-
?�M]��j��X��mo�~��Pe�uX��=�"kW�Xub��<$F���.�1�<ϩ�7�F�q��͢���[Ʃ�~��l?q#��4t�L�Ht�y'p-*��: ����2_}� �Ղ���өc֖[���Z�;�1���Uo���A?��CC۪̜x��kd�?:ZW�H�u��;��}�џ>�2S�^���%�gF�@v�w%1�WfK:���Z�8���e#��V�U�ZX�绋�������3]p!�9�b����o��S���Q�$�I[��ixox��%���#�8oO�ȟ��l� ��lRA��(O�d�o�}�)Œ�P�kttD��j�\ßQmt�`��8NXHSr>&��!��^\����vX>]s�?��V��Z�IH�\��a��m}�cNn�!�+q�g�"c�~~%I��6�r�A]�]ﻹ���if�g�7ˣ\
����CŘ�}ԣ��mm�-��j��3%1��q�w��ڣ�K6���$�ؿ�@r��cRP�o�7��/��^3o����20=t'����F�u�d3
���|���:�`U���(�6uqH\`l���!���
J �]�:�7�T�n?���we���x����:�󺛪��6f��Uk_�@���<Y��E!���|��A�8��HI�Xq��g��Wj�bn�fX���}ɴ�m�O���"|�����>;a�7%$P�E���K9B�P/�G�B.����/ν��Ca��p{*	�GJ�4��8�Ǡ��>��wk��a�h�5ԫ���=n(�7c�E�u�˻°��-�P/� �F��hv$8�% h�n��TW7�p�$*��Ry�6	7>�|���`�M�0����~��99�얎"��eOS�b.�?u��흷nRҤ\ʁ�t�%c����C3a7����dt�@̉����p�h)'?DV��L�Y\-R(�
���$�Y�0�p����u\49Ϛ�"�4%7�:_�g�
�Ý�i���׽��Ʝ�z+�pX����E���l�R�oǓ&`�b��Q�!���gsR��#��CnP�%���Rp�^��eӴ-/w�=�Bx��
w��e�!N��J]�$�fƀ �)���O���/'	Բ������eI6��í�
2�1x��H��u�f��d������U�m��=�8�,�/�k��5�b��K����D3�9�f��`�|r���g�f<�����ۡq�x&����#�.	�Ҁ��T����VI+ƈ�?zF�G�;��_w�_Ɔ��嶎��8a��8�^F#�)�7��\�|o�� wx�� ~>z�*�;m�^�/�X�$�ן��ء�6�?,ѥ�q��J�����4bݶ�?d!�o��BN(r1��蕭,������c\0�+�8�c;Oӟ��g��'!j��f]���Q)�4د0-���H�(��3���iO�k���㉇�
��iΰU�TG� �}�P杮�NQ�n�ɏ9�3v4�uji�К�|�\L�ZCNh�d� ���%P��uҴ�[7�!i�`�=��\�z(y����� ����+GM!e�	��k��ASs����>�C�;pz��n�;�l"@+/b*�c=���� 9%{B���Q�	.y�����=�t\v��|A�_w��G�a9�����?��u�eStvHx�^R������5Q,dI$�4hpt+��i�ꋕ�t��+��Y��0�	B{�c�?j�L \m�(��k*+=ݗI�ۦ�_�UЧV�8H*&���Bʠ��<ʍ���A�y?��9|
١�
��5Z�*��o$+�獯�-�fni�LHy�����ߧ��ڷLV4-Ni�u�!�/0� d�����X���A��Z��AeQ��zGC�ک�o4�Όl
�N����X�t�,s�F,�^�d;6�Pw�S����Rp$�Rݍħ�o80�cj�b9
��Q#Y6�pG���nIi��R��4�w�?���u�&��|Lt���Tc*���$X����~<d>%2Q&��Ո�峺�a�˜A�����'=<�"�W�=�pyF�[CBG��o�h��d�[�{�h�G�-E��p�N�¶dv�;�.��� �RB�t��͛=#�C�@�����B}� _S����f��cV�}	ݽ;^��ǎ�h�.E,�V�X���bfJO���0i��L���D"�����mW-Ö?	i�"���q��GB�ٝ��z�6��ε��&"c�r��75��8׭D�%�uTA,A� p��8@��u=�CZ�	��Y>�S����J����n���kH����od��yTm�2n@�<oA�P�D��.��� h��$0��rA(���S�2e���"3�X�7'@K6B�d��BTO�٥��� ӨHp����Ӟ6;i�/��4�B%C�Y�`gQ=DN+$q�Yz@�wV���5��N�-PD[��t���q̑���d�+x��B������zj�C+�3Xq�Cn��@Z֕� �]z˛��%�N�ԗ��f�����$V@	e�ǘ������{�|E��\�,���f��;ֶ�s{*�'�+R��fAf��Β�z�%d��*���e��jш��hLq�L���j��g��a�5�5�(%�ں	I_��l)N�$�I�$ҥ�(�*�m>6t���d\g�ة�[�Y�iN9�S����P9;F����LrOi���>����A�D�����?X_ޑ�zB� �Y3^�������/��,$Kz&n0�V�0����G�9��E�^(t�i"1��5*�!J�K>Wk��q������5����9��xf�Yr�j0���͸�h�)�i����Z#���9�'O_��ը��G�V���+֝�LBv�*s�3��i��.��0�<�s�t�X�3Ny��]���k{���Q��jQ�4@��z���q����Ŏb�=�G����|���UYu�\�
�6����I���s��9� i�ֲ�Hko}����y4��wv�|nq^�U�4��4�v����q���[����ƭF�����	bM�Y.�*�x4k!�b��m�ǒI���&�o��h]F�!�0��]����c����k?qgS�D���c� *'��YI	g��!~Á��ȃ���#9��e�xq�/+N4����Q4L�U�Vqʡb�����,u�s^	[]QͱGӯok�t��l2	�*���e^��{��_ɉ�$6~_�i�+���X�P�E�w�^[V"E�˟K	�O�?�+#_X�t/z��YEL�켦p�G�F�3u��1�aź�t\�w6/js�LX��_e�$�U�e�����y�O25���@dM;k���+�t�s��?3���@@�+Aʝ9ǣ0jZ7�-�Pv�BǥK�����EACbτ2�*�-bd1G�R��S亘R���ȝ�{�.�{T<)����z����������[��<o��I��F�ց+��a�����j�u�	�kc�T��!�9p4k���+�܌��ҹ&/z�`��-$$�����L��Fx1Hc����ۣa�;��?@ ��,|h���H��p�F��n)�ĩ%�i�q�9��mS.2����q"v�j��5O�~�w�B�గ��d�3�L�(��������Yt��󋕮��^��������',�_;���$e�W��B1z��>�('=eߟr��V�|�6xkZ�h;
�T��{%��4�e��V��/2iNeF��ؒ:E�V9��El���1��:���H3�()�Mv���9�-ݔ�\��|���}joa:k<�4("d��;�ay-�I�Q!c^(D�%�}�Z���-
�:�N�R�����j�V��ɂ��	k5	 ��[�s��RD�S���͵u�=�V�4<�кVu�2��U,׬��wrY���09���	�	�X�@�/n�3gqC���9����|ĩ�����(�Pe�Jғ�DfN�:9��O�)>�Ù�};���r����6�5�_	t�PLM��`,q����e�=_��b�d'�������t�?ev(~n�?�F�hL�n$8���גqQP�9���m]`�\���J-?Y8�r��5�m�W���u�ܼD�)6�*.Bg��»V=o5�䡜�Hֱ'�C)^���e��cVW𧻓�ѲI��_&��qz�$4N}�c�\����[u�C7Y1\�4>P7U�)w���L�U?Blt9K�F�p��<���wA+�I]�n��^z���SQ�% �uI"q��	0-	!fj}W�Ԇ*��PUjG�M�7F����W����A��K*M�Q)�D��W-)���֯9��_�H���(��B���#�77M��,����;|�l���)6>���S3g�%؟6�4���}~p�ϣ%�L�)�%�:-� M�:�\1>�Vv��^]�������� o�gu:Z���-�s˷Y2���;���N鳜�?�}t����K`��.=�a[�tg~s�,�}�_�w7]:���Fq�R���m�;���]a���фVV�k[Zg^�M�p�k�EnM���jF�4��z���c^��5_	 �<�8V�"'%�Pb��#���B��` ����Fсx�ZTw�6wE�Ww��~��*��s����z���p:�n�f��nD���Y�X<��l�4�i���;�j�M�9~.�N��~d��po!D��!H�㇉�CI��V�rh2�e,'U`��.4�2X2S���AP���]��6���η큺��=��J��$04"iW�h2���f������"{y�}:]�k���@�6<��_B�k��P�P��I��8�5��L���)(Q���V%ѻ�-`��~B
a�P؈�4�A%i{M��_6�fD3��y�I8{=?�T+6��"i��t`+�z^Y��@��r�=RM�S
j���P�v�lLem�;�h���}:,�vJ���V_}�v��	�L�+,h_)����ncE�*�r���a��1�Wqk��Q�>�o��3���۷��x�͉h�H(ɐ���WF����wvfX�9��y�w��U�r�.����1d�Y|	�Ǐ�O�$��s[E�����iTi�#�GR�<{�x�ʢ)ӌ�m�0� ��M������	g���%��h�($����PY��c����x���p�f���p��γG0ä�N�A���Y�:<PSsЅ>�1��3�i�\�E�*��ON}�TA�x�?_��]�{���6n�"J��Jt��uVWO�%�X�k���,8"c����:e� �N��A�DT� C��L�x���wf6�B,5r���|ꆼ�'�f��P �k�>ږ��[2�u:� VƮ�i#�=v��E�)�����t.q��g&��A^���_!OSO�R�c�'{y�8� P�[�_8�vI�o�i�e�&q %��z%��I���CMA� ��`��ʸ�֔�L���>HŌS7 �����|�I����*�̴��4��uz?�{uc紏��Ul�M�%-��Quxj�"��c�a�hk魖�,�+����@c��c�Q$?}���N+�2[̓����Y+8*i�\3 ����3�RɌ%Y�=E�S*R�'�?O�}-��N���?.(�7�+�T�o#�5AQ�v�*�ܘ�U�F�DB|�N�S.�K�x�l����ʮ��)�T@Cmd�I�-a)u���;&[�O��"�4*�{kR�Y�މa%7:�h	1���f�Q�����v���E&������qæm~Ny���|۳�$ #��ǵM��=��;N�GfM5Hռ<��סV��	�e3��_`a���˫�/<`+PP,$y^�ȊPo�xl�,_��6����A�$w?��r��	�z�_�lX;K=�1����*�X�k�`N��Q�`bZ����4���iVB�����#�4?�	��,�<�@�X���ˆ��ci7�Ή��	�
�J��އ(���� ��z�nsHR]t%�T=f&���c�B���%%˗k*9�S���$~���u�����!}��WcT�}���-�37���(�����/�a<��0��Ό�۫�Y�(d���a?䶿O"�׈��DRsm���bR�dg��Y�B�u�i���ȻD�˜��M%GB���(�f,��`�x��)�)�zPPMZq�njƽ����jT��Z������������Z�4-�v�ܞx���P���e���5{��E�����g#�ۚ���ֹ�\U����������4"婄���$���t���I5��(y�^�Fȣo�6>(�+��X����mS���m}Ʌn�W�>�i��*]��4�ϳ���������2l\k�M�~y�'�7H#��+5�Q�T�g�}ujw���j�1�
Nqa���f����"���'qZq�@{��[�1!W}����F_<8D�)D�1�v)�%�Y*��~�7/��n��rzB0�}��M�T�n�c2� PJ ~���{�s��$M*�����㭭}�	�С\ih}���N'+�J<���P��M�ܨb%?M�C�:WW\7��кY��Dr1ӻ���d:��Z��V�V�{`�������L��H4v�J�#�+�0ȁ���MP�d�u��<��A�Rmsπ=l�*�e dZ(�f�]p,ezywā��~^i��gć�ϫ`s��ˢ�_Y�S`�ma}�P�C����䬃@Z<�3�lɺ��s��	�S�;R�02!���@2�L������C�6�8�����-6zC�V�|�*���r_�f#�VB���|9~���є���|��?�w6�̧��C��	@���>N�}%�c�մ���tX=�˧b��n=���'�"i�#�!*ה*ڰ �	+S>�n�0��Y� C��W!Ȩ&@ځH�v+'yO꽊��C���a���KN�ҡ�TZ��#E%Vc��ȷ<���*Ht|q۹T���j���j������KT�����'H�-:kp ���6��lm�}��5�!^Ū�� ㌎8���փn.<#���������ID��G$S>F"����6���m�"���t���.mlr+�CTƶXy.
��1bE#���v�8�벵�Q��W��B�؊#6v�n\,�i�Rq��U{sf֎_=���'6o�"��N�>��XRWw-q���Y>��s{ئF�f��C�a��4b"f{%�ɾ��/�a2�%�U�Љ����A�d6����=��.�c��,U��D�^%{��A�ͷ�]'�sv/���L����
��;����?�}��\T2BPə-<�$��V����1�S N}��W!� �ǘbm�wŎA{�ڜ�mPQ�֗���)�d�@�
��Y7�q�K�.N�����n�:q���ւ{^>�B[ڳ�Rφq�B�����ڟh��ް�d ?j0�>+�:��s�{�����˕���_>@����Ζ<I�Nmt)ȸe�?E\;w	������ԑ!v�;�O_�p��J?"	������0�2��G��XE#�m�6MO����k��ۡv"g\م�������e$z�=#��{���.�yFQ��u^"2RDwf�0�^b��a�����Hf��"���r;��&���F Y���M�2~Zmh�ף�ɦ�;��8�2�iiL��ްY�<DG�-�~�b�[<w�Y���LY���p �����3�8���Z�Ch����¥��H�t�{��@
����o����8{:��yqߖN����KK�Y��H�G��[�� ��s��W���M-X��h7M�?a��{<f ���t�a�W�bp�۟�]��s��h���k��O]�(<%kV�R��� ^U�M�}X_a�@A��<��Z &�����	c�#��w�*��۾a>�B�TB��>��q�x�m��J�~ƃ��JL6m������@c9�]�V5����fR�Ȟ��E��c(� ����y�(�`%{�h��<l��\wS7�X�-}(�!��&~١��l#^�Ǩ���ok����w�V�A�!c�@l˷������v�52={�^]�?TY%�k�E��o���z�шc<�j�n���1Z+��{FvlGN��ߔ;�n���kT)^κ���k�kXl	��%��MH{]�]kg���Ydeý�M:[gَgY�"^Ɠa��2��qV�_D�f���t��.�(0f+c�8`&��©-�v�Ă՜ӎ�I���l������mS�"f#Y�X�.,.�g��n��S���J��gB�i�H��ʲO'@8[0A�!�.�[��En�Ps}x(�K3��o�{�^_�v ��'������}5&f��ء�"�w�P�W�O��,|T5�'�VA��G��9e�%��ۅbZhv��]���'_V?��|d�C�8Vd�R:G;R��9�a�^#>��O���p��CM����@��h���`��M�(�[���&�/#�cJ��H����E�0H.ZY1x=�|ĉ�5ʦS����b�7���m%֔w�����R/Ar�x��,E��C��_R!���(@+3Tٴ?�R�����uu�LD1�����lxZ�/���k	�t�7�"���2b�*�҈}O�W�!<
��M�!P
��fԿ�^M�(
W:A'�����*�S���6����Y,�:;�GB,_�ŴS�a`�H:�����Bs(P0ϑ!X��Q�:�(����[e~`�W�.'W�,_���ދ ��'�	<1���ǟV�LF��Y��*呲�$D�Ķ{�|�[��`�tC��cUbM���j:=�_ym������y	\��l<	-�S�.�Þ@W�$�fH8+��&���a�f�� ��Ln�E��PHB�֡vh����X��1�J����u�7/aN�1�W�P�Gk>o��L�����5���u�Z��0�����ҩLL�יɒ��FR}�R��7L~z��Bp�:��C|W���>r���P��):��L<|����an�쯰-�1Ժp��6�VcL��o�b|h[f��(q{�J̌��a;���K�k_@���{�kN4U{�ቸ>�J��Bő׽���c�JZ�{���YOzk 9��K'Y	�G��*����Bc�$9`M�m=�B�ߦx֍o-zbG���K��1~ԞOٞ˂Ό�%Eѽ&�]ٕ6\hv6l�.�Z�-B���+��xC��SH��[�R	���X��d�xېv����2�3���F=�������4�~K��#�F>��( ������ȣz&�_y��]f����I�RS��)}�eR�[w��^�K��Aۆ�6*�\ull[��cC�+]�%в����U���X�;�0 ӥO�:q�<�ӥ30V?��M�.yb�Kqi��Mm=���U������q��1�O�7�+�fI΅�Z����7j֧>����C_�6�E�
�l)u�l�{��!��kb9���9H�e�����"{�>�WR��x��Ď`��fo��~|��FlHd
B��fkɧ+���e�5h�����$�����(�&��%1`xk�����M��߉"��+(* \�h��!,↾z#�&�=�m�7'�,ɲ7=Y�v�']�����:Ή3b2A&��-��#TR�5{KĎ�����5�����=ޡ�mA���,>�]@&�545��>����gV�i�q+5��>@X������L@"z?6L�8�?~��)S2���UG�g��`!<	���\�I'��.t��j:#l	rYOgj�i9�s���l)X+WJ���37�U�� Og��xkI��Ϩ#��,R��q���){9�S�|DeH?�Z�Ӈ�2��/��K�u)'�� �K��K�r	��M&����ra1�&z�Q��W1@q?d��Gj�v�[^F��ߕ��6˛I{Љ�$,H�b���Hΰ�<VZ���+^iI7��C�X�=�l2��EwNA�y( ��d�i �h�@a��I�F,ή}��!ս���_��"�rv�����2�����~��n��kƦ+�ѱMr�n���&M|k��raf[���)��������4�>p*��=�|�z �s�X|Z�Ή�\'�k�s��v�!3 ���ȽUO�P�l��-<��������S�rY�6$e��Cژ�j����9�V���/h��53��M��:�q�ל��9��N�ga׷10��@swH@'}�Q9A�]I�S��Ror薞�f*�տ��/���C��.� 2H���	f�����x
_��JX��l �&|�vk"."�_\����:�R)ŃF���uЇ����jPr��)m~�Y�qt���L�W�^�������5���=sk�C���2]'Sa��*å��S�TA[��_��bE�����q����<�~KӚ����X'���y;K�p��-fO4 d]P'J�G_������ڡ+�{��~���"3���ٕ
��8j����o�6�����%�Ѳ��y�^�
��� '
�|���v.R����Í�'�"R��H]�8��HN�=���|�!���Mu]�Ȏu�:}N�kg�!jyLx6�l]ت�D��R{0�qEp�t�i�w�mB#��?�'t���u�
p!sY��S5�HJ᣹ ��;v���P��;^u�*NE�������X2<�=Ȋ0�J�^Q�&&XJ��w��ߨ��%d����5QB�����֘	ڭJ�'_{c�+r'�A�[L"�b�^˸MS��i��^��A�"GNX�ᅡ�zoݾ�	e�62��/���!N�'9g"7�չ9�u
W�M�[ �Kz	6
��`��u
���?�A�6wP-Kr䛬P�C�1c�T��g{��Ȱ*�J_�৓Y�??�BE�H�Wh��2FK%�h��˼9�v?��ӫ_�M�z�+u������=�5��26�
�*JI�A��۔������D�Y��{�CS"B�����8�,�^ �r�9�TLݓէ� K{*f~+������C,U��l��;��(�L�zy_$�u"{8텚V[�_����Nt�� �>#�Kc|i�3C����e���(�Pf9Jo)��	�����;��s�ŕC��'��M���Mƣ0�m�fj������+��|�i��cV����c�Z-����{�����W�Uʀ����CZC�k���tWhQ�6꜋��9р�M��}<-@39�t]'���5����eP�AK��L��ïQ��%S�t}��Ҙ�h�s��P�w�]���������ֻ�J{:����yà.�h9*>�ס��LpK�zxݗ��lwI�Z�`�]D���+2B�R����Y��j�,����e!��(�?u`B��b�nͻ�/���C֮��v��\��y~zaۆ����<�� ����a;��?wk0z5S�=Lc�?F�Βf�C�!D�b�&م��s���eo�2y� v 	�BH��� �K5�4l�6k�¤�ג�~2�34���2�(�CᬦG�ߡ��!'��F�5��H�_�F����a@�� VA|���p�*$J$D�z�+H;V8C�Z�M�SX?����%��+����똖��F�m�`[Z0���Efc��w�]T/D.;�b��b�.����j�5@�[����%�g�"��C��>�$��5p����%���V��&5^eG䧾���Bj�/��̜xn�b�  ��R�h�T|D��'�sd��ڜƭ�5���03��[a�@h�����-�98u��JK�Pv-�=�[�)Q�5���>T�1�j�B���y�w�2 rZ	�{���O�FH4���3���%H�L�4
�i��o�h{{�a��ff��n1f��"��� �"�֋ݱ��W,s_m+=�?69A��e�v�:����̺��ZZx�k&uiE��T�ڈ�\HC�G��.��?؉
�ۂ���o�o�\�e�2p������V������8�Hm��	[�
��`�*���)�� g��Ь� k��*K�ټ�R+���6�޳��o�M�O�&���P$����*�jRe�f��8:����;��|�~��ތ}�³�oȇ7_���N�m	�Ri��(bM!,�(���j=�Xo?	7.���na�d�]�r;�؇ji��	���`�E?@�������-nh��o�d- �8t�G�{3������$*�2�[�}�on��'Rֽ��5m��������kpO��:83$��5
#[�]H�&.5�H-��u$:,@�}���7���<m�҂m�%��cJ�'$:���d�yf㡌T��e�r퐉=��؁�1��,(��)�Џ��*Bb��yӋ�P�j�HǸ��!HNmH�m�5ާ�����3._����t�{��ܘ�f���Fp^�w����T��}�~R���)xU��!�"Tl�߃+`�wk��P�u'���
3p���~+�7)��Y',�Y�� �q�%ZD*�e��PK�;V���HÒ�V:ɒt���C����$Ħm�4�<K���۵\�-��^�$pqj' ����G�7����F�3)��G?_@��� ����b}j�Kx���aɆ�y�d?0��R�̝[�Y��a�Z`�5{f�R��!t{؉	(\}v藌��6�: ,H�o�� u�p��j��ZW��W���y��Q��UonV$Q}�EԌ��'�Y	טo&�ٳiN���ulr�L�ʖ�rt�Zl�x04�5j��:��kD����1{�&2B&��w�:\z�8����V�Bt�`�2�S��|Ʃk���:���7��DjI�m=W3��e�R���x2#���0R�K=ĥ�+�F�m	�ohټ�S�W�aY�U��V��7�|�����(G;�5��c�w6yI��M��� ��X��Q�R�J���X�:��E^��}���g������Ћ���0�̸c���P74`������"c˻X��h�է��L���()��IT�����4��S w��b��SoM�Q�OR��g(��oS
`I��71�@��l��R5N\}�5�����'�j|亰 %!���Gç��$:��ܒ	�Eځ��{/%�G��c�R�̝zID	}n8E�.�R��x����,�2��|����.g�Բ��^�5k쥅���q�ݵ����>�����о��k,��$�^uR2
7S�fJSR�db4� �5$����k�e�ք$��	��^ށ�䤆�Pc4�K�a���7׸�;!��B�1�ʵ��0�:^u�����ɣM�D��Ԕ���9����Md�ޣ�B��x���Ҧ1L1���5[����iP�	:��5��A��d���B�;c֊��Я�F�|��I�
��C���*鳕�;�6�Y�5��N�'N����6�1���]�\+��5�!썈���Ϳ�+�� ѐE7Ir��j��^w�t3��z_#�T㨞Si݃���nČ�p�6Bt�|Z-$��F�'��|�
X#����ڰ���ƒ�Y�L��x��e1Y�NyI2Å�5�XަG&�5�׏��Os�����\�2CJ�g���!��6�4wa�N�8�:ust�b�y�H�_Ա��ra�R^�3u`��v���tE!��l!Q��x��I��(��q�Lշ�:��	�A�)�xa�`�/�{n�\�r+�[?��R�\��[$|���k��E�W��㨞&�O<a����F�#��;-X����q �Hʸz���	E8)�ڵC~��2i���&ϭ4^�9񆦝��X�P3�^��a}��@��A5��w��w�����y�So���h��A���z��=_�HH
v�hKH˱�{�<=���li5ʤ�;7~��+&�*ޒ~��6Kp� ��8����U>?d���w�h��!��y�~�M_Ӑ[��+`��׃d;�|�8M7^�i�P��8iP��	��	��&R,[x͖��O����Ԧ�S �B�V�[X�g�M�Q��k���ad%�d���p���'�@a�p"�C<��kg̱�X�tK�^� ����`9�0I�C�3%��o�X������V=�� �UI���f�����˸��;���g/[�����z��)�.��,}��3�N����UE�!M��[y��c�G�?z�������hi���"<���e��G��p���ӟ�J7s�F�JA��+(��X�}٪����j����p�;�2X����k�� ���e�}���s�`[�t4�z'L��|��ƴ쥅'����@-�K2���]n��նa���-����q�Z~�fd#O�ce;ŉ��6�+H�'�xG���{�`�H�i��i�P�yh��H�d�u_r�P���1��;��/%�\WH�v��}*i]��B�\�����Ȫ��+1�ۊ�$������a06�*��M�Z(9<w�g�i&a卌�耨W�IG2~9���%g�ݦ�gМ���ʙb  ��WiSzX�M��l�-��8{`v��TBF�&�%�>�U���W0\���1`�H�Hs�:;�Țt�2��H0�ڌ���5�4s�؊Kp˗����@7���C����8L5yz���>m~$@�#.���d�ql'�:���YP��mK�&2=���kI�<]��`��>G�O�������%�#���n�V�T���C���##�q\6��/V$�������,o��o@�f ��DAZ����@��<[�TҒ'�	SL��6��xu�T�"�%���8���a��3w��`F�f�-�� �����+Sժ;)�v>x|��܊U����%09�-5�Gq$�I9�Tm��SXQ�o��	����Y�:�D�o��s-�P��fדm,��q&� ���M�͠U���jS�c%���	���t�sô����cd�tKA��=��;�ܘ}���eG��_�>Lo���^`�r�4~xyU���FA��G���&��Ʊ)�?C�EO%J��ǀ-;U;����d�+E�Zod}bej�($|Ž���\�&�f�i5*��<�h�d��
>"2���atR
�6�����Q��]�˃~�p���T+��{;�:�%aG��Pw\3Omt�`�&{݌$E'�������cL��b���s�e'y����rp��G��li���,���I�"m-�W�h�>�g!��e�ߞ�"��~�l�0�	GIv�2�k�E*{�QG�%������ƃ����h����U�- ��nB+���s��"y��������u�o|j�>K �A��ز�2�)D�k�T�m��i��Ն�0�cv슾Hc�(찷0�Ϛ�����~䚬-8|ز�P��o��P=�����g�1��?+^0[gT�nd�W��q��z�������~����HJ@8D��!G\��~N�xḟ�������-�W�\��pڢJ㭙I2%y7��2��Z0=������^���Q���;� ��O> nXF��<kԫ�蛤�ņ��ApcK�!�쯚��.�YwT>����"�Kq���52�������r�9�f�o ��Ũ�,y(d��w��Pc��U2^(CN]�>��uKD�*��I�_���qu�|����ܿ2���ryT�'S#w�b�v�k/��A*ڻ�*a+Еx�f�*��G3�"o��� ����-��8d
*i��������{$Lp!��K�9�/m�.R��jo�׳����~w��o"
�Ve��OiA����\}�� �B�@��VUR�L�����@ �z��������UF��w_����`s/����hC�~��A=ɀ@(��n������H���5�n����MV�;]�ӭ|aU����1���-�h5����8�$��9B�pi���w��L����&�G�q~��"���.ݜ��2C'|Y�tX��i2
v�m�=�N	_��B[�-��7�z���$�/�V��ߚ���{H�*�Nh�I.~ާ�"�e��9���#bd�}���IT����p��:DRq
xQ������v�������7};f_n��#�W�lA$�#sXW���qX�'��$ ���w�'�7��I�r���/\b�*Y�T���5�-�����+��@i��
��i��@�x�Rɼڇ!Ŷ�%b�LTP����y���m���:l'��?��5�ʃ %ԕ�hLg��������j��N�����!r��;��2Ĩ\�i0�{�T���.嫲} �Ǖ$=Ц�g���(�-�xS+��ƶ@hgg���q�q\���NM�K��Rl�1��X{ly�M;v�F����GR�PP�;ۡÜ0��]�q���2�g�$�uB��p0RX��^O^e�K��V��%:�ki,)�T�|���pE�����:+�`xw��Ǵ�!瀉�9��_��Gt�f�b�}�0E���
���G��� fI"����@�r"� T�|K�ah5�/1� .��P�Ǖog��9����r�Ӓu�n�ufЄ��g�$ݺ�<M뜐q�[�#[���yY��VF�'���ݙ��گ�߳t�9�cB۲,�����*N�U&#����NH ���jK�2#�������ib����VV����ど�~y϶�������>�mꡬ��
�N	�u���K��*s����H��� �	�<��7�7h��)�y�R�e-&��dYoMM�ʨ��n� ��_1&O��KETb��eUW��|�!��˚���j�sx���F5bH����x`h}���y��˦�"�Q�-jZ�.?7Kt�pv�\K�ѯ��A�n�:x����0#��X��w@���9����=���M0sJY�����1U@��7G�֪���'s�S��l�D>X�-��q_�,Q%��������� 7�Ю��MX�F��ח��Z��5̈́�_/1 ,1#�ڛ�>:da0�����<#�6�����v6Y���Z��C1̲_�SƷԐ*S@�$��v�ꨲ�]Ɨ��:�
�iQ(��ƫ2^S�7���g�q�m��#���g��8x"o#-�[TZ�fl �b�+/�۬c��a���R��ɦ=��	�?�jh�+7|�k����mӚ�^Hfu-~�Bp�6Aͅ3����r����-%o�G��y�k#�h�u�Ȣ�w�^4"�?�b�Թ����峞�#�������GXp�$=)�g��24����J�F_1��#2�=1t ����Ԧn�ZK0�?f��5�;:��<ƚHL�f��K@?�#�!�/�,u "cb'�;P�>a0�H �>��ϔF?������ɫG�/ɲpG^���x��c<}�����;�@�ƹ�_�h~�_����B��ͥ��h���иC|��/������8�-����:�M�{�:[]��*Һ5������s�emu�er�&��=�o0�]gy�H4��H�ט�_;�>�& ʡ.S�i���n�0��Y���]��\�52��6�;�|E��p�&1�RW�"��@��g�8������Շ0M	3���\�s�=[�39��R��	w�ѫȖ&݉��5�hP�C7����_����K�M�t�M����v��(��쪩%�"�_��65��hk���Sx]���P�@a��[��$�d��#����bӉk�Se^�[��OKf�7�C �����N\��[�9$�y��ђ�쵾w��P��"��/!���ăy�9���4�a$��!BFF��{�4@�
���$q�m'�%�9��ea����";��W�h�Lw����sK��� )k�N�V�-ڭg�GQ<t���̼���6���+]��,��4����%BK���v���L��1�Hzܫ}���87N}�����;�"����]���&c��n'����֩{���/��͹��	6jS!�Σw���s8S!��c�~��q��!��64��D��}������ ۏ����'��l���\k3����A�!�Mk�>���v��G�cR��ME+��.F�6>�������Yu��_�Q6
O�[�����י[�$ר��S$4�NK6V棬�R���3m��&hk�v��o�ʡ���sQ�h]��cvy|r���4ן����g����_�k����H�����Y���V��R����MZ�lޑ���UU%F!��&��
���?S�N�u�G�����}�� t+�
�S��$��|>��,o��i�ú��
�,�B%�\�
��o`ޥ�Z,�0(���e�82DI\m��B�<}*����z�v��lz�y� ������^�!d=P�Si��a)r#w��\mq|� x����;��>���>%$s�������?`!����������.�n�����,�@U���a/��:�'?:0���z%�΅6����r���(�v�3 �ڻ`W��@Ā=�5��B�QOuE�c�N;��=�%wE��0���*^�� ���S�	AN E�w)2����@�j,N�@$Y�Vۻ�9;l��c!���{���C�����.ᶜ�1j��A �IƼB3�`/���Z�o�X�@Ǽ�DV)��|�蔲�!�W��H	7⦯�`��>��6��u)���4&EAҦ��s���'A������߳��]fa���2-�4ϓ�e���٨7�V/�pU�3���)�ӻ�; o�4�ړ���SS�~n%����B~��t�@4��P�7�F�o0<x���Z� ٽ�O�d�W<d�����Fb�D�..mM������+k �Zٙ��)����7�\��<c��12+�g�ǉ? .�'9� ���i����.벐���|/�����$i�@K)�S�%2�n���!�A�7�T]���ul���Q����Z#�Ѐdу��u �ͲQ��S�F3�ᾠ
��w�� ���r 2.q�lE�,��i�ˤi�����ߌ�@M��JHhB>x��c�P����=8�<��8�8�f֐����s�<2�
��z�#�kߢ�i�kp�c��?H:�K��߈�E�pn�H�\`��e��� �>Lebm��U��C�:;�orө.U^K�dU���A�ƈ�[q\����O/���nok�� �o���M��ݍ�K���'N�����F��B��;#~m�w�z�ZB�ё;�vM�������T�*�t����\������� �\l�T+{҉����w����!X�R�QX('��E��Q�#l�Q!����l8�)�9-J��݈�80e�ej|_�X��������o��0u�G����p�@oN�����w;��_A�q��R�kɷJ�9�a�i����2��/�����yh�M���k���g�HL6u׫J�[��0��(0�wV�;1��!����Z��GB���;N������ٽ�zX>��{*+��*dx���N5����BL�8Q~�`����IF����7}-:N/�B/����o��ϫY1���Hsg��~��1��D��i!��w��n���&w� ��{��Զl�p�ֹba�ǻ��52�#������C�P5s
���;�.�4��P��.`�� �e0k�/[���V���đ�����N|�ƒG��JH�4�>�B�꘺y��6��<*(e�M��V�
�W�ƚ�J��Q���8�R��D;tl��B�2�[CQ'\��3-l�X!kx&H#�޿v>*z�!Э٠�}���� 9���BA,�Ғ��PRf�N�C���˿a[76��*-ɴ���v/��!��qb��Z�W:ˈ�جF�&�^,yR�R���;�e'?�3��d����u9`˲�� ��#3�{��rIs�H`�-�0�v��0��"VƾKݲL�O�}�F��yw��`;ό�sZQ�
�v��1�r%�Qf}�kP?q �n(`ݜ1��/>��1���:����;���Ef�a�zDu�*"#��~�I��J��X�M��4�Z��Q ��fl8�>G�p)�I؂}C����2���lUE��;-�<n�d��8�T	sB(u|'�ݢѝ�^/�G�<�rBa=��2�[|��t�=C��2yx�y��i-l����c)�\�_d�zUr ��N�32Tj�z��@$۸�q���&��j>a�7#-���<[�_����u)����u��Ub�=�R��Ǔ�jď�D�� �G���E�D���g=���r'���K�Nd&����6�l2280/��`ǽ�T�粮�v;De[z��)~�Βވ	�TN���"��/Tw���G^���֏{�H�I�9L��,��C��_�,g�m��C��-Ԣ��WL�]�A��x���9 LJZ��>�d��{aF�83`=Nz,*�tb"��0!���\m2O+�����w�!ĵ�'|��V�l
����R�a����#���5�� �8HM��T2���q�c�J��ׁ��qk�!�g��
� h6 MI�N�Qsp?i����/�
�I�����*텁�� �C��I|�1�|�3��00��V�A�
p�ݳ]�QbU�9D,��S�o@��l�{w�����,!`����]'p-�N�*�םЙ�Õn_")���&�P.��"$���<�)�h�	g ��12�ge`�u�N�4o� �@��!�<�	 R��@�\��aC@����X�2#�P:(��V�[�Y��y�@>��M���{l�2*�_vO4��]�Ә�5p�ӝ�w�lS��������� �����0��F����cM��z'�	 U�|�����;K�����vHb��6^�QM�]p��W�w����C��H�{����3b	�B����4�Z��^'g�&�����~2��<�؀�� ��ĸs�4�skPEw�o�ɖ��Y�kg��&�a�6� �V��{Cd�m�6@	8T��޾e��2c��H�y��"�C�Wa�ܧ˓F�n-,f�i,y�xj�9_�j��J����h�l���V�rT��^r�;=�p��IK���e_Hc��[H�m��N��	 O���c���c`��$2<q��7�xK2�L�T��d=�����˒X����z����<�5���_q��*D�.��A���3m>1"tA���g͇�B=�v���a4	�v� 5��YB8����*�c5[~�|�k'W�m��K�ڐum`%Iћ$�W.R���*.b�P8��#�4���8��#��)T`�k��	g:wɸ��շD���3�k�����%�Y�Ͱ��`��+��Mƫ�������'�r\+to�ɑ�7c����o#�"�Ʀ�JKHC-��#��iԽ�.�ɗ.A��Ou<�c ���A׌��'��B�iB6(qT�~8>�;ڨx�m��R��O��:����K��M/X&3ob��+�\}�g�s����DDͅ�m�.wv��y|b\���"�D�q3��Ǣ8.��� �%)�K��7�2�Y"��T�䰑�(������<Fx��u0�H���$<�p�@���FY�n�
s+R(�_ �������8yw�g"��������W�����霼:���1u���@Զ��z����g(W������p�Ĥ���`��߉'�� �o��<P��lRh� �b q�Ƚ|���@����k5�D�ĺ��.�*�]`Q2j�&�{C������[�*��������8/�����'��/b]2Wٴ�6��Րo�iSMU[��2Έ��u�b�R��D�:�S����j��܉4r�	�,����9�_f���bcrž�;��+�V�@�,� �U��0rf�L�L6!~�p��و.�0h�" %��|b[�v�od�Qm�rؐCD��.s�7���p7���smq^4ӈ����c��o�$ �Ni�*�!�e�#�a��s����Pr�>��D\�r�b2�(���Lm��?�3�F(�9+�b���/�V�J{�D(���^�k�N��F���.Z�{W�W�gKF|��\vRr5�9��m�\/Iη�\�]���������/9�ᕇ�6�o�$%��Ic���?��"����l�#�1}����:�Șr3����5a�������v�lWg��2��218��w�At�h�s|Kۃ��}ha;�j�W�"m�{���L"�/�|�ǆ��:O&SچXk3�<'hK�
�Hy����uW&h.&�M�/D�]w���{�[�|�ZS$���_6��=��jwS�����Z��k@�1��:��=?�C��TM��?�}�wN�|�Uh&/?C��+���e�{[Q�Wo�,g{�.q�h)ئ��U��1+5�8W����8�	Kցo�2E`���������/qg�O6
C���jfN6���8�ibm�	��l;�t�h��B���o.�s���]f���!J�&�R��"�oX����5�pe��U��_���8O:�.�G>x^s9��ɢ�H}�2w�{k�a_OŬ���8YL8��̲6"�v�:���$`��U"5
�Qw;��t9x����V�d-���w�|�{��'<#m�HN�1U3g�z����Yp;��s鉨A x%���0���d�d�ߓJ�^����a!��-���[�S*�zH �#3�,��2��}��Z	�H�
�����Dgd4�:�i|g���j���L�9*\�BB��ۣ�;P�:�ZVMZ�R�6jvQ1@5�DAT�[%�ə2��BJ�$b��D����쓎FDS��nT�j�䘣qM�2��"Af�ha"�����pV:Th��&a$_g�W5V �Ŗd�E��Y��D	�j̗n�c���RV���k{
ف��j���,��N
*$��ߛ�̄RK��<��ꊲ�%'��YgC�̖���^-�{-m�P\��dP��x�����_J�p�G����z�!��/��7�WQ���\�?3![��tL�x��c��[�xҳI6�F��$��Y? NΉ�1S��ɵ��ѫ��JR������+1'g�u�Bb�䶈���=[w�4[T&0�!d�:��� ib�ޛ�_�-. ���H�'e��#�\�¦<]Z1��Yr��&63���>>����^���6�=��w�5���0vT>J@�(,�Y_8��(R?���,���o+�IA8tk���kw>���Rhh�N���2U�fr��;&K2�t�S�ɗ�6pG�!L״(,Q!���Y�:�(V���z-� �R���|^H�N���s�E�I�qP[@b�w ��CV�H�d�M���u��6>�"�-G�JT�,q Θ=F/�Ђ��+��Ka�]?&�d��1WKti�X�O�ʏq������/56R�_r��u���G�\Dot�3���f<��5��Ϭ��<cY�X�����1��}J�jF���S��FL��5�i�j��;\�����4昲�T	���0�5k9�<QM�lF�eǀT���)�諃C���L�dֻ6!�����q�����v��]ds��\��=w�%!߁Cz�4T`-~n�����ɝn��.
�a|�3-.�w�����i��������aD�!��o�"V���E� j8~6��F���Q"�I98p�mw�ZT�{��@�	A�"L�-\�?r���B����!��dP|��{ʓS%�9�kn2���.�Y$=�G��s9��+~�;G�����6��z��q�Mi��Tz�ԅ{n�5j�A�N�X�&1�����d]0�:DD���z	��5��%dm��g� X/�,���[~��v
I��w�;m�\O.��Xa=ܩ�y4�d|1-�t��D�@_q�{m�s���Ђ ����]�����w5�~n$%�4wY�h�N֛3S��A� >�yey)�$���-����C���ܶ��@ ծ���_����dp(�5��J��.�bke�		��F�N��^���B!�Q~�Ự{FW�!�'����?�'?s����jF�_���ھ�R9�h�>�A�A ��$��SA�����*$u�a�8J�]��n��ՙ�S�v�З.�}�D�d������i ��Eg������r;鰴�qi
������'0B���C�t�՞����H�0�(����rRwQ�� ��W1Y$Lz̡�޲U/���V	��B��>/�����LQ=]�[�j1���7�pF�FG�g�H3*@�T�+��Z<Z(�� ���x�"�*��Nb�),��F0<�C��oə�⺬��Ѯ�~(��}�c�`��
]ܔ�l���7al��F���{N_��9�^��s��5�}uc=ڕ-^g�ƿJ��/>�^Z���4s~�&��x�n_}`Qͻ`*w=l����+a��+�3muz�w�qI[x��
y�a>l]��d���ʸ�M���k����LhI�F�Zq$cp?�;@+�>��^I$�Хă����pnEI�nL� s��e������Й*�SJ��'���������蔷�%F �_/��<�L�`Fp)��@>�#ݸvj�k�J����%��Ϙ6F#ٛ����S򫃰�xz�o����M���2Ǭh����m�N �-} ��lTJ�P�*�����3) N��R:Ҭ��ѨA�l��n��`Ν�w�>"VP���)�����N0����8�i���Yi����i��︋},X)���{�t�䩲'�޿�0$���{�d����b~e�C���&�X�C�\й�����F�r�S�C��B����%z�]a��6P�E}��2R��S��\{B��m|���Kh�o����i���f�8.*�aԳP���ń�WG����#j�ѝpJ���Qu  �abY^�~$Z�gWh_X]D]��r�3�_�ỹ����^�K�݁��dܙ4?Ad#�Ƅ��G�gs�n��(�#X�!�����u�Yo�G���O&2O�5�N�����-���Ԅ�"1Έ#֘)Fا'$��>�CI�+9�Z�Ò(;2�q)9�N������c�礵:GT�1cWJ��*ԧ�:�I��*?�zF6��噿q���Yz����:�����2��>J:jk�F�sd�AnI+�{#EC�5�r�Zb ����y�ź����qJ�e1�Q<nHzCM�����.m&�n/G�Î�8-|��!Ĺ���:�c�-?�L�V��R��V��T��.F�}BƋ9��h�W�����9��D=���ε��S0��N5�l��x���{�����'���q��r��Z��R��������w��j�=��9�y�X��V<��sr����a�)���xg��!��f O����D��y�@r�t\�������V�[�uׄ��5�_K�t����C�bTծ $�;���j����	���!i��Q(>=������Ū�#O�n"��F�U���^ʔ�+K�Ν'^tpa�q,�yˌ�+�\�J����󋜽	�� ��ui�+!�L�(��f>��@pH]濹���\!갅�^�^�Y����Ex_/�NF[�{�ʩ�*vݠv�p�AW��@v�CTOl��&�>�1�0O�t�]�Q�tP��eR�;����P��Iȡ�ur-OlQ�#���Im�*�e�n񫏱f��T1h6��hT	q����ZQ���ĐHl�Ft1I�d ڑ0�[9����o���Q��>&�~��&�����yFF�p�e���aFW�-d�˚/����
�O$�ʕ�0��l#�鋪E:Ũ՛�l� ��ͶO���=���a�Ϫ��ʓ��y�#�u7Ԏa���� �j%f��B{�L �����o�E�nE�"��pyxY�76P#�������Z*5z�[�Deukٟ�jd� �X�Z�j�4E��^W�������kT��;���ki5�j���Ս�Pf���Y�UH
Ť�Eܜ�#{ސ��'�%�'��q�W0u��pk�M6�(B)�0&�qO=li� kT�u�O1�-�8��dQb���h��e8Q���������A�(˞�o]�e5?�����a���+;�7�ؤN��h ~M�,P{�h��sTP�m��M�[%�:xC�M.�+O�8��,�+� Xu��O##�ժ���4Ye�AБ�6v�1��q�|�;���ޙ�T�:�SaEhͯ��.��w���"�M��w��7����<�@e���,T�Nuc'�V��\=��m^ƽ��vOc���~��d�OL��l� �6c�݀�2�L;\�uD�g"�t�|��~�i6ҹ1�H�HRF���<��x2�C|o�ڠ�C�by6�����G&l�|ۤ��J Of�?P�Í�@���{<=��Y��'�0�_)Tb���ګYecZܘ����Vd@��(aq��a�oA�	"�h c�p��o�ǜݳ�,v�8�x]=���V�@���p@�����h����4ҏK!I�}@�%|%�����4�A�s��mET�9B���l����bp 7dU�``Y[XrT�K�MG]/�j�u�"&�Yj<<�N�!*�O�- ݷi%����ZkS:4�GW�9F�W� Pc˃m7X]��UZKGLq9NE�f��Ѣ���u���DD��<��x�4}��\�XV�93������/v�����=娈[*IvꂰTo�+�_й���"̸�Ǣ����e(��%�����H��Jf� �Z3��-濝\�d�"�Y���1b�fc���s��؊����'k�,W���|jw�o�<7i ]�ܬ�TဂE�Of�P���L`�MN����]��d��>�C��ui�Q��2����)�8���A,�c7�K��gK*�Z��|�e&����$�܄�:{�-`g�]
�S����2��Q�G�B�("p���	7v�?�]$�j)�G�l)f��`�jP&]���(@m�I0�q���I�pK�b�#��׬ە����eմ?�n����<ޔ���R3����[�$��wZNP��6$^$�ٙ>��t�P�1]_Aa�4���4_�����ML�k,���;"W��r=�
W�k���=��KΦ�D�� �p��A	g�[�B��MlDsş��9���#�UxY1r2!BD�K���lzð��ռڏE�N"IzA�7�Ή�h���%y���B^�kƴ��0��'���y�����k��ctr������`ق�pū�t�m����T`8WȊ'���#���뤷9�u��{,a0_&>�[&ܿ�g�Lcs��s^-DW�Ƽ�7 ǳ���iKB�'c.'*���+�IBj;�����]S��J�*�'�t���gHb:�e�����-��j����il�i�{I"cu�N�=��Y������?uzRC�z��N�1�b3���{x/��.w�M�-�s1(1'�e�@��xWD�;�ܗ�<��I6L�Q����u��2;k���eZ��Us�E��mMkZ��բ�̢

�����y�n�G��i�S;#���ڝ�䍪Q��n�|�U�*I�>��)*ڒ��婕f#̳Ms�3I�(�u9����6��f�l��d��7c����e�.d���:�~��C4l��bF8��9P\�X�����w�>�M��֣��\���W��dJg���"��e��@��qE�:h<�S@<��_=���3mů�������#5A�=w�Z�ZxK���~�����Xc�!�At6�Iu[�t2���`J�R���:��\֍kn�ϥ9���e���}J7�����:�䁞
�3�,'KcڭX�s�х|�z���p����S�fS>,��x[�0 �zD4N�Oм8�aqO;ى�l�۶��{�iv$_/����X/:�"hO�6��n�zSC̥�� )}�P�3�y�Жb���}��X[,CܜP���JVJq|N�������D�� 1����c�}Lj�}�D��g���6�ޕ)�v�|Z&���X�Ǐ��RM��[�h�f�Q�Wk���Im��iQ���)6\���so��W''8Gim̖w�(R���3)�r�-���� M<	�U6-#k�5,�r/�3^��*��\!�����|@I(g�A߱7G�_N˛�6�UpH�Tl*VV}���xT�����T�[�_=YK�,�Ԇ�L�ۇ�~�1}��UwhE�m�J8ƏÉAps_GϥPYF��&���1����L��g�@��H���(���8G�[�9lzӓ��7���0��{n�ߋY]E�]Q����74������h���!���5ɻ�B��[��p��R;!�j2ݶ-v_�Af���e�%���-�:�ָ8�?���8��Et��f��gͿQ���ؗ���{��q2D�R�8��Iѽ��T�s��#حJ�E_��Q�J�<��YN٤�H�2P�o!R!��{�>{
ڄ�����y2k�-�P������
.�/�D�Ӫ��m���綐H���d ��s4@c"ÿ�I����u����ԟ��׮�t�ē�@��\ �W3�Ӿ�s�(��5H�{�_
�JCG�,��㳰(	Nx*�R0�.�`>g4�� N��1��@��W���i]�¿�G��8��2|z]B�NOJ茰h'�:/��5�|^=�=�ߎ�T_�o���(��Y���=��H<�<��c�,a��Iǡ�ʹ��+x�A3�e4}�R,F����_��m�n���>�x�M*ي-�י�T�S�<X�#�2�龼W�Jmⲥ	P�Q�ԡ����4���D�Sa+e��3{'��9�D�6m@����o��,w|���B�r�Ӻ=�t}dcB(2CGȕ	*�1�sq�$Xሰ��LW���-<�:���l�^�mr��Cs�]�{����I��7{���9�D�wQ@rmND�N��ˣ�1�R���D@=?��&�8����!��y�k��K�k�]�^
"��:�K��S�f���	yA����}+	}��|��sz�G`m����|���p�X:ӹo�U��7��$Zѳ��Ѱ��%��}xZ��?�[����Y��&�Ju&Py��u|R/�f W�Jw���f��3�<��+ 9��]sxf'��j���p3�4G�\6E�Y�#��Ȩ��0B���yv�O�D�� a���]�B"%y|Q) -�3g���ԭ�;ǩ՛y��1����2rQ�0�N���V"�}��w��⒘$C�9ۼ�iu��-�HQW�}�]�+�Vӄ�3E��ÇY�j�'=E����P'r�6������Jj"[V���/��C4�0Ȕ*1�0҉q0o�����Ep ��_tϦJsӝaI��������C��?3(؀�*����i�[���k��Ҋ�eU<��&���&�@�`j݅�ual�u�S3��jWBk��?)@��M���A	.c0�E��V8���X��`���k���39W)����g���m�ս���Fo�_+�`���p}�y�>�|�#���}B��M�P�h����Ӿ��k0�q\6=@5i>A��H����|�wDų%�Tӗ>γ��㔒TiUY�[�d}�(Z�<�������G��uݺ&�ڇ���
t�%�|�a�}��>ɶ���f�]��\�l�#�YL��r3h9*|Iz��܍���h|M�U�Y�Yߝ��j��]�X!+I�s���.8�Q�P���g�[�X�A��.r�^6�)X*�Y�{���uy��U�Wd~&����rW_	vLVD06(�o�y�d����v9�4A_���34���g?�e��	�CGxY��Gk|���.�孀�=�ĉ]	��e��IFܤV;��u�Z*���e�	��qē�rΖV���򻇑�V��2��Z���C�\AVQ\�7�D���}�Z/�bb�>eθ&�����2�4u��B���媒�0�����%k���8V��������}~|m濠�H��<"ЏR��qV�ԡca�0»8'vO��]z��Β�Kأe���jh�d�s�{�n�*�s*�1��q�:)eE}>�q,<y`�^.4(L<5�V�����LޒH�P#�;0�Z­�O� R}�-�F�U-�^(=�@6Er���,��7���c�d��d��;_��g����ڙ֖ �v������GfD�����ù���iK3=w��46��Da?��E��@"\d��sAO�c�����'�HK��M��}f|��[��Q��[4l���F$ .�X'kԗ��<�.��]N�q�v뫙�O�6��J�&h�w��>�1�w��4�_��!�e�K�,�.��{�V�q�K�D2��LL�iE�q���l2����Bj��¡ޒΔ��֗����Ad��6��m�˂7�lt�tl�]E�s�ӗ�� ��>�ZRFY�!�.j�+}���Z�I�S���M��#L]>�P*�-�+Wm�t��8�/�+j%+"��)��,<�sc$��$����nyUu�9B��#T�L�U�����=i�0�9���]J�t�k��,k�	4v�a0zWb�}U�|0h�."H6�ھiL]*7n}>\�,xݐ_���}�ʩM�v�~�0���߁X�Ռ-<�ދ��ri�a��9
���a!��R�{����k*a^"��v�m9����/Q�vwaM� �����b�&/Us-��I�l��W��������_�B"jLS
�u~!��g�d�����|��4�'͗��,���|9o�V�y��њ�͑��N/e���Q�l#����Ul���(ȚU�w|�ň,.Q��9<x�x D�-�W8�.z��� h'�n@��7����hrB���؈���9TI�g�d1(LwlԨ��Ƈ.�Ww�%Й ^H�<��,S�����]@_��ayz����גܨ�Z����0�I{�`��2%D�Rj��$!�1��F�t��ݣ+|��CU��<��.2#�i�S�5��E�+��B�����!��K� �1!���V�!� ��w-�6�
 �vB�&	��ѧ��$ȳ�dѦG��MT-T����\���.���j�p��]B����D,��르���.h@�n8�/͕A�m�h���KZ2NJ�8ZȄ�$�_BT[�12�J �~@-|5�G�I	�<�k
���
);�N�� q��*ד� A~@��4����S}�1a�A_�/T� �͢��0��n���.�,3�j偢�W�� �q�K�*�	��S�ڕX�HI>��A��af+9v>R���m
%%���ξ��C�����K���|E��@Ԯ�!�d��0D��v�}�G��`��{��e��S��9<p3��IE�����a�ǘ��wQ�!J_^a���������hf-�S���W|���_�B��_� �\���.O�Ć�>p}�xZF:m��Ե�'́g1��	Iu)��?8p9��;��	�u�� �|hyӛ뫃�0�ژ���&���<���\g�g����4�a2i��Uv��Z�;Ƀke��j�gA�����Vj{�'����)D����OJ>���<㪛�=a���*X�Q���0���#'nP� Dv�� R)̇[�*�߂_��n_�
�)?��g�Ad~�*s&	)�&�i�0���ҧ���+g�-j��x�~O)�����OdM�w�y�:of�*kϏr-�:n�&�WZ�O+�@k��RCLoB}� T����X�3&�w�b�+�u�q\�z}�Bc�@�2@�}�(��ӂM�jǹ(4ݰ�lS�C�;�Ai��h�.�I�7`������4ԁժ��b�H�^;y��1��{��f��,�������KL������T�߲AF2��z&Yq�!����:uj���ON��D�}�y��=%��Bn����<O��Ɓ��M2����芆�L9 �-j_��l۹�/O���>{�k<T���sn��J�;{�x匀}�����.q�OB ��~��g-�iaQD�#�%���Q5�
E�C�gl:�л�	�=`k�J��q�ԁ�Z1�I�.�`��d:qa��o=�i���qc��S!��f݈��@(���&��C�lgX����O�M��he��ɍ�~�5D7��k/�ʴ��I��:`�{�S��؍�:y��Zs��0W�`/B��$�ko��&��1ff4f0G�&ʘ9��y8h��ߴ� q�B&�G� �m���.a[�H�sQh?�j!�Yg �����wQ�C�����M�8i.y��m�%k�9����.��+�T�%��V�K���ǵ��U��A�ٚ���ndW@�Kh�2v��Y,��9'�P��ml� �k�9�Ҁ����(������{,Y�AF�J��C��[�iH9��[�#�Q=j�~�8���Y��֔���2;��P�\�ՅG�4N����������� �	ȫF���ʾ�Gy�٠�/��j����yo��m���-��%>��&���`���RTځh�(���E0�
L��01ƱYx6̀.j�s�W�F��"�8Mjv��nN�'�r����{i�.ԣ8t��7�Q4�8�1p�،1?����G�ɭ��J솯{g�*�z`T���6V���&w����?�u��GP���qbS�XU��}��Ȫ��=[�r���b�uA#�J�^����EB�pK��4��_hZHh�t��M��$�^��{"L�>l�S�yo��+����x�l�3������7�<G�����RȜ��[0/ �'𙩅 M�z��~T�L��R�H�U떊��Mn-[�3<:��z��b�T���[�][B�����/5�z��[��9IQ\��4��կ?{�׾�����}���}����[�z_�E��;W\@}���ض�x�<�vt��nB��%�J���Ȓۋ�H:�W�d��Y����?�F�[0��.�U���s�ǟ9'����R+��n6�"΁�h��o�-t�*�)����ҽY�90v�5�:�">m�`Xt�ڂ�[��	�$�����w�rL�<%��e��kT:hש��I۟�Ⱥ�q�tlv�%���u�i���L�Tх�=` 24�S�9�wKb,��):���%G+�
L��ɞ���Ƕ���K��Z�3���f��+(������[��b���Y)/3j�X.ak��#ڮ���>ڞ�K-�}�"���|; ��~���Ԁ��F���o�z�*Ki1����#y	�n*���\R�:e7�z[|�z�Ӥ!?��\j�ֻ�g���Ӏ������lڳ��4e�B���ѝ���'B�m�W����-��i�7�o������"q��%"��T�s��w�݀����B��|��Jy����uL20��Sjx�מqw}��T*���w`D�BN�$�N:�2^&N� �)�6H���Wƣ2F+����gT��)F��̴�F�6���i�. 6?���X?�㦰A+�&�b(����`�����ؐeQV�� QM��d�������P�a�v��?�┱ҩZ���`A`���
�\�{wY/��73���m�/v��YX
)l���nmj���ǖP�/8j��^j��/z�]ѓ�ጼE��xia���(�����GHS$�_�/oڰ|�`��0y���L����&�ҁ4�^���6�z��g��?��98�I1
&l8(qq�sfr�W7��<&~��}����ESK��#VY�W1�1_��b��h�X���x��j+?c�>�,�%lv�ɱ�/��!qvnW67���ھ��5�6�N�V��*���Ǯ6�^^��#L���D���PI[+���&��p�W�̠�XR�j�NEi���c
����w\ś�?y�}�70��O+W��0����j¦���L�p���|1/����^#mO�rG0���7 ���1+|�K�-Շ�?0Dy��:���'�ط����p�2?r��ʗ����G�����}�GR�)C��t���������'av����z�_i�,c��8U�{�W��o�t3�>ލn�Ђu���{�y��%&�A�;���6������:��"�8Ѻ�,Q����b랩�2�*�6P{��*<V9́G�7�9r�яK��D�"��qvAt'o������������+��-jn����ٖ3�����@����^~���CI�jlʨ�����[���[�x��n��*����8a����]�y]mϋUO=)Œ+D�T^�	jf��V�Wx��]"b��^�EE�țM{~�ڍs�=�u,'��yF��� J :�(�m_�΢?�p4�W���j-�R�^��F�`��2#��9/�OlՄ���nJhKe�����-��c��[������5ޞ��eAO�H���3&yA)߃̫n��/�l�~��J�
����fs�Zv �;��m
Q9�ME�:U��Q��,����.}��=:(
>$ow���b�&+-Èn����D#Ø���N���_=B|)�8:�+��Wִ��C�J�*#M^��8=zC�M�&GW�?W���	6ǐ�����uv�HZ�Qմ��܌�[���g��^A3��3����RkHFX�1�X�@���T�����lc���OKy"
*�+6h�M|����}�MOY?C,l�'��fr�7P��Nиj�ݍʒ.~8r�(`��d+9��U8���h-�_�E�ȃ	�����uϣzo/����>�ߚ�K{���Nk±�x��4@&�e�9jZbH�����lV�*f�nl@�0k;j7�nG�T��
�u֩观����)�Y@�F��:*a������
�V��� �iT���3-��qg��ދ�z�|S>T��$dƂ���D�än��'?$��#\�wgE�Tw��g���V�t�F�k���!ōZ�ګ��GY7\���ŀg����R����6M�©.zAĩ��1/Fg�\��!��v�X�[��O{��$&=�ɍ���<��c�\���N�b�	6�.�X~+r�!
��G��uj/bV3��
�����8xC胲~����H��9o�@� >�Q��eb�<�j�,��9���U�m�Kuޢ�&��,&"W��O 9,]+݌�:��HL����~L3�bb�ܙa��2QLb.�Er��K�`�B��vy��)�/�9��#�b0�/��j�p<�N{
@���?����N�#���ͳZ����Uw�7N�.�~�"�~���H�z���, p�nn�_ �3/<��lz�ϲ.��ac�e�F���G�l�e������v�?e��ѿ�K$�Z��u�D��'lW�A,G����0���	�d��n)�ݓѻ'�n�Iq��Y�"�o��$�Q^�J[����8�㉸v.������Y�K	�pK~;�w ��Ǖ��)��Կb�#&dR�7�~��a�w�_�|(�O��<����_*�u��&��Gi����]O�L��n�G6��6<jS�w�Ƿ�����'�W+�Qr�I�ˇ�KM]o���F�M̷���q|���p�L!B��o5� �����Le��L���[mo��K��8/F�i럽/�P��c����0�(ew�v? =�0��Q�w�3يݚ�nm�쪕�\e���M_�x�Ģ���e'kS}�����{I��n�7+��J;��b������9��}ж	sF#L1�sN�a��	�|Ȧ��Ԗ�@��v��%l�CFɌ���ɦǔt	�q��)���{� ��7/ �^���Bs�e��*��};v]�1':�0@�i�7�J�g; ��WBhTo�$����2	��^]I@亁�K݃�f��ƾ4ӥA�.��r��D��M1z й��|<T2	"?ӧ*�~��T@���1���*��Pv��-ab}�{��}��!'o�vNF��J��Θ3b�EU_rX
���/`ag��5o	����g�G؇}y?�i@/���*?��܀:e�㜾��\�r��iD���Zu����H7����e����T|����Z����{��`�@��v�#�Y�@�]j�[,dt;mu.��ih��*��*C��x��ς������e�<�C�-�t�l�Ȅ�L��s�4�g�K:|���#��e��Iz�#�.\`5�B54}'u�+>�ϝ�>Ts��%��_NWtQ�={��vH�F�F�%���@��LƋ���+� ����} ��R���$ �2;�7��ϕ���D���&�P�q/�,Dq�D,��A�B��I��c5�Kn �4��$���,EUr6�W?ߤ�J��H�[��Rkҍ���J��%�D��X�����E�n
H/�u��u�����Ke^��Rꇬ	ߜ����m+aɰ_~Bxp��퐒C���!f�!�^x�St���u���	�I�&+�X&�o��y�o�����<�j�l��Q�ºn�L�N�V�b1�֍�6K K���f�|x�`�ה��f�L<0b]ۻ4������T���
82)MP����	���O��]���s��k�Eg��( `�N�턿�U_a�֟�K�l���Ώ���ݞ1��
���}�)t�l5�X���28������t�bJ��tQ�F����r��c��>���8D�^!��/�Q�b�����ƈ�4T�%�U�]a:6�^�Qķ/�6,כO�e��(I濨��R�⨂��F�cGW'�S�PY��:r��o��eM/�su� ���1T~\�ƹ����u<�qqm%�9�P@U]�,�=\;jݑ^�����#M��Ki�A���B�z���5�����$�Gx9��~�"��u�P���hHE�~KTl�>���ʚ�~�=	���6E 0��6�<Ϥ^�m�I�}��� �t��BK����vi��+z+��c�*�&� (��ޭ��1���+Wy7������ݎ���I"`c?���F����ٽ�>��C�
�#�p�!�N�7C�:�5�m��6.�F���L�&q�������	:�g�X��iH#��F!�j
�uy$g��u5�Ei�%]�Twf���m�=���&A�3�*aN�O����cH�L��׉h�鳉��PWKx�d�a��%N� �?R��/҂^w��;�,{4ً�,��D�ɏ�R��x%��\���]�K��'��BgDۡ�9�%�js>Z������/!���'���s�Nr=Ø����W��M/��0��5��ԣ,)J�{υDy��	�y������_c�D�n\8������̅�m����,7Ȣ_���"gD�'�v��Ȣ���5�����?E�3�/{U"�w��<����8~���׋AO��iG"p/��f�U��#�P��@��`�4��z�}Cj";�\Ll�~��1�QTw�,�Aa�܁�`�<Ǭ�R��8K�"n^7�w�+�v���Ǧ4�R-��m���ѥ�V�8���ӣ�7@���bT�s��y�[*�[Ȓ�E @
rm�!�8/���9*p�ћ%�"��dn�e��j�jY�Y�V���>�j*WH�����u]��w��}�����m���k�Pg��<Z���ē�H�+@T T�"��a'abTjSu�\9�T
��xbu�H�m����é��V�� 
�gM����x}�U"�]�7b����)ƌ�]�·�� �������W���-���Iя3=0�"2T�kA���]����%g��:�8�Њ���d&]e@a^�d�a����f���-RI,L��n
��}	-#ɾ2��W��^
J��)����ځߦ�� x�[\i�1a��Ѓ� ��%�NU�� ���uu�tC �rzRff2���z��'��� �랄���Xs|��=g��켫rov�="O@A�����/�oxp�6�Ų�n�4�����w;���A��&l��Sg nߓ��w�(�裇�FQ7 Kx�b��$�]������K���]9�%��!b�C�\x=cU�#g�<�#�ϗ�(aZ�²��ݕ?�1��ӎQ��z��,��{0��o6+�����F�!�Gg�* 3������)�XS�^b�c�O ۟F���k����U�[(T����(��]�\p6ZY��
�g�&�R⫕*.�]�����Qr�{9�4e׿�"�=e��V������t����dG�F��x#���!�J���1�Hu�+�?���P֮rcx+��iȘt��'���g���7��Mf�./� q�!H�kvț�{pQ���On�V���&p?��I�$~�m4��Gz�Y�%�UY$��@C��M�{h�����I!� "��P���Q�XjI�����9��������q�N
A���o��B�[�h �/`1Z�"BB������u�)��|�V O�O~t� �'�'a	gR�i�t�=A]%����ks�_ۄv�*�����X܏x@:\� �h9�F���,az�[._P��T+�2v8g��B���� )Cxb��IKz�>|��3 Y��<(3�&	$����fCΣ��@���/e��MM����d�;���@�U�ŵ�.���8�����CQC�8�Y@:���d�������*��V�gΰ9"��JyI����B�)��*��R~��n.���%�g��wZ����[2:.��hH.)���
�'��@'�<�fZT���̪Ze���y\[�|��;Ban��_�#EA���wq�r�hbAbiRvѵK�u�����bZ�j<���jL�,[�a����i< mP����.Tb�,!j�~G`]�ta����VC>屫[ϯE�Z�
�e����m��͞�7K���|�6�R�y���/$��d;c�S��Ϣ�`QP�dߠ��4�����~���J��K9�N����
�!g*>��p �>*�Z��5�����Gr�j�(���#������/.I?��ik��`_Qo��nxm4��-Y��4��^߳�(��l�8>�2?`1$� ���\�����Ԏz9�B	M#���a]~����;�T'n�����3w��;�� ?L�HJ~��aUn�b�f��	�����^1 � s�\�Q�b�k}�z�p5 ċbc�^���}_�8aH�&� �M����?��tQ*�~�_ �Z����T�s��쎰�$Z7�|K%��B�1��O��u�aQ���nF�� K�bΜ����!��,:��P����G�:�4�o������@y�jĴ5�ߑ=ҒS���_�<�L��/��0�Ϛ� ,��JO�3��~���~T�9�$7M�aM�.)��K�@�1�ö�ӈ{���t��Ԛ:��N��,�1;�IT�����1�"��J�̞,��kb��G�Ͳ}�~;��P������R���7rϻ�w<�r$��:���Cm����L���h&P֊8H�4*"�l(.��t��7��*�wɢL�aK��BR*G�z�U+\#��VJ��J��-5E\Q�߲O� Y-��&尻[�ԓ��ly����:��V�=�%p��4T��3Gu/��\y1jX��?�oY:�B����s�K��p�z��X-����"Sq��t���H��jz�@	U#H�cr �\fն�Ͽ��ϼY=���r�3�;��Y��7�D��CkB�(�I2Įe;�B�$��ǲ�P������.�b)�H�m��Hy>�\�1 �9Ue��[F����m"��8Y'�iT��ZpGli�5D��T��"!�!�5P̊��	@$qb'�|&MOrW�%���)�~I�\�P���g�Y8$��?�t.��{�~�Ś�0�ujV�����O{�R��e��<G8�W���K9vٵ����O������ pճ?0k�J����"��>����ϱW$M������Jr��#q�=�lI���2�u-,`�p�[,O,�)�|S��ˠ?TjI�育� ��Z���BT�O�m���&�f^w	~#F�"��5ρ�ݬ�2D�����zx4��-�&�<0w��ߨ��e_"y[�lg-�'2��)��V��?��/ڲm���^ �,�;���Dco��@�X!l��r*ڵ�l5Y���	���R��vA]�"�-�o�蛳�(����P�&y���w	N�"�ˑq̳�}H��h����
z���� �V�CFE�i�u���Xod�������j��N��*[�Lo���1�ݿXZ$i�r�:��F�����q��XK}zE���!*%�d��+o�4!���`�мxd]���}�so�lֿ]b-fR�<[GP�In���G[@�NP��u��"6_c���N?�]��E����㸩��� ib]�>laqZc��?�US�`<�� d-��#������3�m�A�:�7%ʥ�_*�._[��I09�U�38b �/+�I/1@l���o���	���=q��	w��5�Cȧ�~�����r���2y���u{�b�f�[��V�^t�׾f��?���Uc-8��l`V���1bs����k�ԁ@|:T�#Z*E (��w<O�P2-T�)W������ic�����N���R xu�
F�G+�亽��$�<��W�:B�݊����hV,-I�(�af����U��0C�����JY����^��)�PYIEDyjY.����Jd&%���L�gjqaug*����������m�tb��f��<E�7s���f�.� ���L������N�#�w&p��	7�"�ɻ9�������<���	��F޺�\�J�bv���w#�7k-m���~��[�xW��'Ǘ&���l�p����������>7�ml1V)���$܌pT</�oe�P���ժ�ט�#)�>�|�@�5͍���ˁ�e�5lhYH�8Ӧ���>'��,%��a� �ل~���-���wA�����@���V��u���Z�@W���'�,�E\Чu�)2y�<�M_«�? �yǗ$�H��bnW����`(o��h�ӯ�d0l*U����u���`�����8e�ɋ�<5cQ�֛$t��PCk@˪�e���"`NJk���@�1!�!pr΁�)y����ۘ������˖���X�8fx뻼�߯�H��%��m^A�P�k�)�FB�7{z~i�Oް�{,M뜰qg;g���I8�y�� \�������x���r��Ƿ���b��/����˝Y��a�\5�N"ً�m�,*�G4�R�Т��
m  G���/e�������q�5+�g�H���buʨ�I��ud�6���CT�|����Hb�c���YR���R�62Bf�������;���������a%���'�Ы��E�qV܋-C�W���_�Rr�`Q� ��6�H�dj�~�Xȵq��
l�.Rܲf��Xԅ&v����nd�4\�`�e2V�~�J~�`A���_�i.�r�[^+�e �o`�������a\��i�M%E��D���
&����8��{���t)�CjkE�I�)�'FD�Y,�!�����5y/�M�
�	)%�׿&l��F^�׳�E��r���sjt��3~�`��[������c�ZgX~��ٯu�ŽG
/w2R�� ��w����끱�D��@Tbj�"��2����� )�']���،f���Jbh_)���� SK�������D|�A�n&(�Ɋ���H_>�ģ��֖&��g.�ooD���{9���`@���	D�bW�؈ۢΐ�Yl��P���p�[��RB��$���T������$Ʋ�O�Q�$���r�i�*Xb���=t�dPt�9�[0_r��1�Un�CO]���n��<H�f
�!'7�5���Y_G�i�=-+��܏L����q[����7_H�����2S:[���L?͖?ǩR�ݎM�������zؠ�]q'�q��<�����~�9A�{����X�Of��<� �v�L;�p��ca*�#��Ӌ�h�_�����#ec�+@j�w ��6�C���m����\�ݝ*�Sd�_H6�&�۱�p�p����W���L���G;�R\Y��-��C��W.�-�b X��{=�%� G��7 7����t�lR�l���P*~�?o�ތ���:1���~��K���]���5��g2Ts��0*3_$O62V�mR,8z��(J��p?e��1|s��N��4��Ð5L�
4韆=����/�[�m6_�L�^���h��7#��JJj����[;�ZE4v"`$��|��i��m��\�����O����\`e\kzV��lt6��W��Iq{Fg��)B��[��f��V`	r��/`t�"���T���b���ro�Oӹ#!%�7r(�ߔ����@|΀�9�*���y�(�W���v�ٝp��r8re|�,�%^��Yt�������JVm�;�L�U��7��C�|D��i�Y~SݜSd9�.� v��ǽ�I��%��������<vk��P]�=QAz�b߃�-c[I�����:�۽��C~��/w��+TLv�T7#A��l��r��E����7���j'��\q�rs��ؙ3a5* �A_��F�澛r,���S@��3�3/����pL��$��oAP84��:������g?�s2���A]�'����K��U}y	LVO��3�iLB#\�����ڎ-�BC�'�j��ܜ�×�Ԕs��Gۺ����[���@��׼��[`ײ\��V�Kζ����2�9�Z%y�����4gyTɛ��*�=|:�9v��<������=J����-TĎ����4KJ0)����2e�W�w;|5�_o�=zu�D�-�&��6��z�7��>`f�$$�yؖ#o������J��"��i��Rҩ����<���I���K��Wâ��5�r��ֈ`8KYD��Lr>:"t�*H����I�������wkӂ����4�4��M8����SnԺ�!���T?���*:�Q1���%Y���)+/c����i�:��*�{��:��s�7��H��j45�!�ɇ���I�� 5I2���8����OB�0Kn�1�\�8�*�i�����2���'&�mCY�����@oac
/�֏PY��Q���x>��R�D	q;��܋!�tO�Q�����q�O������%z
���
	�7[���#���8��$��c҅�c��S4�^5�8��:���j���#}��<%�쪬3�z�p������f*&��A�Fp%��q�5|˹'y���7<�������L�<.<PR�H�\	ϭ�Q'dM�B���Y�g�Ln�i<��@ߍ�av�L2&9���l�|�Ű����K9�Ѧ�ӏ��<h�L�Q�5�܏DK\�����8픭R^v�vÛ������u�G�*���ք��Z.��`�5@ËXR�~B�n�ݬX��N=P����hJ��v��+:�)+p'"^d���1:�6̈�`�!q�ISu���'3�'�Ux��ig��a����U0ayltLF�Z��Y�{�Hؗ�BhͲVa�[J׌��I�M2u���_;�4�Xy��Zgp�^��exb��"�(�Vƻ�|�R����DQ�;��1��6�'ф�夾�mv��p�Z�}-O�t��Or⸨��������\��W�
�h�J8ġ���2�ޏzJ��򽺎aeu�:�JR\�l°Wc˔��2��L�!�Ul���j�^��}��~֣	Q���(q������@%��}��h�ӛ�(A�.a~*C'�yH���f��+z���3!�V���ㅇ6J�Cq_��gvXNJ���Q�,��x��Լp))��8�2�J���Z�ϴ��2QV�W*X���B��X�����7�0�,�}�-��x�j�Z^�d`)Z;�g����LP����?��o'@�"�B���ѥ��u�{������z׈��$�C���7_�.��Q\`
� F��>�NK��N^�r��tb��%�֑Wa�^�tCŭ3ueo|̉?�(�y��R�ZD������e3����c$���Y��]��'_ì!Z�~ %P���?�ޑ������J��FL����n��-�
S�l
 ,���ORo(� o��n��֮&�#�	��_�|cb�Վ�$G���X�)���7Gbi.��X.��%����$�w�p��{ cü�;�"���M�3��Q�{���$��oL4A}�:�~��;/A�_S���_�/;��@������n�@�;���Г�9Mu��l����r�]�7
e~_I���I�m�l�u��$L�K�i�J&j�AHSbzb��i���p@�o	�wIEX�fQQb��Y�f�
���_��	_�#D��;ť�Ĕ��n��c<��Q/8\��E� ]������~�':Hhl�!.F\KK3��jC��y�U����0�o�!h�x��I S��m"��v�%�u��$��)�iF�|ڄ5P~�|�E�eB���Ha�nI�\�f�6��p=Q
*WbJ?�+`��{�R��)���C��$0�N����/{�j[�v���S���ؕ2�v�`��׹`�A��6�BѸ�ИK񄗴��!X���$��߲�;p�����跮ĦS�=��?�M⽤���R�M�/�S�*�⳥�����l�pt����ϠDx�t3Bpe,$��'�*�}���=��sbk�8r�}��@o�m �����9��T�/-��D\z:3�mHQ���'Ye��������۹�7`�t�\cu����y,�ܩ��R{�d���.ޏ�?2��͏�n�F�w1fb��uw,{ ǣ�
��({~=��8j���V�;��/��(l��������p$k�Pg�sy���ZEy�:�0lH!f�;�e��!j]��k�w��:�G�A0I-�c/��>\K���)��x	>��d�-����u{����� ?;	r��N�.X[u൓N Z�\�W�ʡ�J�3U��w�Co��
&�ң���Џ{L��؛��oP��}�h4��^_b#C3����(��'����χ�Ĺ��3U�㿘y3R����	~�s�\�#0�ŭ?=Vk���1�坜���Ic�ꝷ�=u�^.D�l"����ËfՈ���
G�0��OD�h�����k�G��D�Mx�OZc��	hL��ٶ�P�Zv��).��H湥	�&��w�����Ы5��p�|�_Y�_���Nې�S.�ئ;��}���/&�vu��`����fV7�M�ހ=TU#*�1k��P�\�z�O����¿#+��4�&b�{�́�5?�%����[��1k-��7��S�{���J����YC�U�"A��\6��YQȗ]ۅ|���	�Ywy�U>����>Ҥ�'�0l7gx��J�f�Z���`S��8�Q���(��}��O\Ҟ�/
	�UFf�=U`a&(�	�$F,U�Т����<UD���y|��˻�����-n�4�d4���0���_a���� ��5��vu����j�vy��@h��%�PNh�qK��h�[�'F�y�p(���	}"A��f�Ɣ�9�(����$P���w�A��c�U�X+����JL��7(��F?o�*�7�\��Zjxi��if&�,_e@Yѷc��MK�N4�A��
)��!0���<��}�}�=F?:C8B����q�Q�����+C������w?��hc$<Y��C�����ڻE�hȰ"Eⳅ�h�/�C��	Z��m(Q����,���Iö�%�P��������|�J���?�7����e�Z#>���;�h��;FV��QF���X��E:���X��G�F|C�4&�M}�:S�0��f�v�n@��{�ߥ�>2vt<3N�\���9,��o6,$�ዧ���s�V������a�D<}��"쪪�@FD��������a��CYrr"R�� 8�Q(#�am��������"��9�sH|���9��m��|�����<Bj]��"]�p	�7~��~G����չH/_��,�3�f�A� �>{�h
�֦9"��2�\0�2��9N�!�pʠ�Dq�h��MM(?���o,���r�;W��0�S�?�!2Nj��y�s��*lʑ.f�6t�����r��>�?��s��a�N����p�9�RJ1��sX�:�o��3�a��ώ�䛜�}�J2��9�	�8�ۅ"b11�u%V�H�S�Q�~ΎO�/,d�5U<
�	��c>�U�I,T�еS店�t�d��VE� �~iE��y�������P%
�JuwV�X)d����c�o%T���F������|�'�y`�� 1n���?2��[��O���r��D�V���7kV&jvJ��%?gd�-.�2��*���p?S;a�������D~e�u.r�g, k��m�7J�e�)�?�8����I��1�A��@r`Tϧ�)����S��֎��f@v��D8�t�.����^	���I 1��1�P��"��,no�d4`ll���6y����f��oy�֯ω8C��@p�5�M��s�Wu��Ǜ���3^�����A���Q���(���'È]�Q�YS׈�\�]MG�,A�o��U��=�"�!] �Ŗ�ւ�`%|t���6:i"�	��	�z�T���i'������ăo�s���j���yT[eC3�H�q�t�u�KbD��]�Jo+5.��
���%�Wv��֑���ޡ{m��p0&��>���\�z���H�Wf~�1�a���A8��=GW6�eZ=�ݶ���SO��5���l�����`��h����Ji)vy��6$MTK�|�zG���u�"��-S����$�t3��0�l� ��'��ʡ» ^ĽSU �w�'��5��<m��hԞm?#q��[��r�ʮO�ߤ��xn����"[�^�*������a+���v�3����cm��,�Nb����u��j%
�`�����%U�{�pÌ���KvU$*u:	�X%n�^�a����}�6��?ĵ�������M�� �2�G&Y/%��I%%X�_>ἠ�cp}~�K7b#�$Qj#������Կ�c�]�!e��o��z�z����SF���!��s�>8�{	�G�cr8S�j9��+� ��*��6X/�3|�ʚB�tF�)�bDъ��n�����F��r���B�����Tq#'f��Bڌ?O4��CF͝�~���H��޿�pm�-��k����H+�/y�Q�eeES����6�h,��m��s��L��HR*D�<�ɐ����q��|���i��]�,B֭�¨�����kc��f��U�ke�D8�j�Y������ϋ�����7K�������T������z�E	���)	|%v��o���,�IC�����"<C*\�nQ;=�kH��_C`�*�:!��A,���:��Xp�S{�&i�5S2��o�B��Y&�3=�R��`:#�����,�>9���������p1f��+��D�{���9M��#�����@|$r9�΂���.��oM`?�@�p�^�<�ڕNG�:�t������hَ��d
���&k*�=��q����o�w�r�rr��4I\�^u��J�B9��FT��J	�+�"X,�J��mX>������)t?����s W-�x'ɰ��7l�t�f�u�#l_�@���~�1p3��0̡U�M��*7�'��mu�沐!�P#�^�t�v���5_y��{I�����~�A�AU��MK���o��+��d�F#t=�����T��hG7o�o��I���TOS�}+B ~-�X�6%!��0�ĸT+�E�m�������A'j�.�����*0.��bcd�3D�y�a��9̙혆C��7S��d�
x.��M��V��g�������	L^�	�!2E{��0`�<y�YC�����紩���Qִ�.��Y�� ([�^t�׊�{T�C��d��C��H"K;��;�N:�/ ���-%͹l�,��QǬdg��r�
�4kw�<H�+K���^n~��z5�~0��WS��"{w-�j����T��X�����`N��i�9��xw�ha�d��u�ǀ��>n-Z������`�M�Zˣ2UhTȼnQ�0W�6�?%QGKF����6�W݃��NO����`o����"C�� �W;֨з�QǛN�q7�-m��L]�Gxs�w�z\���A�4�Y��)͠�!�JA=
+�9[;�s2(�|�C���Y:���4ׁ�/p�ο��vE��:m>�0r��o���ݗ�O��@��؄��<c?ٴ�nLz�uEYW暟Ɉ�7�t�C�U�醓�V�b*�o����#_@���Gf�� ��[�S>��t��5�����Êcx7,j�����9�VL�e�2rdG�ƚ�D�syL�Z���2�K0tD�u�����f�-D\�at�M�S�̭�(f[c�L�QK�e�@�����?��sI�e�_��K�ꃘ��TI�ᩒ2����^B�b�S����`}��?����G$����^{�.��P��� 6Xi�S�˸�.�\�t�� ��=?����_�T�Yk���8��t��:F��d�Z_�I�L%P2se^D�Fr�5E���T�"qW<zV4M�_)�4�������x���
ǽ�q>�|�"ɻ�(,߭�5�vwg@:@*r�@	�ս<�N7��֞�J��Z��	cS��/�q9�6iw����CC��*��6�[},�csq#_��<�a��x�)Ԏf�a�/�AM�YȐ����ߥ�
��Z�9^5������b}�a��
T�b	�̡�Dw�p���q��dt��C[�%//�J���#��4w�TG�Pp�v8�v��HC����9e��{{��6Z�	��険b��V�E��;��Rs��+ގ�wg�li4��{ �u���;�
s��=�*t�6��TW�)ɿ-!�stՑ�"O�u������OR�\����)3��]ŷI[3�.�"��h/g]��[�X�R���5�.��EZ�����Kz��ss�ʡ<Q�<aK��#��+<���ߪn������cn�+��q���m�UORI����>ۀ��d*�Mj�q:G�'��P!�^a��|!�!)�Cl��n)�,Y��:�����E�`���Eq鲬#����\߯P�w� �NB��"��4��V
�}��5�k����~�$��Ƭ�-����M�%��U��^�Ҷ�8��"P�Xi�`Qe��JV���v�ė���֟����yD�:6Elou����� S������-f��T�N�!Al4�#���}���5��]|�wN`f���fq�B�h��6.�N�~��B`]�3�M��Y;�`r~a$�,�2�Y&%�dc��TH�e���&|�����5�XA��7���3w}���a2�],;�����~JbN�O�k��������c����w�֎u�$?FÕ���C�ؖ�-�4˨�i��*�ă�џ��K����͈���f����Q����֔qH ���K�j�ڽ�~�,{�9��t=��q ��)��s��n�o�x$a�O V��!ƪ�kX��^_P�x�1�1B��P)1�yO�C�%�={1۟��!�nO�&��pB*���EW�%T���aD>t�x&Iq�i5d � �r]i�� �M�ag���讽{�7/�.�ȣ�m +�Ǉ�H��{f#bR�:��D����W�+&�`�xm�V �E�ێ+���jt���������q���3�4!O?;�k]��Q��?���	�f^�1=��||�.�OE'I������L��(�R+�qOW�`����i�}9��\�`��ަ;_\�����f�� ӓ6Pok:A�a8�)����3��ϑ�QnS-+�.:%,]�q�\h��q�F�2�p�sK:{�΍���*�v��U~7DƁ����z0>�)Yg�+6��w��B��p��,���SЃ<���Qf��(а���]F9�]F���F��&'���ױI �O-�Ӵ�B4O�%�",9��م�m�& 7O
��b�Z��۶Ùw)�rnaw�����+���Cq=�J��n�d���y����>��`s\�[7T��+A=��{o4��U����\�e�%uiA�v���(Z��*����V�us�	]v8i�nIV�\��@?�I�9��>��tf�E���c$%e����@��cTpq��kFr���D#���P������+`���Ѭ�MyrD0�d�XO7�"jJ�ܶ~b���հ�CŃu��p�,�l�V_��M�8�.&Y�Z#�	t6"O�� <�����P�K��<_�)���!���b�N�]I4�K"P1ݤtdš�l˅Ӫ�]���5
�,�S�Z�W��;|�:L�'���?�N��Y�?g���_���9��$�O���J���r��8?4��#�WRqE�ݢ�x���Ą5y�O=L�b�/���o&�����s��|�+�o3�5U��9,�8��"�&R$�����<���GM-��ڳ��cL�F�GW��x�s^.�s�g>/������?���b?�g�L�)t�Kx׹��	:b�7�]����[-}��i_��i����VDy���Z����ĺ���b��l��³�g�5a���k����{x��1�o�(��G�5��S4�
?�U�$+UE>aa�4b�LAl|�T��W��i��ayp��A Uz��_2��A�krH��w�9��E3Wk���QxI(�gilI�T�K�"�x�"4`�X��m?�ů���B�3��i�x��I�>�<����
`S~�
Ba{�R|)��+K��U�YF��7� �z/���;���&�y��9D�uR�0������iӼ�}ǧN��Wpp
@Bg%�\&	�� �B��U]`�ZoT��m�����qm7=�8�/�)����W�P&z���X���s�D�����E&�^���%��a��ߓ"�����>�-�M�+#i_Ȧ
#�����Q��)41c	^�3䛗ĨCM6�Z}��S�涞�5��̑+�%��]CY��{b�(�%a��ґ`�oh�ިhO���ւGk�ވ[���oe���Y�Д���r+,K��ɪ�����NFM��H"��x�t��k���Q	�\1b��:o�ڹB�*΁�$��l<�;L8J�z^$���$���S	,x��܈ �5�槬|� �cW�ѕ�Z�͖[V��3�"��<��q�� ��Ԃ́���G�5�,���5��6X#l8�~��.��4���n@(�Tͭ�t�	v`]�SF߳q�	|�ߒa]�\�
w5!�H����{	�^0"O�� <M���YA^�jQ��3r���V9����i�s�3�ۢ�F\�4��uQ���Kޢ������F���¦�%J����q�����,|�t�i又��$��Y���
�W��0��=V�^G��2�6����d� y2�[!A9F�x-����u���aa9K�����b�,.�"C��j�߁�0� �'�+�1ϊ�J2ɱ�=�l�R��2��ѭtQxg�8!��F,�d�̞cˊ`)H����R%l-��A?S�*�Ka%�gt��6d����ɉGT��5�Z{��;�`�(�_F.ُ�u����?z��l�^���ktuXP;��� �X?'C����ա�&X;�Q&��񕁯�#H�S]��oH��c��K�����q�$mC��Ց+3��c����h���G����ǇbH��AU�����F�EI�L����#	�xnhC�z��7��2D�^�e�1t�l`z���+�Z�0G��;�h�0�B�QE���l+�v��یvI�*�t@�h��Գ/���l�G�;;R���^R*�L��S����*]���{G"8�� ���Fl�W�h�_A�R�.H���&v|�}-Ɔ�aPH�^ȸ�,âe[%U+s�w{���a�"���[W�m��������e�Cz��J��*NV����z,�IszE�*4̓�nJnz����Ί�F�#�5MGUe��])Ѹ���MUBu/7Ƽ��Ő�4Z;�~}��'_W*Ȗ@�-�(����
�Q�o���,��7�OY��Ǎ��"#'c_w�W����M��P�75^ ����Y+jh �i�AG��y�6p�еd�� �O<^3��$����4+������^��e��DZ��xL��|X߭������(�Gb�}8$� |l����x7��Nu� ��0����������<x��E�������A��G`�����BFѼ��8���<i��z,���`��JZq�I����.e�w��d(�����9OB��ވCʭ���\��2�(�����x3Qo-��T�	�׆����~V#���;�A:�X� �삫q�B3��W!
tJ�@#�1M�8�-�jj�EQhV�gAVw2~t!K��I w�������UP� �Z;`tK�<wǻ���.��\�Ƅj%lU�S���+t~Y��uH�tI�E����� �{�����T;`�(e_颢��\Z/���K��r���ț�0�Ξʫ)�3i��G���Q�m�9�C�)���IW�<2���(e�{&���!'�/M��'}�-��~ۻF��C�$��o�a�}�U-R���pc��^)���p@��c�mG�4!�d���]\���ĵ�RsXX��^}�����@Q���Đ�ZɌ�W�I�W�ƽf\ G�-7ۏ*��U����c2p�{'/��@�Ю�y�0�P�C���ڜ�f��S��rso��-݀]��e 7��o�� ��wv+�i�mגy�bN*[�SО����ZM5U��%�W�i�[�Ǘ~���Y����� �,<GJ+y�;�k�G�4֟�|�?	����=m�k@@���ƍC/���Bf�]�H���&${ �zm��sV��ݍ�����3(�i�xξ&�0ך<K�XT����Ϻ޼;o��y�v�f��o�r���%��ca���:��in��G_X.�&��k�G
��rqhhGod�YUl��0[)�:G}`)��4�4C����ȶm0oe�x�Ǹ��Xi��
�n$Vz0����+C�u~�9@A6AB-F�&}&�.Av�,�3�So��+��aVA��f�{�W:�����̏�-!��tHĺ��D�,T�LA����X&h��'ia��}�b�)�3iPة ��U�G�o��5e �t^���KP�_D,i��DLLN>磦�d�.nU:�!L A�͚���+�.�6�E�c&$u�*u��j�4�V�DtN#K?jP]n�"O!�Ĝb]�DcKE��vӇ0_�a��N?Ⱥک��/@�+�+�Ч�w6�f�z^����A�S�X	����kI�g�=��q���nSuF �D�����tOG�b~6�wV
ԉO߷��gγy V�V�a0BD� 8M�L+S���I�Y��Ť�� �飈��#'��������֛ V��`�5ϛ<:t�Ճ�����T_5(dĕ������[V�]��W�#�As�z�]�4�J�UY�YV��.���<v��#b����WK�drk���k�̊Ի�s0'*�����X�W���:	�J#S���C�����@�MN��ЗB��,�������''�|�K=��m3�\�l�pi�G?Kו�Cl���<Y����0���y��N,K䔖0[p�KY��g�7��޾�Ej;Q�è�� vت\7:��%���N��a�2�*��7��m�DF�(l�x�'��Tr��u�0,(a�4��;��5���ą���zI�v-Kk덂E	�����d���QM�O�4���zE������[_�;�P�?@��q�_ω`��y�����&(���Q&�{�W̒�e�t�O��ܗ# R�5�2ۛ<X�� [l�s�hlҡ�yE��u@���U��4�V��~62OU�C��1��S��3��iQ���g��G#}�C�7&����!} ���q(�U��]���T�� Z�|����$�����n��H��jIAS�.��_`_�$&Q�ڊ��,����Jw=~s<� &hM�_��"s����%|ܫŸ��մJ{��3v��fY|X�-_��(��p��ݢYr{�yb!��$ֵ���ʲ�2�U��Ua��(���U�09�U�`�}���4���{��KIXvoH`�؅f!����cg��������綏ʇ򾒈�e�L)s_���K�
�2Ś,�3�	Ʈ��&uC=�O��Kg�Q}0��=�Q1�d}�L��*��ԧT��m��|�M��$jikݢ�h��$�+h�Q��ux�|�oe�����hQ�E���f��T20���#m�I�~�����J��dh��ǹ��e4ߒ$�M�/1����s�d�G��X����o�A��}(��a_-!�rE}�$�$���Ċ��	���{Gs<��\����k?V�CY�Lt�T��2ٗ	[Α��]z.����O/��EĘ��Y{��)�o�4��'�`��̉�hK�R�ڏ��{Xzw�k�\X�J���.��#�][��|��~>�$�k�4M��p#���Ǐ������fmZ��?�A3$�g���=�;�&�a��(�4�H�C��8d�&m�MGE!W�ǰ�UQ���
ւ�����4�Q���i9_;e�>KEW��	6L����N���A6g|�|�9A;?���ؔoo�)��)�&ه��δ�v��h�7IEL@��� ��MS�#{1<fl���H�<�a���!k�Q"�8fѾ6�w�����4�����絽)�ۿ�����Yk�=R��Jl�H:?ס�7�E���q z>�t�55F�$��b�+t&��&��m{�c0䗔��ꋟ�=K�� ����F��~-��(7��o%���S�&y��ә�q9���b�>�KB���z�v��d�E剒�T/�_\�hX��"ލ�S�W���
թ�D�*O�=ֱ��Jf�IG�Qs��#{��H��͋�0��h:�*m�ODR27j9P����k����"k�&@
^ĳ?�-��L��xMEe��U�xK/AUBAZHށ�٩�i.��pM-V�����E�S�h�ժ%
�/'6-D��`C�� l�]Ϥ�pC�:q��O�[��@���uJF���hT��/�3�^s��o�C�ƻ��0m�˥�w��!;O חF�l
�Hk�mt%�y�����Ho���E�w������ND�_\f�H*�\���� ��j8� �����a/|�SV�: ���倦��d���y�6WZGA��:D��1�ԻS%�5�?"X��78�aO�w2s'��h��	�*Nה�Ef�w����`����!���ńza�|M��?#�_�@�fq���jt]�W%��N�4�K��r�k�Ŀ�k�0��<�o���E�j���)�����		T�b|N����m@�c��9�R�k��0��-��f����6C�j�D�He�c/�0ZF�:M�R&3sXk��"���7'A�g�Hz� >���dO��[��y��Z-��L*���p��L?������L���+��s�\�`;AM�3ZIQ�Z�t��5G�VTje$���Om�ƃ?ލ�D�F�zԑ����Y�Ɲu4��N�c���_R���kq�&G�@CG&}���Y}X%�	-���[��\�k�R�Tȳ���*D��̍�+`�h�c�m�� l�F�(k�}�v���7� ��5nmG��p�DF���rZ��Q�|=N�׵ڥ��z�[ˢQ �rh�}�5���i�����G�>C�?ό�N�K���6@I�f�i��ƃX|
gPE�8{��I�'�����^�>o���D�X�V*H�{0����T'��3P\�p���|���\(��X� +�z@+|n�2ᴬ잻V��u�9�GFyW��M� lt�18�L�\���1�T>��5l����w�]S����*�{bvG:��@$q�2�.*z�CjX��E/���11$@����j�x���],��ʥMo7!���j�Y���uy�U���T%�[�n�y���`0��}���9����m5��-5���q%j�9�h���X���+NԔ�PѤ�]<���%0]o�CZ���Q���[A΃���Vޘ�2I	"5W&���q"P{�<�a�ͨ�9��EL9w|��Iݤf���?�\�sdʓI��5M���r�9�o��:<�� |� ��"�����⬺՛�n\�l#mF���5#p��AAN6�+�_��; p�f�Xe���������-F�_��vỊ���X����{�Ua��j���b��u�M���73��j�5�MC�� ���LJ��9K[��6��:�������8n����ȗ'F���r����&��۾2�>��\�K Ll�Ƀ5��������0R�a���*�����g�|{����ZJ��{�Ө�:�-����X·H�K�mY�p]�W�i�ӊt,�(F���I�� �˨ͽY�gT���^B�uuhJ�*k��]���hS�e��I����䅕�H����p�����c���借H�_�p�����yZʹ��,��U4a�8uReW:�j��Zx{�:�Y��*sd 3]�E�n6.i�*��I`����FԖ`��X��.Z��M��&L�j�o��?|�`+��U���R#3���/Ή7|d�<�!`�T�3p�4�l�FQO23���:=SL<�
�_�.����+��ՑH�E�'�: ��\�7�+>�zVa܍��2��yg����f��v}�b"�h�@-�O�\F��بۺt~����Yg�T�'.�+�ł�]�(j�Ǽ�u9F�2�npY.DZv����պl9Ԋ� j���׿��O]lR�x<�J!�Ҧ�»�n�jG��Tp���$�q���X��i��r����o����HP���i�o�x.�5�t�,����r;�Vq�<O��T_?�}<0�7��f��u<4����*�͞f'�6�_�}�������Wbs�;�/\ʀ�\�ߓ4"��c�&�@ir4��3#�˯��Zj�V� \5ڝ�D*_�Ϛ�.�N.� K�`��ã�|�3��!CG��ZH@�ڕ�w8g��.�I�2��_�˶TΈl��^4
TNsض��g��}٥��s�P�F>��#��dF�CĔ���ӓ:_-cȢy��f10���|"bB��W��R��>aXM�@��|��M����G�*�A.,�&3��p�|C;e��i�,8\���Gya����`�]Gd��惂�E۞1�n���P��4Eo����1l���P!��D�ox��,&�Q*�9�q��*閅M ����A7�i�Ɩ7����^��^g,9ܓ�N�$+���QD0�d��Mܜ�^n����"+C��m1R��kf����_�N��ERE�����NrA��������_�f�e�2F�:�I�_��*;��tioo��+��c�Od㇛@�%���c� �z��~I� ��󓋩B��,I�f�uRj��9��6�gp�գ��|6(�i�a��؅V��vc�~�$e�>��s��Sy�#"�ez�r&�b�Y_5�<koL��5Ӌ=.�^Ph�2���+ٽ�A�M��^�Oe�.��-�Ѽ1�`�W#d���(쌡�dܫz�`�>3bL���|�S��z�a.�ߟ��fNL��C�P����&��~�a��
�������e�ɂP�5����l��ªD*v�k�8Bй�t���<["9X���[�+�h��� U.��W�K���e�Xg'!�6�1k�Xgln+������D������ ��۫��B\>��k���P�f*�-m:;��'�:�~Y���h)��&d��S�i0�I��}:F�uc��f�� ��I+r��)�a���A4=�q�������R�k1�nԾ|ro�g2.�"�oך�:�T�$S�A+�f�O_~7�Wvx���1~������#r���~�~0ӹ�(�b3�����;�q��޻����P�_���X� ��i_�>��l� -��e���*�V��i��o�R�~]�cV���`��	�hU��(���q)Ω�򈪎�²l�X,��#��zVزWPd̛����lr��>H~[��)4�&a�,��D�"����DNL"�r�o�/N�G��$�Ȉss	GK~�C�����zj����q�GZ��g.�j���'A�	ɚ=A�=�7���!�'m1�]9����V�e��*ϡ	|`�<��k�E�FGkT(��If�4&��g��.��(��b3��*��`vg��!�,�ZJ�kp� R�:��Qx�J�k��R��Q�:x1�D�:�a^����D)��&���o�0�U$�N��X��ʦ�ůݢԝ�%}��^���02|k�rO�T]y6�� �Ν��A�dF���� �B�ka�$\h��=,�W}�bL�G��������	��?ax�)F��v@��gW���<�o�TKv�/���v�� �5�[^�W;\֬�����|	ZC�?�#���"g�hi��.y�ks���=������N^� X���Lh~W,5|���3��3��r�0����nT���1���^YU6��rH||F�$�婕���Vū�(��m�UW�7�?��L���a��@��W�y��9�I|��g�#��nB�-�u�D�[GD�{Z�;��Ң�3�XX5��|�fPx'��-����ɳ�M�1٤��!�sE�i~3$��S>*LW\s?W�)]H''��bs���&��y�!z���U�p�J�.�~B�bp��l>W�4۾pG&��V�]�pa�8�J��.�/:F9J�|2^�ԩ�[8/����䤒���:�E�+���"�EZ�RG�L�|�&�Ğ�DXZ�:ŭ6d���Ί��(��|þ0�&!�?́�P�i��3�Rc`�r��-���0�; O�	aK��|J�
�[��G��F�Ƕls,Π�Q�C1xQ�~�{����f5f��R�2����<�\W�`��c)W�?�� ���б��c Tm/u�lr*��d��ؿ�G~!ĞD����a
&��Zx�������B)9`�
�u�Q�*>�+��;�}��u�Y�MThG��r�0�=}���$�%/dD̕�
�~�D>
b����X9��bR M�Oǈ5���އ��~}'��߭�y
�ďw��
&r�N��R<��UQH11���p%�彩��nѡ,i��9�˦�@���� `Ha�a16��W���fh���L�`n�8r�`%v��U�f�`2��9=� 9�elg]��ս�j�!�t�9���K�b~��K�1��MnF��4�O��#�z1�憭�h!�YWj#�
�Q4_w�����\ʹ�+����Q|�X�I�|�3�XޕG�����AZ�T<I�^ّ��:雓ϯ�������x��|�P�G��P�up-��l�u&����e}
�'�eO�ct�k�AH:x-.�*�>�a�JL2�����@��|��Ċ�'��ZO)�*gTW�W�7GPb��{s��Y��ð���;f{X�!h2Ԧ?���:E �Yt��]��ă3�a"z_&�j#:�g��@��p�c��PgM�?0��X�Q-x��@�l�a�:���������P���ݸh�B�&��(vF�_��u��J���<�Qa��4�v!�t��#T�h�������k�LƖ4��=��g�e��'�O�ѫ�N��j`���a웺���#�V�
5��|��?uH���h润��lZ������� d�o�oFRH �k���%Sv9���!%���=y��aso��T��D�҂�Ǯu�q.�R@�A���be;yTȧ������-|k(=-�.�Ŋc�v�/hy˶�*��D�
���$�Q�'����+ I���ɞcB��`X�D|��Vu���?�^�i��&O  �A»��3�n�!��:�Y{�8�c����+��:�$5�����5^�,C"���;�x]���+Zq���D��"8%5�Z�b�b�q��U���\�)�tpIe�nG�2���nJԓ��7>X'd/����\�������`A	XϡY����3���'v,�,���a �>��Y��9�(����Жn��y7B�kGn�
_z��;?M�3���� ұ�/�@R����(~�8YZ��6^nW�EZ~ݡ�֋+�czS�] ��3cVS
G�GQV����:j�ws���k�˞��2�
�k?h��H�&��-�Di�h�bt�� HnסI|��q�
z��~�+� ��z���֎��Op�b� �^&:���@]e�hNxe�����~82��@!��F�����RD\�y�����ˍ.��������k�-�Y<ƾ��=�:Ԩ�F��ԬIBI�4�������t�	N�)~7��c���]Tb���+B��L���I,6d�ED�q
�v��.��S�L�J�m��2l�����Z������]�\R�5�<��棶A�bM�2M�67�E\�;�t~v@�ϖ�����^���cq)F�-'�B����_5�3�{�]r٤wf���neޥ�[EB�U�k�� ���]w=S���2�����V�����<��p�4��J����o�K��0Z,H����ѧ�N�z��p�C�j,�(~?���|�)I���?u�"�����������<3�'�w3�1��o�[��'6)`3���\�AM������1��T��&�`�.L3�q�x��8�
W��͂ω]}9�C�,ݛ9d�ė%�@��\��~c�6��(�5a�;R�����W\��n���CQAg4f`�(�0>O&���w�-�9[T�)�O9�$�ԇw�?��`u1���0����DO����ĽL{��!S���w���H�D2}
�ݓ�YX6hn;��׾?'�����2�������ӽA��������;E���D{�[���S�o��<��@�0��U���~������(&8sy;KդG=�.p:qv�����P_�<�e�(�dA`�; -_�+�/�xM|�����!��;he��>(�Fvd�l�d�<��2����D��!���_�"cj�pz60�N�^C��kʾH���;���5@o��Q�����_��?ޢ $>�K�"�g��{3�ӭ�KJGX�^]�א~���_	l�6杻��`��[pe�)W�$[�v$	Ƕ$�'��c~`㳿M�y��?�/(�~�t��y��c�4#���C�v&���N7x
U����Qf ��B�����"	v�n�*��o�-U�.0�)���ٚH~6�f�F16@΁	f@N����\7)��oc�>b.����zf 8����gl��)���/���oiv�S_~~Pf�M�+�b�kĲې&�U�~~6S"���R>�g%�� ��<6s�n�o:,�uOm��,hˑ������ Yh�� V��Rƶ���ET���$jR����L8|tוR8��G)_P�J�+X��A�C�]�?���l-y���^����:wΌ��د�������:#Ey��ך��ľ��ao����}����>Gev����A�a&�$�g�c���uX�]���w��$!�e��p��:?R��W?\��}�>R��ɞ�PHޫ��E?I�i��;�5�6����t��o�)ֶ�7{$���{ٷ(�I���|	Z���	*+�,�Wr��hXլ]�X@<c�ީѳ���$2�&.r�[�� ъd'2.��X*!&�U%1.a�����T�>�i;��l�a����fL��H���ob8��7WǏZ��s3_cԪ0�{�o�F�^��!���-���:B�˪��=,m��oшM�6���Nhwm�v�(����w=��%���R���R����4t��Xi�R�#� �\��2k��:�N�Ӗ��z���=+��y�k`����N�~&^@o ��6�5���:r�K58'��' �<E$�eP)0�r�TB��g�Cp{H/��u6�:��ִ�3�����]��%��4?�̖���Ӧy��u&c�Q�4-U����/���4�)>����f�4<W�8	��I�(��^��M��"�h��,��8��@ǿF'��H��mX�5�ż�z�b@7	RHYeUM��\xn�,^mK��1�_�ahU��`� �N�P�V�b&��)SOC�f-4�|/(��#�I�g��&����Hom��Ѳq��
R���d �
�s0����>ͪ���8*�kKtx�A�9�RXwh�����总(�xp�/�ʬ��J|�Se���+c�j]�x4"��%v��R�vN�aZ����_9h�fuhx�r��D\��E�^G����,�rK��j���7h9�*������)1ϊ�Gqh�^
�b�@cq��y)������Gj��Y�5��=($ӹ��=z�?'::VW�q���9�����H9�˽�������B¸�+��l&#���7�2�	�#�tX���ӓX��iݜ�ī �+�J���"�)���z�ݕX�SXA��7��|.ګ.�:<�ʠ�{/K��^�?��D�1�W�e^o���..hO|F�IL�2p�ϴ=,#O)��r���T��U�w�B��[�/����A��桯�/G�:r���7:_��6��(��\U���/j�Am��隙���	��ۮt%R�.A5qF�8�1텹���@?Iv9��\U�ᆤB��'�OK�J��]R��]/�8]Ы�u7���.[�:lg�Vp���3�����:b"5�Æc��W{�8��f�E��2A{� ��;G�)(Ŝ����"��h.�W�8�T�] �{�(z��3�;��<�D��_>ˣ�"�X00�M�qˈ���$����a�: �#S0C��s>�����*���.��j!U�y�zs�[[�!,���Z��Ms~���Y�dgy�B�M�=<g�x�z����hV-l2J��c���~� �>.�ǔ��������_�&x� �?��>�	�W.R�-!OD�=x��]�=���&{sk+F��ZC� ��Kn�7\�G5���O\$՜PMd�Z��-%����s�a�t7y�g�{�m�o�
�GC�)zO xq�b5��LŦOgX�X�W0"�*}q�[Q�fp���َӛ8�F�����[��'ƪ/�)ɪU>N�f�+]8�fr��ng�c��vvB�p��5O���nh�XY	��V�A�A
"���#&�"�U���������iވ����G�*&��پ�E���X]"i��Ym�?�s�hQ��o�w�{������O,��pĳ��%F�<E�v�*&~�܊#/�O�c�%˽_gpH��[�j����K�g��-�W簰��$yobߒ��I���h6��9�(���B�w�_0 �~�T��愒O��r�H��p ˤ��*q����M�P�g�:	��xfH����iw?�9HTE5��}�����E��Kl�`R��hUsS�#F�l��g_C�UV����L�*L0���fZ_N��B?����Ћ�o��)"�Cx��B�E�<�A������`�ɥAP8�4��������j�pHg�����ya�C�TYq������.<���P���7y�"]��������\��z"$[��z]�b1�x��h�{�ӵV���r؍�6���AAT��!�y�ַ����';EN�R�K7y\����Y�^ ����K�㱩�v+W��E^�}��~���΄��tb���7�Y(/���ir1�5
��gh�!"�q�d`�&��_��:3��I���+�ɮYn��5��Wx�sƐ`�*�_ _�2WEm/k�'P�U6����	1��������a���5�Ȩ�w���1{��|���A ��dOt8��U`��5SK�gŴd���%>�+nOBBmp�����j�f��S�#��� p�(�rRG�_�A�2�	�.�_n��}g=������C��S�Z	�_4<��B���m*W����#J�^��\��-~c#�u�@ڊ�jo|�~�^{��/���y^Yv�@��0�����!� y7��D^w��_{��]�6��:���2��p��.F�MX#ge�p�p<8��˾w�� ��_�a����4s�%Qb�(';��q�%���"v3?�ʵ���6�:��ˣ*� J�l"�e��H.����U*��l��\��%e4��@1Z#��[���y��o1Nn2�o�r8�KH;�A.7�|����$#�� ~o$�9i��jQTq�������A��i#A�hJ;�)9�^:���|�BҌ���ԁ�Mp�2�CZFWs��-ه��ii7� �c�C%���p�|أg�Ɗ�GP����w���S��Aw�;�	X�Ta
�I%�]�e�a����c{�p�R�q.���z��:��('b��d��G���̣uiǴv��ʷ��vg�8�a&�Vm�qNmO������B��Ζ��;Y�*G�Sjb���$뺵�,��??2^�����-m}(�w$�2��#�b�v��4������)o��B@R��'�3k
A;4ۖ
���u���۹��$���-�T�|������ sF�Rv�grz��y�0����62��J�
���-�`�����_�\�j6��H5�]���d��||�&��M �5=��j����~��G��%Ocd)�n�7W���p�����޳������g�f�.�óH*O�� 5��<;B2 _��x�4N�<|�1}�,��(�[��̫�[�y�s-B�oρ%}R�ŵ}d�1�o���5N��XfW�a�$��A�V��`�M��R�e��S���i��c>%K�����`:0us�P�;2_�'��.t��O��t_o�!EW�J�K5��f�t@4���$ʄ��z��k����})�HJ>'Nw��OTs�����&$��9 �0�:}�j��j��ӫ2��H�F] ��	zt�p��q�uc���,D�� ���)�-췕öt�D8��^ˉ���y�݁Y�/E�
8��谊>ޢS~��|fk�k*q�R���O�����$�Y���-L(�6[�_��՘	�G7�g���6�.��.@��%ef��!��-����]�ܖ���y)y׀%_�o�k��8����Iik���ٜ�u>F<�:s�H��R��I��y��/���f@�Yh��GZ8��[�cm�%ݟd�Μ���2��k�gl�X��6���]���U�	KF�z��F��n�y�אI7�h<�9�xܢ�Θ|�����^j?��$�~Z{��F��4���$�^
�3�^M�^|,)
�!MH�A1��i�i�v�2��`)���nu,�H�9��U���������M�(�ץ��!�Z��wi|�]�;q;EXfBR��e�����l���ۖte���}3ZY�4����
��g�_����_����z��<��j�M����9��q�*��0�ev���j&:>F����N����pw,~�QM �i�2�l���(��ȭ���vA���ֹSj)[ui��&S��}R7��͠l���X��T� �����L�wH�-��ᨤرq�0� �o|,\�.�0x� �{�:?�5�
�:aKOZ$E���	q�m�e�ohn�{!�O6�Xtj, P��>����h�yP)�1z��c�4��8?�K�R|f��(w���`��n��f���� �m~e*��2٘h�g��=#"�hH�j1{z�6���C�L-%����|nm?t���S/�% ��f�/��7�`���T�4W�1��;$ȧ-'t�,�t���_R^����0Q���O�Yn'xD/�k�/�B{�jM6�R�OK9̨U+L*���Ԩ�Z�m�Z`�C��D|�;Xf��7��P7"a��8����21n�00�
+��x�W�~�,�(��3h�i2c��m[ؔ�)����3Ru �1}1�?{�Y$��ʊոjuFoX20-޽X��=||}g�\]�Q�� ��~f�K�Rc�8# ��*0iV8���V��";�u����j麰1	�rW�*�Q1����cU���Sc�_#�K+AQtZu%_P�bO���@��=��鞕��D�[r�^���1>��QP�O����M4����wī\Ar�kA]�9|��Z�Bчp;�<pfR��3�HA�"ʍ!�fL��=�r�k7�% ӱ�l�PK��	]��چ��:$p$/m����."���1,4H�\*���63"MlB�v9���&����c�4R<&BSl��m�H��[	�U�Z_ҿ� �X������{r��9�*��,#�e���W��p�|P�=�f�<��w���f����6�"��2!b�x��Y	��&A#>d�x�s��)|h��1��2�k9�N�;¶�ч	g�!�G�U��#cD֭�6�F�YpL�;vk��"Y��;�&��FD����ͲDu�H��I��B�� ��������f���<���_�Gm��#w�k���~>=h�$���(ݧMR=9.6�\�9�+���,{��_��v�����k��39x6���qCp'2b	`'�|s�bm�S�.�ݽJ�C�ʴ?�&�h	N!��[ t�����9��S�ůx�����"�/)N%�b;������S얏~�����9�{�p��_m3�P�)��?`3�NE��pזc�?�ۭ�i>�`5<Y��=#l[χ�-���[�+w�=R�p���3���	�n�l��S�gLPb�3�c�����$�g}<)��R	Nk=t\�,��a��(���:C޶�( ΂��6��o)�pJD�1��{X�!aێ{4��
�)xGv�%�ŏ�<JW�Q��P.�4�T�w l�eG<N>_�;��y��%�M�;f��T����=���\��	r7�\��p�Fr�Y|�x�@q�4D�S�R�Q.���~uO��]�ᇄ�J	
"�`Y
��{���S0�戇ו�N2� �ш�5���8�W^�~P�z|ahFqŀ��h��ҍ7-���xw�,��ȿ����7����Zނ$MȆ�IU���-R�ىi2�i`=�u�B�����B���z��/�r! ���GoA��O=9�@��Q)h.���{�F]�?�t�2�qr��m\IflB��$r��4&��+��bR�F�@HySs��jw=�^����,"��� ������oO� AM�ebbB�鑞��*,�.���>rk*�����$M6;�?H����Y4dnme��-uY��O�k{2㡘��5c|�A53\J.�Bg�ӳ=@�NO��gP6KG����'8�."_�Z/u�ۆ��A.u������ǥİ��	$֨c�E2i$H�^A�B�0�@��)��;��#�Pa�g��kBqSl	�i<�<!
;bb��d;ʾq��H¶�!4Ξ��4��-�MJ���}l��-��f��r�/׋d`���5��U6�x�MeH��YX�
$�ۇ	c��g��bP��@�0�f��h	���sL|]5�류$-�Ҫ	��X��lRIN�^��š�6U%�˞�g���, �'�@�H�[ԨQei�	�b[�-~^m��9�Ϡnww�0���~�36���@��I��F���K�W�����3N0������F���S�6�sC�0�灾G�
�!-Oy�(&c}5"Wo_�]BFd<sAL�I(���KM~&n�"����a��/��eش�F��S�(�I������<��7�#�':�A���9I���C�P�p`�gl$�0XP�����K��%kQ��w���	6d
���T����&ℽ�b."SR��e����0�Snnp��Mtd�Wp%�;��z:L՗��x��]����(c��Ug��[�jd���B��46짏rP�n��I�._J� �g�I����b
z����yP�1~��@�6�_���!�z���!�jN4�;HPqY��F��m.�mq�����<YU4A��]�I����[,irYlSh��Hj����
��C����ܨ.}�9��6�E� ��k�j�E?H/3���#��c}���������q�b㫩�u	�35��vo^"���!�1����^_��0&�N�� B"����y�|���p0s�`y,�Q��`�KA��V�E���ʞ����B���_oc��ɫ���'(cc�l7�&jd��U蝷~ٻގ?9��̏���Z�Tȸ�H��q��"�eT�Y7��o`�1y�ʝ-�UN��x�V"�֎2#{�a����K�rUr�9�tZ�"]_V�va��Es@�����!��1P�t��
�����l��Xdr\����}��ƶ8q�8�/ȎC��?e�u�~�|�P*�5)-�h�v1�w���9t��'��:A.���1�\׷�p~���=��|��G[�ϫ��ƞ�1�T��D+(��[���gӂ�~#~rzl��+�|��Z�MS@:E1��-
F�R����1M����]_tA#\"'F�[�pcn(��7�\�]�����Ѧ6a� �dq�f4L�!B�F�H��u�,~�7#���y�E��@&�T�o���= |��E:԰[=�E���n4;@�����٥��8�q5Ӏ+ g���r��W�0�䬕-�+<@��zB�Z*���C-c����X7�<d�29���B�k�RZ|����'��K��
��EŤ4�a��K��=��ُ$~�����5�$�a.pȼd!K�4��0+X��s���fL�S��$BT��0�3��u�^.f���\�9�0Wc�ʓ�h�v�d�|d<�n,��j
sϬ<���wV,'U}�M��M)Zd��8s澹��w5�QC�X���!f-~��AAs���d�F�����3��u;�\�+��FA

`�J'�!e)��k�į���Ԑ"<��b_��W>�RI�緭2񸶒ڷ�"�|�`kEf���P���fV̬pN�o07��(1"n�<)��qӧ���%KNd;'�=�4��@p<rz�Y	����+I9&kf(�{`�5�1����#�i�#| ��!��E|�FT���7��:��P�b;+�i'�7)xտ:E�l�]&F�;\�)��I����	 0�^�ھ��\y�N{ELnH(Y�gJ�����eB��	DB�����jN�#�˳�㊯P�����ڪ��,n�b��8J���[=�ڼM�;,���3V|������1(��Txw��9G���054��Ϙ&=}�H�6���<6@�_0e�)C����*軇�(�f{�XM
�f#��d��kV��º�8r��i�n��z~P)=�=�<@�!G�D��}���n�-��^��i�kxj�i�#?������e�%��$������4'ى�Ur�-gFMx���xٴxF ���Ƕ�]��i������ ����չ��JH~�}�\�LND�C��M�FUa�����~E��:�\Ɵȳ�M���+$P�3�Aj����'+� ���#i"Ee�R�ͅ�a��(Ǯ�#�Zy,��j�9g!�+c9?�Nk�	�1��ޮ��5��������D�O��q"��<���9zp�I���О�<mꙘ|Y�U@d�m���"�~����n���W6Ά�p���d�u�H͛#I��E�i�e.i Űݘ���b�zo!�5Ld��n� ���Ѽ�ɀ��&䵳��)�JG�I�8�'Q��VSP��W�#�����T��s1J�:��z���ïOvjTr&Ԣ�Eۏ�}�ƺ<����E�g�?��\V�8��Fw�����VK�xK<�NS�#T��>�����;ݡN�Qx��X��Z�!Z
O�B��T��u�<c��u2/���1�/���8��`M.���Q�����=�[�G��2(�!���ߟrQ��:�%o�=�8c�~�Ón����H�t&l.b'�h��o�������]�Z��s�[�n�
�I~���Vdu�Փ䏓�&�A�;��+�̉I�^xR�͑z��������K�8r.���`0mu��x5<1;��;IY�^�ĩ�Ї�]�P6a�K�r�+IU�)h�J%i{�)��c�&���3�-�$"�R�P@T?�����$p���$+�)_�*9U�c�M�Y�sʸ:��I/|s���A,f�b�Z��*�5�Y��K$dh��eV:uY�{)ңq��e��A�И������6���$�|�?^"�ģJ?��y�k���р��Rn6�[��_T����a��`2�Sq�n�]�Y*.�Y�V��}��0�3�BH4�-���>�tm\�W6	�ʒZ�����>�g��c}�$|�\�K:��I��ֹ�G��O��F���܂�����v�/2��\�6���=&�%�@������82-�ͳ+zF�e}�� w�Z�$����W����)�M�D���OV���<�UD���^>��_����|�x2�kR���g�ن1����P�h�}����G�=�n@/���k�:�kI����潋d�c��K�iAa�0���
Q�����WC�����ѓ�O�o's��"AO��ExA�殻�R��e�P>E�3C~��E�^����5<��"�V�YΚ���-��\J�a�����<E<[п�[�#1�f0x�si������:AG��������.Lŧ�kN$h�}����H��Շ-�k�<p���d�6��6��/&�M��e�ј�b��!�k���'쒇�VN�T��[�!ނ)Z��@aӢq7c���5/3�B =�J����'�T�3\:�8K�����V��=(�\Έ�!��͏	�`G��!�B^���1F��87��J7�;Ҿw��%`�*�`Rǯ��m%��e&*��t�-�@	��v��b	�p�|���+0.,N9�q)b[Pm`sV��3���_��FGFm,�g���G�t�B�G{
1������m� W���E��|]�������(M�׽�?�b����6S���u��6����x���yk}w��2�i�yr����F���Q��e�(�A[��,(�>��'0�!02�h�?�{���-jc7��q�I[[�Gp��dv��h��F2���x2���J�V���Xt��|6��d8���i0h�ߪ��y�]"��p'�2�+<:� v�qj0S�3+���*���@�}��Qnh2�g+e��=(|P\�r���?D�!�]I��n�h��f`����U�Ѕ~z�Ŧv���Ԉ��>�_��c��B�2V��������'��Qm��>���f2�2|!���(�URAX�ϧDv>�^������9�1�A�G}������B(y��1�\B���bO ݐ΂���+�_��@�#���>����=���D��l����������Z�H!�� �����׉��\��j�Pv*��x뉻���mZ����5@CE[��o1�n�`�>�T�F����6�>�]���(0Y���;�oef%��aG�����S��{���ْ��P�C� ����f4m���ÞQo�c#+/J$.�?xϭ���>��Q��{#߃��[�ɡ^2a?�E7c��Q�֥���W��� ��X��&�opR��yynRH��b9
����Sǘ��d�i>Jq*C-e6\A��N��R��J��=�P����dC�GO�,-�;g_�_$
3p�G��Z��1���&M���<I0�<rB%�7͎6}����y�M�k��3v���V��ji�=	�t.���!wF(�л!���!L���$<w���?6lFo&��@:�L@jn��8�!o�@ā�gIW���yYΧd@����MYi�S�x���
��C��z&5}�_׌�+:�����cI ��5�2��l�(�v�
���[����Dcv]��یތE�fjե�Pø7�\v�X}K#�ư"Ǆ���pI���k��g�@�]k��4l�>���4��@�YC�ߧ0�n����]͠&���D*������!'��?�2�)����(��E��
u�������,r{46W���X\�[�B��y!]4')n�Sh Y������i�_�
��f��7�2c�ơ�m�K�_Ql#JOZ���߷�����W"��`�c-v�d*�jw�t�8h�/hv��ª����Q���K�U�R@J6v�͸�߇��?��WEޗ�.
ü��TY(�;1��?��������j,�ݸk-����\��2͌U�w�K*�같��p�0f����C�4/�r\J�񜱄c/�S�,�T�7�����Lh�i�A8����Zi�����5�:��'�Բ�wA��͚������JS"K��[�j�5����|��EwE�#�q�Q<�:��:�]��ӓ	G|n����u[�v��}7�]��C��#�{�`w�N�U�=V�{�o�ˊ�Vn��:/�Ԁ�}W����~N�ݏ��|��<��p�f�lb�)�a�,��ME>�4��y��-l�h<T�����q��3�|Lq��цdR�u��Lq��!"�CA�8ݓxD������;����tN .�������K����	�oz��"��#jwt�h���請03�F����cis�smO����؎�)bt�(MP���'��7J��,"HA����٩z� {�@�ts#�HO E�t�ޜ��O:��^<ূ�D�΂t4�n�OZ��0I�����g^�	N�v�@�Vx�i�2]���v��<�D��Q�\g��:�|�|�����{gPN�Ҹ�9�k�|WHR���St2Hj�����-��1z�E<��T:�ٙՁ�߹��M
���d�l��P���dk����F���y\�I��� �!�1��J��/�«dKB6<+��/h|^rC�]�O7�ʰ��eu��6ô�V��z@quK������*��2�1�Cۢ�$Ι�
�Ǆd�F�R�x���'�$��
2�~���%�WBm6>4���A����Y~�H���l`[&��	��.� ��̧�4n
����L�b?>_ �hh��'���#s��8�V��4r�F����v�aF���Y��.�K���> bx\��I��:���hþU��;��^�6@5�M��dwōY�v3�Y���#u���7) ��M�N}<����y��t,h��vN@n�"�А1�d�z�Sߴ݀A��<�oW������M��B��Wb���-�.url�!glS�p��[����!�ޠ�p��D0�	2$��mg�lKo*�=t�2a��K�,�lvBl+�k�桭f�WL>M%���ٺ�����m:2�=��KцlKsmB�֪��G�g�dP�&j6۪�j%���6z��E���S�������LW�h����q#�hi�i͔x�]�72	.���65L�!�%{=�������P���N#a����A���G�n��&�c��RYGJ]p�r�#)/�m���h%�s�ϔ�-1
O��٪y�V�0A�⌅��VXY��X�G��8qa)a�>�(��N�}�����'*�,��y��g�B�=h~�'�0��ŭ��aY���,h*��呉�<�oϠׂB|�"8�)�Ū��Śh��`�T:�3�/��`�3�zRu��CDIyh)+?�ĩ�p&
�{���Q�7�����ǡl�+�A^֥_%��Y(Z"E/LL����:�쟕�1��'N���9Uj���k�/�@��_�����[����=������Z��N�:h�A׻3t�o����U^����C�8g�k֘C�z)�ߡ(=�
V9�V"ɿ6=���v�ߍ�5v�Q�D��i]m���S���ߧ�2�:����Br3�Ac�pA���P�}*f�$q;8��k�PpH{�+�����������]���1�U	�~q��fp��0��҉<���B�n��?$0}݌���H�����n/���Iz���D�ɱ�����R�14��Ѣ�1'���	he�N��4X����bӃ��GU�C�=�V�w_\��b9��y{(h7o�������OB�)��q��m%
}�����-��1!	ʳ����-�o�����KD�^��,�ϵHR�,v��ܺ�Ϫ?�1j'���$H�,�|� �;�$?����F�.K~(*6�"��r_�4z.E��Xn����p3�����Uג�ҳ'���4X�M���'"�|z��i֝�ha��y�:����c-���7�E�4���������0I
xÄ���E�OX�}�qZ���l�ƴ��e�~
jm��%�xI�4Һ��W��F��G�%��~����� �3�f�@G���w����'��6��=�>Y�|0F���Q�V0��R�� K�H )E[�)�%>�ݘ��pl�GOb���j����	�۫K(?t�> �Ѯ�ڟw���F|�������ܑu��F�ؓ+q3�6
yO~���]
���Ƌ�@���h�Tb{DCт$#�E�&��loB�?��C�uTCHjĺKλ06�Y�������Pȣ+=�]V,��8�}�7+ҫ�"֜$��uR�����ӎ�᰺���sK�܁�g���@��D����D;U���T�G�����n���X�~�����4��R 'r�nlz&Eռ������]'of���e��7�	��Xa��٣ s��"~�><G��j4�}-�`�dU ?d���ɲ!uh�P?���T'��I�S&It�I�oρ�A`j����*�ox���#%V���Ѭ.z��;��;�r�� 0�}�6:�8V{�:�8�K�o, 9Ĝ��m��c�VJ�ug�}O����(t�U��!ŇI����4��K�s�c���v�_#�()Eb7}�_�pF. �v:�;�����)�3�?bR��"�X�]Zz���o|���
?�e���0(�
�b��L��$��Έ�,����h�M�k���=K�KƊ��5�=�:X�2�$%Fё�g4Ӥi�ugߛ~$b�g���R@47_�O/��R�V���T�<}t[|��(����_����	�l�m*�v�T_u�,������4��j���փ�VT��=T�H?9q����h��=j���[E7�3Y��Yl�6;��3$�V�#�@%P"fYmYf��sp��4�ʷn�<Z���3�i�Z�a79�B4�_j��tξ{�l9b�6�J�{6��hE��;��pO��Gu�.�̃�1���KjqY�����ᒭ��P=޲�tHJ����8	d]�$)ʟ�����{���87$�������"(���T�����F�\���u�t���=}�чɒ��t�Rk:��"2�/���}ͮI��@��� ��l�͇���o�P+��-����C?�U��� �5�9��P��ʋ� �CW�]xB=��Hi�g~�6+��K�ajw4_r��m� �Εp>�$2AXR�."^�55��1�)y9P!If�>���0��|z��j���Ӥ�A��^d gU:\Nb��v�!%��P�KW@^�̈́�YX�2V8�R'��6^��R0���WU�E���\+8�B�̒�[1�\y3�z��p��{����k��0��%�QzӜ��$W9���7�<��Pm_��T��Ҋu6q�"s��ܦ��x���ސ皷>�:�ɠ�]LywI%�!� �'�Y���K���K�,{F�6��!QJ;�~��*d��uP��`&G�f�6Aw�-����T�ޗCv�=���FG(�������ݯ���Jr|���7�	Qbm��
ݣ1b ��`��k����̓�\ہ����XY�9�\�c�i2E�0����l���ݽ��r�{B~{�G֯�Ą��c镒�9{H��9�g�u�&qI�>-����'�+o��}�|s��?�(`Y��z��:\h�v�H�|��!t���v�#���ph[q��_QL�*>b�:-�j� ���Z*2~�g�"��_1Y�<ntq~�4��ɡ8�/���m����>�THA����F0�@c�$Y�wg	4��l�݃(����{%�Iy�����3k�|�����/1y��m�?Vƭ��F}p|B��D�Z��Ⱦ���z~��Gϸ��vw�c6��6\J���(���BO���g��B� ��[m �@�ܞyB>!H���[@HV�dL�g����L���F4�nM� �])L_C���^��C;�22�m>]b�_�X��/��"\�j�z��3"p�B@ӝ�^e�a���"E-� l�#�-�a0�gT�Xf��\��2�RS��������"���I��>F�{-m�oWy)Kᅴ���6��@�����)_i��i�X$.)�n"B2Z�u���C���ႅЪw)MLTr|
ȡQ�Jm��u�S�'�@�NHF'���Hm����Kt�9pd�	>�[�?�S��GJѹ? ٞ�C��s��K{n�u�z���K֌Fq�
���S��m^qw:���-�Q9��L5��{?��Q�sn�����_K2uB�����tx�K�6�
�X�B/m�!�EN�!�)�7���U�[�`w�B�Ѫ@�/�%�v9V�>�:��{�������ir�Od+�t��e�u�55�a^��ǟ������_�t1d
Fc����:�?C`n�2	�ZS =8>�Rc~Z+m39��i� ��b��9��p���$=�ȓ��T�g��-Z|JW8">���Z�O�*�()���g���>�|�ҫ�nT�E_#��b¾�O[n:��n�RVko�[�`/ΊEV#a���+������V�$��fzys�L��-�A�ӯ�8a��HCkxx=#M���:�i�X1X��^4��F0��[_Nf���Yxz���vWeY�[�-�٧Qe�[�N�u<���^�̬%��R'��0��!�~���=L�����rm��q����s��iVk(�u�Ku�(�ZU��j9��ܢ�4�r��XjSdy꬈FG����O�ی�{r���ܽǬ���U6��*v���#��k��v�����@}ݕ��:�i�2h�t�bK�),ʤ��������~�u���(���Um5{V�E���r�̠�� (���0Z����έ�q��R�_B_��'�6kla6uT�r)e����vS�3���)n��D�5�8����@�hi�b=(���r�e$��?ʕe�� j�Z�P�ho�:rdC��:�C����D�nΑI�HV=H9;����Th�b���a��K}�I���<����m�
���tP"�7��g��aڏ'"m���^A�,3r�(� �`��������𺘆Ĺ���
���N��0΅�5�Wɜ�o@��A�Ks�[ʍԞ�0�+*�,�f�>u���w�0��MC���|���F�\��@XF~bC6�oD���w��a�{��O�PӒ`�%�H��5�Yʽ�����?Nq�PJ�{D�V��~,x\!�h*1eQ4[rI#�F�Z?�rɦ�OˁJi�� �b��~�!4��a��oݡPۄ��?��[h9�`)��E|2=�v.'�N��b�g%��*z��/a�*�+��u��Cs�m��O,jz�G8��d5:����`�=�p��F�E�:�<bp4	�F(�G0�TB�c��|����6���y]�ܞ� e��h+ H.��h? h�ua�@5Z��nnқ���X�'�j&��_>0Pk}�0� ���U ��V�K�(����v3��;�˻J��~l�a$����^���
r	�n/�B~��s8��$Cv�!�������`-��ۍ^}�J����q�٫S�j���0���Z�[Qt�9%84!����K���T�����?e�X��}]l��}��|�Hq���ƟMUT��C�s	Wz;�P����gE�g w�棽��������(Zw U�:�--LF<h�*�ԯ���{:ح�<�Hc����M7�:��3a�?RpA��/9���1V�`�3mn��"ȸ8���j@T��^��1{��M��J�bm�\�z��D�s�<�{G^s5Y�RC�ڻ�'J����1R��RDԃ�3o'�8ZVy]�G�D��C5��c�r)���U�D�`T%ܖ`Y�����Њ%%]6E�:����>��2�E�������G�#�K��Hh-/Q̦��r������A���*ϴa���p��|�k���t�y
�w��A#*&��!(�6�5յϊ��S������o�PC�ƲlPT�	�����#'�
�N*{[}�yK�oW
����O�M0c�<��A���s0Z{��n �F?Ə�n���z�ц9�d�k�q�И�q<Eg-i���F������l�G��}�+�"��{�Rդ��e�h2Ib��].�vOZ�lO㜏Tt�o�k{�P����p�E�n�ʹ���TWa������ux�@޵��VTe�b�y!���3����n�~����j�sx�<�zH{�������I��z���}���xw%��U~��¶J$w���Ϸ�V���h������P4g�	u����ت�Ѽ{pw4�g�nל��ul?5퍉�.�v߄=������[n�h:��0W��y�Ѹ^z�4�j�NV1fo��"&���<o�ep��W����S��()�x���$=ԧ�T��q<U�_V�N�;oym[��K�>1ʊ��3C��Qeq�]�J	N�e��h7�ry0�(�ԓ��z�[WK����~ð�'���;�J��8w~)/d!6"���U��#�q%P�]C��L��A?���c�A�9=
�>Y�!F�>N49�i9:��(�7�MI>�ѫFs��[X�Omn�H�	��7��ԡ�.Ǡ�:�a��߮�wwy�R�����0�ܲkY����W^ǯp�9rRMM�ů����򮻛 D\�1�$�2�E�W�"�3B�r��G�l�h[�X<���a[Qs+�}�Ƽ��G�P���	�0�@?�[+��R��sz���c&@n��}�w qT��[{����X'G�r3�'�[�spKa�&����cŞ{%>�`Q��5>Tc���Ǥ�h��L�Ep�؉B׸�0��O˼D����g���V��P#�	ay�m2��%AE��c��D{���xQ�ۭ�\�`�J�"�ߡ�ל�8���2�D��?
�`��oհ2�y⼰��cr�Q-���vU�(W@uж�J��>�ZY�.K����)��^j���RlmI���J�h_�%�&�W���
��B��']n�#�1lfd�\�v�f��gd�5y۰8�m{�a������ՑA�LP4|5���jC�<gg�L�Oq�K�W���
L����+�(i�
��F���x���������y���p�4jp����E�&�JZcf���s��H�����"�4X��5���*�1N0��_��?��a� �.�Sma����4��L���H��u�P�=�+}��(J�w<J
ͷ�<Q����:��^�N����5f�x��1��s�C�E��0HIj_ρ����B���+(@�~��������ϲ�x6|�e�����/��>��~� �$˰�*nǭ��JHe�V��y[I:��I�f��
(C��R���N� ������֐3��;	-m�Õ�Ե�]Sg�U�j5�4}�-q	\l���⸽+_��u�:�Bכ�e��.�Y���}�� �I޽T ?���M&���l��!@ɝ\W��F�zo�!�$���܀�I�8�J�mzCYY�jCo��&|{��s.lS��2��r�0�����rx^ֵ@ᔔܾ�ֲ�0P��6�%`��3G��j��P�����\�����w���*�/d�AY��1\��@�-5��˨��:�Q�o��騟�(������8l�N�|�)�	H���x�J9�q��꭛ָ:����
m��@U/�,�F�?�P>"�r��p��]��4�)�r�a���Z��TS�AW���S�V�]ʆ��^J%q흔��&�,>��X=7ݩ�1 qz%����V�m���qzp��=ј�@���)���".�!^�	�#��I���1[�w�����?�E��z�P�ɻ�x��y�!�(��>S��(�B���?�a��~�O���i�j���8S��̃�3k�rJd�>VE��<bVH��AP�P~B�չ߼E����Ĵcy|/���AF�(�T�n{������e��s�J���i�4F�7ͅ�cp�F�� }t��*��d!5�AQ�x3�=�7=\�q|�5:�3���3��t�r^5@����W5��%� ��Jݒ���6@V(<�u��+n�G�=��ݔ��T�c�9d�D��Zo�Y�[�d�&\v%B�w�S�,��vg����&$���`  ��t�L�O�=&�-��/�n�oG��>&,=�uE�?�/�ɖ�uG�?�X9L����q���dӀ�x�4�~���'� ��U}2��8����=�1p��9�Jxh��'#;����lR%�v*�\���MGaZ���D����!�&�9��%Y����&Tl� ��+�`B���h k�5�Ct.jp'Pjg��+�5�L�!M
,�x�x���ʆ#�m|�fL �=�j+�qq�9g��-���YG��T�Q�Ϩ���7��z�
_`�Ʒ=KP�$)C��K�R�4NA9J�OJ&�Om�3E�� ��1��$Z�GY`V����&/�J�}���l�� �ZPS��Y�g��d�d+�pv;�π�ۛ�H(�qdKt�J���p)�6z"��87p2�q��5�g/�1�����.���쟥JK��[b(� ��{�{<�:�K_Y��@j�!��֢�ȷ ��9�>*3�:c�����[?�wґV{� s�@FC}~	�"��	iv1/0"�s�Y}�������Qi~�7+=���0_�>�h}.ץ����3�8��Z�e�?�����uBCby�iKٙA���KX� ��M�����Ou���B�F�����s��,������+���YR����8)+�@lZ�bz���Qm߻J!�~�"�ܬZ���-a�LIs��̇s	u���T���i\����Li��yu����b������K����k�ק[ed~��9ٸ�(k�y��u���2�	��SD~!�UT�N��N���N��������M��W}6��]:��{V	�rU�L��&{�o<��A�dtՇ� @#�d!;p.$j����m0�Ǣs������.�}rt|��ϯ�BL��A��>�o�4�d% �&�D���vӡ��d���i�?xؿ}m�[��+��
+�N�\��ϋ||�AzI ����GkBr�`d��Y������;XI�+1uԐ��bqT�{��n+�̈/���%�G��T^�*������}{�gLB��t�#��N������B�����X��KTa�[+`�۟pe{��+A�2� �(ӅH�>���rEF�6M;��so�w��d���(,uJ����c,vW��P�1@X��g�����}ϿVq��۵�0���	�Γ_:x2��j�U2���v~��1��kH�_SĈ�x�� տ��I�]Pښ�v�����q A'8d�Eo>����? ��^�>ش��:���X��򝢓��3��vvw<���
�O��iN����竓1�nc@�����'�YTc����Ң���p����m:�S��n�*9���)��[�~���U��X���o����5P���1(ԧ��9^�rwz4��a$��;�����Or����;	 �����z����%S��OG[�u�i_��̽1P�G�C���r��$�f�][Ć�X_��R�tx��=C`���q��]�S��l�0��jY5������3|EC���զ�Żm��pR���/<�gMS�)�I'\��Nm���&�����Zڎ~׀�,�NP!�jb"WN����s����f�-FU�0�X�e�A������������P*���}L^�N^Ϟ���$܀��C���6��a�1	�	�+����鳐3����]9�:&!��\�X�{�5f��Ƴ�\(sGFNa��P�SJ
�˖:`r���p�NPJ?Ui��H�	!tq�π_� 2m_�'�S.��ֲ��.�4i�Cb
�=��1Q�*]}�A���[p����BN�<�����ֱ�n�V{a�}{ӺV�g�z�"�����D��z��`�V��,4l)����)����7���k29�sk�S^Z����I�3��7ܥ�Ԩь���u��mip����Q�K�1�$�ͫ�U�{�6:�5	d@aNq�bBd'W��G��juA��=]�f�1�}���&.)�/>4�|zw�j�zZɼĥ���}ث�)���m'�H��@�`\՝[y����!���y�p����Qd�׭\饱�Do"�H��r�]�]�9kk�2��#��f!baw��I ���6p�J��]O<JA+׋�Tg�됹��Da�pR����rm$�����MI�e�w�}����;`�mN���>���I��BSB��{��V\�#��F�3&P��Ks9����,4�:���,뢖&%��h.�1�1g�1�#ԒM	���m��b҄0;@�xd*�H�n4��:��j]�.�#��be�xK�+��o=1�=f&�@�DMN��5_�~�:e1�;�x���M�����O�s#Ə0S#���^����%��vRb��u���!n�G7� Ѹ[n��ƣ���B�Vhѓ`�f~o��"x}S6&pcj���Ǹ�:��/�����L�L6��<a=C0�WK_9�|oц
���dS]Dw�
�"(��[�j��l$C���$O5+l���\tU�w��;�V׈�?��S��Ǉ��{e@��ň��R�
�^A����`a�g���#�w�d����-��Ȯ���ԭ6i�M�}���?���l��'��bƟ+��:� ���!��,����������Q{�vd�=0��ۜ��E �jK<�~��!\?��E�_�I�	=�}�~9kC�t��j�x�7��MH�ζך+Wu܎�Y�0��m��ꅐ��l�r�]�����5$�dL\^3k��b�P.p�ym$J������q����N�]L���v9�ڍ��}��qֳ�)�:�u��nb��������fޕl�6\�M��@^t@� �r�O�*=a(TgP��&M�
F����pB0 ��܊��Q�T�+�e�\����;H���*3����IG8���/6��O�z�}�M�k���P�]1�m�Z�wVs`{�p���X���G6�a��ZM�Z;}5�ctЗ���b�|���i��DG�b�{��J���y��y�|��k&�0bH ]Qz�H�k���kP�\55Z�\T0�H��&�_�Ξ���W`���a��we �PD
b�/�����֚��`\�`4(����-�8#
�$���7�Y(,Hv�=̾/�����A��q�/W@e��B!Z�*VBVMv�O��S���1N�̗�g��A��Iy���A���r@ʩ�	9]��m<�BFF��a�e�;ZN�3pbsO�-��U�瓻$Ӝ%xo��������ɿ��!���x��,�=iF��N,ß]b��` �5�K �^�\W!�]�}���u$���WG/%ts���׎�8*K�)#�ie��)x�i������>܆�ϛ�BY�[�݊��U&%\]ʫ ۂ� �`F�F5i�i��
?M;��.3phC$D\�(��f�hAu�)�UYv�$B3�N�Sh�#Ń`P��6b�=��ZG�cWʋO�񧄒E�mHc]J�����A�iG�.b��y�L��Yb��Ow9!7�g<^f���!�&#X�cs��������əG@k�-�uC�ji�=�;x_��
8�ř�':K�P|�
��oN��3:����$&���К�o
��:D[c�^ap[�Yםy��υ��A��Z�Q�X�6�.LӡOV	��	��D�{Y�HG�^���Oܛ<�ʒ�4����71I|�[�������@y�-&T��@AΆ�����J��]����P��u� C�"�_&"��T��jW���u��Fi��{h���͋���~�ȏ1ؓh�H��3�K�x�j���i�#�j�i_���'T��FԎ��bU���5Qb([uH	z��|y��:��X����d�a�U��|y�d¥��t��5N��6С���1l2���JG�&?n 7Sڽ��$����@����,~o�l�!9j3-��/�M��j��iZk��|�lO=��>$�A�(�0�$�k��<�y\|�O��?A���Bk0�E��|�F�*��p�P�a�4K>S2�I��,�Efp��[v>�p�|њ����qř���U�����"v�^�����^���}���7��W��s-��xj�u�9椷6<@��"9|����hg�EJ$��|�%�C���S� 
~�}��,)G��N��Ot���䰣?F�;�#62j�&<���.�B�@�>S\�5;���s<P�J�%��ʒ�Pj��:ࡪ���lt$$�^	&U�*_�-q����]��!�Y��C㾘��"+�����غ���L��!Pjbh�.�m@��{��a��.��!�#-/��&�D4	~!�2�	��챥p�7\P�N4���F9�u��OU�g3�^.%e�{��ޏx1�NC�!3�"���]�!|F��s��k]���� �9!"���X�����w���8"��ό��x�s�š��U��8�&��F����|M����#��d���i,L#���E,�/͉X����h�[�ٸE	��3��Y"r4.�W���J`�r��<�Tm�*��N99��So�A�;���'�c��4EcL��b^����&���.$�8��Kԩ~�bג�<�[^�j��A�:tC��q���V��3����oe�/���i���6���^����Un���M#9潏v��Q��E�t_V ��E�c���b�����9y:�j���J�hJn�OI�a�vMp�eG�,��E
��ӡk)h���x�����3�9뻣,
-���ܗ��W�]&�+ry�s��x����JFi�)/���xN�tN�����2���i"��{���9���QN��o��k��[�E�nfQ�Pe���C�5\	�Z���s��er�,����I���Kn��8t��,O\��'B�K��Ds.��G����i+-Dͣ�4�K.g�9���������O�����/>�$X_	w6\	�9Ȣ)��
����W� 9��Z��)R��9��l���dJ�"��-iD��`-E�f�DR�e�0�x@s�N�ٍ'��/���7$㭬6�Oc����#�*�u�1�R�Ua��Oq2ֆRlX�j�:�I�:ۇ�v�
��M�m��阇nL��02ۤ�g*�fy�������`ɧ6�{l�T�2��P�u��]�7������x(�&#�97��L[$���0�3X�:�\����V��o�	�`F;E�>U�g=zs�48ϝXN$|������o�������%$JV$PC�΃������HwJ���6��2�lk�O*���*릊�2�<����f.�!vu�y������*�a!~�tз�a��!�)�%*V��d�P��q�	�
��8��ι�a�l)We#���QX1
H�/�k��-�G3�;U�M�dQ(|�z��Z�.O.Y���w&���	`��v�3̾Ѻ��%s���i'�$�*8�A���n�*m<@����^Z�]��!S��Q\4��Ŵ�A��5|#�4e��u�Ji�0�aݮ��;����7�]��rq�I�dS� �W�Ԧ��rr�ٗ�3�[�)�"�J�.�Y������o=�&nG��o�31�Ee�v��/���!*�9u�S�v��^;��z}N}>��`�%�ŋ����q�Z�欿�!���E�W��>OA��!�+�#������Jf�_%6�C��..�;a꽜�E��_oǍ>�n��M�H�Rh�%�ײ���Z���y%�|����$6�T��BCo� �͕�����k��R s��p�Z�:C��q�DWj.��Q&eh%�M�7��u�|�9��$�!�x��n:�m94?��c|�$�@�	Rp������k�h��$Y��g�{%��Ԁ�U�@��Џ1���f}E
��~G�c���{��f��z�Ք#r,F�	��{�P�W8�L&x;�s{y��_ ����೺5���8�G�e\۷g�e��۟Z�,3�t`G�����όw?8o�-r��7Y�� �m!0�jUb�~�A,��8h���r�!")���������5U��h)��S�ha���>k��ӕ	[�'�m��Q1�$�.�!F���긂Qe̪�6@����@8��z�dƐ�yF��C2b�PB��.C�&*
u���h��U��;s+�Q!�x(��"�����ҵ5�3�a�(g^��-�^�z�x��U���V�;fe{CS!��)Tيb�����V.zN݋�8y�»�Zb�o�d~�M��ȃ8T+5"B�,�If=<����'+�R��I`�K�[��L&�ª\D�%�t��Y|+�;�X�d���l�7����VhVKL}q����NvɁ��Ғ�}a�V%͆�}k<��fK�
ܞGk�K�U)�2�	ʹ)�;�]�l�S�܂=���Mz����Rރ,�>W3@lr@��$f�_��{-Âi��b��ǖ�[x_�������.�;t+��ut�������S.y���W�0��^8���9,��|�BG3~^nC����\[�����i~`D�W�:�}��[I�j"MV�4�	|�_6t�{p]ɳ+	#r�S�s�����[�tK������d�ݙ-����ߣ�f(��|�|�==�(��^�6t���ֳ�li��-h�%>d��8V� �e��~���D����.>4�)���3�!�\�'�5q�b��N�xW W����W9��E:4`' ��&8��a��[ZSi?���<����wD��8A#􌡴$[/n�﨟�g����ډ�3ۭ�E�K��Hη�i<��
�"4K�Ñ=����*a���V�YjM'ҎCJx�O�� ��`#��{=����e���n�"A���:x�ׅ��U��4��f�N/ˀ��=k����[F>�G~w3��� �-�X��_bg�mk����W@k�g9�㾘z��&e?"��uV&��^���WuY���;�{������7�n�YI/�ń�=���(���{np��_��E**PH��l;�g7*��5{��r$�=���ʗ�m����ZU�T�0X;?x�&r�?���'c��M&9��wJ�{UqY�D�1J0�n>��I��l��)����i�.��ܞ8��7���`����O���ʖ� ��.�IN�bA\�U��h�$�O����A�7)��������&�OIw9?17:��YX�*2����{'X�Y��n�*��R���X�s:�7�Y��]��#v��}�����]�|p8��SZV-�!���d�T��5���h�p�f�����K&aե����q�[7I[�٠É.��I�S�:��vG!�i�ǒ��l�����&�"'�UE�2���̀�&x	,u�����2SA��f�X���1�m�p�QY Ci˹�����p�����TVu�ǟ�g��b
�A�+��
�d�����������Sч�"�A����$�a�|#5`��m��y�3KfD|������4xL��!�&�6_qS��@���� ����G�ȷ�e�z�'[p�M�xU5���M�)�i$�Y��& �cm�{�8�5��b'�.�hڃ�N��Yw?Y2-�G�F��O�\��>���F�6�R�{r�~YN�~J��$���I:,�-���(V�.	���n�~�#�#5���׆�"�i��{�c�:t3"���<u$�vAJ�kcXL\r����v��:�ʫ��G�h�eR�V\�L��}PX���F>l����I�?�8��q.�t���� �y��G���^�ټ��MLg͟r7wr5�?K�)�1}b*�/�w�#4+̗�xP���}]�ܫ�e�Y�[lY!��Q:���˴�߈p �U܊���a�؁!E�(��i_>���n�(��â��am�DlK.�,�`׭bڞ�zEv��~�����4�dz(�-����E=$0��?���J�=,����F�-,�	����wCqp��W�$�;	�%�}�e퍪�+v̭b�ʓ���~6#� ΐQ�W�_�̄9F�~�S��X�D��
�4��"�c\%���)�̌�\�Y|��8�f?!�ޫ(���0�#Q��k����BmHR�B���]6&+0`�aݪi4��^�j[b�j�� o x�3Z��>�����P]4Ne�Yf/�4�@͎4&rg�>�U��w`M����4H�h,2>\�7R^�l-s�?	�ku(�S(=rk�$�K���HS�،�/Y�}��حp0�hn�/�4���uA�^�L������hp���p�9Yz��OŒ�r�a�g�d7ݞ��*+#^16|��'.�� _���!G誊�J�F}oQ����q��Dr��!٤t;g�x��U�͝/����|��>������Q�
���7bp�;&uxZ��$=��}�y�*��9L�f�B��{UP��
��SԦ���ů�|���b�+#W�z�wAey9���kt]j�����ܱ.���wW��ݚ�tHBQ3f�51I��պw%�o�`W�Mg�ua�xB��e��d��ێ]���J����+/����P����W�E@f�Vͅ�?=+� w�� yb�Y�XĮ�z�2���|��D�����Ud����t���+�5�f��zV/��������ig���D�*FK]T��n���Cgv
���a�_�|
�"�\_H[lt�������H�È1��<`���T:����a5bB���U���0��';e�xƚa�D"�s�n�}�a�j�kjy��๢��o��T$6�ȶyC`e�[#�܌0�|�@Ms�e�@"�3��{���>d��(?2���wW0����X�K0"#�+�ն����,m�%��&q@�ܸ�/?[�5�Ϝ	�����0��46�F]'�'�ݎ�m`s���<M��eg˧4�X�naZO��Qĸ�P咆�x$�	��'�q�@
��\��.2h蓺=�76W�����z��(� ��$�(�����?��)��Ъz��#��֦X����}�H���c/ࡈ���D���<���`Q�>`��e�,0K@���A�4�r(*:P|��~�4�9:��7j/"Y��"�`࿕17$&�f��I�V�%Q��(D'E��� �g��>w�D�eK����#/�	)[ t�4Ue�ĝw"#ŌߡrH��pN`��L�y��G ?��Q���H�i؄.�&��W�kC��R�3��HV5���O�4{_��#ur���&x���A����aK6�?�1���t���I�9��vW��6�9���4�ϭnN[#�As5Ʒ��qW�wʩvR����m_���65��Ǥޫ|Vi]�Vְ2�\7x=���U%o�DH�c,�6끟~��Mzvxy'۰甞�)TЫ�����^%XX�����|в̬���ut};���y-0�=2����J��3)����8R��-��P �� �\��B�~W�ԞZ�W�GLK�2�S��.Kc�l3 X��olx�Ҷ'M�e
�<'������j�j�`��嗯�����޴��/!g�pg�ߺJ����x��&������J��4�`z�ӲF`byLj����H�'n�R��e�:k�+�H߸<��յ# ��V�t�XV�ݺ|i��鑽�_,�i�A6���ďe�#�Ч����`O��'���K�\Gc�[*A��٪2c�v� ����N��!$o�e�N���lQUm��K����/���8l={��n ���,r(���p��8q�jU���RX���T�R$g~��Uq6����]��(���,�e�޽kN:H9T��*���ĳT)CF'*LD�B`���w�	vV�!�	�;�y��z����x�Q	l4ϱ�Y�0�l ��-�Ū9)�a2v<�HH?D��\	�[�u�<,Z{��s�fg�S�����~D��4
��f�t+���f��/���ԖRS֚g��7����->�Ƶ��T�{LzA~ї����H�=�9H��:�x-ՅwCp�O�h�!B�h 匣�B�:����(��:�8��*��YJ�o �	�{R���J-��CrA�vv���4Tq�o�Ưr�b-f��ܢ��S�U	9	�<�=�P��R%�Cy>���6ׯǶ���s���~�V�޺�㇔o�/r�ٴ9L7�������E�avZ/���t��i�7p���0k
d�
XΒ����[�0M��}:9�7	�5����������G6N��s��Rn�������y��5���y��:5�C�+���Bm���]��{Ws�G�����⇐��]=&�i6�w'�h%;���7��F+ګ���n�M�T�.g��,a)��!�B55vȡ�57_��s�X*W�=� 	��#)�2���h�@�C���mvq�2�%ڳ)�IP1
ojG�Y􃳏��Y����$�K5�S�
^��\�2�� ��Q>�i�;���Q�j��w��لy
��e�#�	�{�H%��5�ZyF=h�(0��o5���^��u@��E���S�ba��e���n�r�_~:jp�r���뙍�(����e�S�a����o�a�~o&eu�b�zK%���i�1I�㤷��>ސՋ�gK����ZX?v-�ST2y�R�ҲJ����(�MK�5�,h����ѣT�WT�7xY��zms>�y/�g�&nc� ���URq�u�� Mx �ۑ	8��{��-)
G�&v���$
_,(K�~�74���p������d%���	{b]Ho���� ,��\�`��9Ӹ�&K\Ȧ3�<�Y�}��+�m�<�X�F\��'��/�7�2A�<,'}��;U�*����/����Ԯ-��|�cgdv��IK���bpf}c�������Q�A���M�ХY�g�m��.����\��-JX)%��~���Ct��B��Ǉ�`&}�>�6σ�PO��y��Ǎ�r����o6N�Ylc��h<����Z�-����Iׁ�Ia ^p
����W�ڷ�`�B�YK-����M��q��j�N��yy#5����0~
��t^�A�[s2��Y5!z��7�q�d�k��>�Pl�)�5�	�K��nTKkj��6Ϳ�4��R�,�_��bAR:�y�°ع4�O��Q��YҞoN�]�Y�`q\�G!\�����!9������H��ζH��ón&�+o��0�S�Ӧ�s�*��ޖ��Z�&�G֎��AD��|b�yʲhйb��m����lM�ǭP�dp�&����D���ޕ���j~�-݋-y�����Ё�^T�:8ӆ��@R��E���8���/Ǯ�"&-8@�{g��R�<8��k��N���g�]�NN��S9w5*ᴁ�p!�@�q�~�vP���	���ڽ���L
�a��-8��驾n]��ü0�n�Q�p�B[ �A�֓�˯�Y��C�ˎ�'�>/I9*�$��Y=������>��ƻ����x�__C|���E4�eo����b��VWd]�Du�`\�|�3|e�ӫ:��{��T ?�j>h��rd�<����B.R̀��2M���_y�3�[�l�3�?E�c�ƺ�AV{��*&:s��3~i�谬E�(��\?��%�s�dZi����s�	�bL5��G&�����Kg&���e$��:�'������=,0�cWH������@#�ݩ>��Aڿo�Fp��Bn�[|�f$�
ď�2�6�!D��I����{�׆���������������ay|�cf��,�(� =�G��1��6�y;2|�u0ځFE�'���Rܔwۆ��܏>�R�!a���!�K�s�Ya~1BRF��g6�ݽ	���˩�/���P���:�֒��D�_R��Ew�d�z �A�=��������9@�a�XO��u�f�k�+N�-FL�걙0��IjR�,��rvل[ɚ�ht�Ҟ<�;��~��C�j�щ�S������㻵~�u�qm櫻�"c`%r8خb�t���-:>p�����Laj��KpךԈ����*���1zu��ɧ�'��1�BA���� I���Su�Z�
�(P��L�%$�2D��*^�HI�S���p¡�ģ�.�S�Q�T�$���P��4�=�����*����a���';5�q[46B�~7�kxq��
=���9>�-�!�Ҕ}Lok`�5'HV�W�p���)��)N.��O=�
��j%�9�Ώ���q�u��j��e$�3��W\�7'��y[=�L?�گ��{oΗ/�Zb�m�wpd�wRP�@�6�i	ĲlTy!Ng��Hg�cso�[�H�.Ew��8<��J����I)n@�E��vl��oO�G�O�⭑I�FW���]	��ff4�+_�d%=A�7���jK����� Mg�F��=�ۤ�M&%���&�F�@>]q��S�;mb��_K��RA������3��Pjl[Tn�(EF@դ(��2�ؼ�1<�����QR$ {�SSsg�BС���m�`����ZLkN�;6��,�Q��3yH�i��.!�*/#�:�����onI'L0�J1��#�h�`ab��ħ,���(���r�q��z?(T�,闍M�d�>7�,��uj�u3Dά��̃(.�����Z���,
vK^-2诜(͈�h_f"b�[:�qZ|L�	qU���˫�ܓF�娊^Dպ��=�&�e�HǢ�p(�[�:�m��%���C�j8�\!ԋ�Ȏ}�2j��c��t=�^�t`"��D��!�a����nc����"�G�I���yl�����kcWO<�簬����	����xR��O�Uw��Y���F�_I�(*�F9;�s.O�jh�U��`�.�s�Qh�u� 4��sP�H��g1\������3ރ��_�@6�LS�7[l�сĪ��F���<�m���Fy�̞���=,^3}c�Vh�.���Ej���@�/��o���8%l��ꍶ�2�}. i�H��Nk|<��(:Fh�d#<�-Ӛ�ln�T�"Hф�D������zY���ǀ�DS�"~��V��"�D��T�@F� ��p7���ʓ��VZ%ҭ.�N�L���'��D������J�[�Q5ع����Ҥa��7��BF��R�C|N��GLU�/�t6ܛq����*�o�|0�)�~��n�6�ԟ^ݣN���H���(���,��*W��z�e����i1�"i�M?��{p\����I��R��o��+c�.w�4:�tQ!�	�S�UδW*+v��t��d�gqP����V:��nǖ[���]���4�a;H�.�Z6�֊��9ᕺ��U��Jn��i����]{A8��w?��.'&ԥ]J��)��ݽl��U��f9^��N-�\��s�K��TY��2���$�B��d~:��z*�,����\8.��N�k5Y�	zf�i���^}�c(+���{o=N��f;�,m`V[��T�܊ٯ�dy8�Yv�~� ���ڀE��+2�Af7�~<;�t :1@�es)�aFb�ҥ��P���τ$JF���J�`�y��Ȉ%o]b���� ZrMz�@<\��Fj�$s>$|��I�_w�[a(}`�Y���8�*�^��D	�)=�|ITm���n)�C��Ɵ��ҍ?�¬��������ܦ���ox�nT$��E����6��p00ȷ�:�ΨB�?��E�+k�\�t��u�1����7;$�-w�)��g��,��D-�zc��D�_�dT+�Cͽ�˳��Ⱥ����W�5d�	��'��*�^"������E�/�1҈aF��-BӺ�]��T3.��"��}�ĩ([zk���S�J����+�M��]f �b]�=��!�^�3�h<Q@V�����Wع�ɱh�{
γyF�ck�F�h� ߥ��1�@7��e��-|�u:l���8��I��aь��35�����'��Z��Dk1�x;n��d�	�
��-�4�>4�Y�N*�'�`v@_���BS骞^��>./�%"Z�1�֖��8jO���t൚�t1��8��o�}8��?�;|����U2Y���t��w�$�S��68�4�F����:6auE)!Đ�`����nc�#��h���tFXi�H���xgu�c�ږp���U������B��I�$ʹ8�|��s��W�]hW�j��sZ��(�LhFHg�>����>?�ɺ����N�\�W�P�$TJ����RP�tq�U�S��ȕ�O(R;�A��i_�5�u�Na 1���Iq�*,�O-�r���OP��[�=-�U��(�|D��82S�!�k�c���B2p���P]�N��IB*����6"8�V�����`��W�_���|��j =Z���ܢfZ��54�&��Q�Z_��~����B��{V2a���u�rw���!�D�i3|H;-E��*�:��a�S�M�#�Y*w/����j`4p��=����P>�9�f��.£�S��+\GU<��ٗd�V�ZC�`�;��P���Oy����	j`�p5�]���H:_g7Q�%>��%��i{��m
�?�z�F����hEca��0�x�9�[�Y;�9 J��l�S��^$!�l�(��N_pg�?�Mm�L�Df�2���"���K৑�lqPZxA�e�ᑭݡj����w���5�W��WRGc����fY�Ŝ�0i�]�>���~�y}aA	�ѓ�Y�ô'����;8��b�Xy����ȿ�50�a|�j���*�u�0�[��.�Q���	���GIf��j,5���D-�x�G���S������P��;��H�+x�1/If�J�IC��mo�!Ꝡee9k��xo����[��#w�ڤ	�%��۝!yL�r�� }��TEMX�)(Ҷ	�4�N�Į!��K�HA�2�nXT�[���r!rʪ�H�r�4�D2�t��8:�^m��"&�
��sZ�۵��:q,\���Oa--�B�w�������*%Wm@��ɘ�9[����:�&7�]��S�;�%Qmۖ?�0�0cڡ8���Q�?t�ᇺ�|=� J�����?�G�8"n8R#� �� z�u�~��8)V�b��Ѡ�@x�$$�N(W���O<�6��Ʃ�At3������1�"8���wp�H��
�^�E��\�!��s����"Ǿ��"D�	�6����%rzGj��2*=���v�D�؏M�MtӮ5�ڑl��,N/���VfN�SG��{)/�jtb�ߥL2� ?��S�
��3ɭ���t<�+�?��-��d��Q�ꁫ� p=�'��b��nv�^�m7��u��'����zf�Jv���'��ngU1C��"��� R�aJo�5h��  ��6�n� ��/c�i
v�P���T���׶�z�X�)�H^-|ό0Aa5N�������,��Ԑm�垾�����l��oK�6��:���|f�D!E1�T�QB��R���ƛ�dO϶sWnN��V /�Z9I�'��X�X��ͱ0I+�% ����1N=eh����~���$I_���"�7wU�˟zM �;�Nm����pu��n:C�-e�%ŉ�������h(I�������%Z=�-��8�k�]�E�Jz��E�T��X���A�c%.D�5���#��w���=�ei��0�_��������m�8;!���YQ��i�;&� l����)UϩT�O9��"
�^�TAc�Ҁd(��t�许���Y��'Gx�kF�5���� K�����&g!�q�>���~_s1�;����A��W�2V9�IKS�{�'Id������+�5����{����-eO�{��h��}�~Ȫ�I����B��62�	ЃΆ��K@9?����{&h";�r� '���Q��M�_��]\�,c�������&��C2z�VG�mp؊(�c��u��f�(L�ҝ1y�kÒow�Q�͑-�^�ђ�OM�{[zp�R <��B򙷙P+��ad��w�<�;�0���R]l3��~%���l��m����D{v������ �W$����
YdKڨ�9˪���Ӥ�ƹp��U8:�"W��W^�����o�����e����.6`����Ex-��)0�����u�	1�K��v���3�l$�4��%�ٷ_@�[j)$�!�F�h�\�$�h���Aj�yjuP��B��G�U���^����ԞY���?��v˥@o��Q�IQ����e*���JDms审��&ꅷ46�f:�|�D�	���*b)�3�W�k'������>Uڅ�,,(0X�F��s�i�w�|��Ō�+�`��k����Ύ��#�y�!�Yp4�ҟ?)gM@.��aV1���t�G��Ì�j��V�q�Rp���m��GJ؛�d4'� b6jb����e:��,iž�z��;�:�c�d�;|R�kn_4	���n�;/;J�����ܮ��=��б�L�W��n���˽e�s���ڲ
�D������p�m;�l��Sv���/�afi�D��|�&�}�G�hP �2)����B���`bwS]���7��k���!�m,�W���4g�9��R6Z�5V^2BhKMD��*$|59�:!��-�LZ��VГPn�V��~��f0Ek��3��_��Z�d�1\��$��2��ūT*ݯ��b���-1�*Z"QJ�E����J"����\������т��~��2��1y��kD;����/)�]t���ƍ��H�����:�ϭ'YT(J��d9����y<�c����S&F{��kV~��ah��j���{�śv=��E���Ä��_tx�:T�t�[�Hs�r�62�p�,<�����*�R���$�jm� �&,p&�&÷5s9��ʱ��(�4�>�(Mt�f�9�Y�S��j��Z��|�9+�T��A�����p@?�]K�[4_�������s�a"�D���m${=���kjaQ|�Q���\���>Ǯ���-,��*8�Cz���+�����9.n�H�6M\�A��hkp&@�TJס�K�V%?�Y6)ь:3�\���l��\�Cw{��ݘ
���5�zd�Tw�GI�mI�<FY0�3K��Đ��'�GNNſ�;~�� �@I�Z�*��|����M�" 
���)���t�XP0Po5����9�R/�Z\H�;���� �g��S��+"�xo�w�w��?QVGL�����A����Λ J���xh����b��W�X��׹V��M�֌����~�oF��w�k����Z�r��]O^�uv�ٕlև����Nփ�m�,�zo�X�#��bi*v�XI��+sIxⷙ�{�P�Ŏ��פZ�j���R���^c:=�v��~��M$1��A���E(ׄ0�Ġu�$ѷ�7w�*K����'A����Q�?!�f��D�s�a
�=���4D���5�x7��P��D�����D�=PuC�B�Q�1
0U1�9��Ӟ	e+G+oyoH�
`�Tj��ZD��=��:��N	���|��hT��;1;�C���8�7[���$��y3+Uڢ��M�C
��$a'Vo���m�\��5K9t���6V ���8��1*E�zzk6�狊������Q����sqְ_ �Z[ �F.\e�B+
�=����X�84�t,�����	�������R�����{�)!}#�U��I��@!�T�p�z�� !Na_a$���
(�L�\OM���z[�z��U D �z�.-5u�rkk��\>ʪ9=����d�FN��Q��ž�yT
�M�4�}\����-�<��@6��,oDU��%��#�� E��q��LI�N\_dyA������t�B�SO����p�V=���e����*����M�h-�Jh~Z.�2�)�8a�+)���NL��IP�B4���(�6�@�s�{��VtUhy�Eaߎ���d��V,X��ޢ>�j�iI�Y2fZ��}�Aė���Bc��y�7C�*���E����b	C�����X���h�7vʽ��I0gy��!q�e	�y�>Lx6s��^�e�4�o�M2O&� �E����Ez�ׯ�#0�����آ;��^�J��	;�()�8Ε����z��IJ�Di�˹�� �]�{g��27�}��+�ֽ/�X���V�#
�k�%�6Y\x�.��b)^���-�}�vC�<u�d��8f�N��CP�c�lq�6��c�0Ч~4K�0m%�E���p�j��dp����X.:���\�L���Q�X��$��E�bkXՄh�b�l͖�Z�Y�[Ae)���#����ͣ��9�W����T�mw������]E1n�B�(G&�z��a�L�A���l3��UmХ�f�������I�s#O�6����5"p��b�-�����L�3D�\���Q���m�
"@��$X� �X}��I�cй�o���s6�J��6�X��<锑��ƒ���_d�쎍�N����`rE�Ի�B���e�܄#�jR)I�����G6ր1|�u�|��4����O�UO�ew�<�K
�2{�?2k�*Ք�L_��y�:�Yu���\�_���Y�ƚB1�������O����W�w�� 2��e��Ӽ�<�4���v��{v��|�Ҋ�&��M�!M����=ڈ��ݎ�Sci�9߱n慽ZO�e�~���"�:���yE�`�vDy9��dc�z�b�i��q݊�S������\���C��m�
� ���_��_]�fOE�(�L�N�?�W�
�ע����U)!��o�	�ۦm����|Eu݌���s��$�h��]aD=�gޓB��8���;�H\d�1����'��0�L	��h�w:5���]!�I%e��!����-m�?k�k� �?	(���lf���I_�/��e� �ul{�>+�X�ޕK�6�q�g>9� x�����?����P80����� ���-l����I�C#��mi���6;��H�_8*^Ȳ�Ś,O@s�o���ڕ�[Hȹ�#�#�ע|r���j"��Vd��H���vZA��ǐ����]�#32���Q����;!�c�8,<��nr�W�s�^]�nS�k��YK9�+zĤ�rE� y`s�Rq��A������,"�%�P��d�J1h�p"Қ�~(�o[L�
j�hm����ͬUvfA!��mC�Y_���̞����*:���WcؐM�EPN��]P��\M���8���>~����!F���j���/q�֩���g��o)�99�9�	LK)�;�x��J����S9m��q�H��q�b�#�ˍK����UOis^�Q����?y0�V�2[�'���r�r}ɶ��J*)#��z�"
 �ޡJS�
<�g��jO��D����E%o��r�tk	�6ζ�������B(:jx�K�U+�}����_�Z��B��D��m��=ˎy�8_��#��; p�b��:���]�$Y�M�j�[@��[o���|X���F�8̠���N�@�*�~/�/�Z��� �h���f!�����k���
��q��a<xQ��ז�V���QP{O�4J���� j��W0-}�<��6�>yA�,k5K���Ji�����=������H%|�(��<����D�%�j�`Qa5��M[�d�<���+�תT�J�[�5�
̄��	�%��6�6�d�ʇk,~������� 6�咆��:O|��{�up炟%<�QK[���*�
���>%���'��6�V9(�h�T'\��
:~��a
7��?{T���(?����g��k7N��(�qW��&2�*�F�,\��E��EU�O��~$%2�ÛE|�_l�+i�˷#c����d�3�G�7�"��A�x0UhWD\%ϵߎI4º��
͗�7��q�N�*	�}��5��0l~V-"c�m�f�q�#�-��rU�Y+���,�񌋐J7�N��`b����h)��Ρ�ՠ�	��T�:ݐ��-ζ⻹@zԱ�ߞ��R���ٝu�p$C�q���=~Q�J']��jv��D��%2���qDA������e����$3�$��Qm�=���c�,q��f�
d��d�iA�o�;v`�%~�c���K�����['����A�ه�=�Ԣx����㗿��]�>P��T����H
��C��1�`�3ZRP�):��AZ��5�2ر�K����+`� �8M�kH�Գ���+��V:XES@��L`�x������f�����^b�e� ��R������R:���0~�̜J�0�+M������>hK���V:�����_2��݄:W$<��݄��dǷ]w�J�o��Q~˒әwv�"������H�X0�G[Z��6�����)�z����0���A���H������f��ȃ���e������/�qX>��G&�O<�5;�5���}p�
H���i�����|
�V�a��v�M�bm������l���\4`s�moU�9j.���8»�M���8u���'��2���u��Ȅ���_��U��vfΚ�B	=�T`�qX-p�+��M�;���Z� z��.Z�m���$]����v�x6�ă�c�w�Z��	�hj���_������s1Ǹi�;/��'��in�#$����B�̹��ۍڑ����-jRP�k]b#��kѓ]FX�W�S��u�	�![�W�{���:@No�F9��t�+D��4g��˘h���n-F�X�k�_�ǝ\�*���W�g��u���I#"�D��sG�4>Z�c�x��mf0	z��,n�k#u+f-�{�qg(:D��\Z����g���H��ѯp���}�]s���F\�2��
�ﾹ��<
�&�c�n���ME���ݼ�����f�<��G��;P��C7�������[���'c�zA"R�^6F�K%����
�^7I��F���t��lǞD�l]S�@L���R8��������&E2a�(Ҷ��^_;��P���C�"촎Î�S~��]~���XENc8���(�Eha�:]��i.C��v�T6��N�ZW|��,|vkC%i?�� �H��<�qڡ|X^�Y	����3�z���_�M¥xI%)����T�>*�%Ha��W�ҝ����h�1�E�W��=�q���E;���*x�ӏv
+-��'tb�E�A@����ഏ�!�]�k6�w�dŏΆ~wand���Nl���Q�U� pt��)/p�$�]J�4"��V5#tv캉�q��͔J_G��-�d�;�3U���{��
s�;��_Aq�j��4�/��9�4��a��m���zW����-x~>��w"L�}dc塱����X�;���6����]������#���[8+��$�"zuU<U�b��3��X;�B�ΎƜ����&?��Z�4<hp/l�y�q0^�35b�<�5h�F�t� �)b��8
�)����\{��M�Cv�oR?��X�|���4-�{��%��ǂ�_m ��@�T�]�Sm������i���"��:�{g���vw-�i8��,�<?@a
^Qw�I�jr��q�z�/��?��9�%�[)�tF�Һ�E�}���G����J����5Qi��>�#�-k��&�2uUs�F�Nw���(���m4�=�;�%�,V��U�7��qxT�q���"t-�n��؋'`�'�V��]|�,)݂z0��m�|���N�⁲S�}X��(�@ىU��jh��"��^����'ѐ���S�Dq���B���w7��Ў�-ۏ	5�pŦj��s���5���Y� Ё��\��h>�S0�� d���v;"�"����W�h�ԡ���N��J鴒!�΢�ڸ�����a+��#L?P��Y�&E�×�E��cu-��Q���m��<��Mٳ���h�i��V�&>i��Ɔo)V���B������-	3��Wd罸d8s���$Ii�(��<ZB������P9�ϛ[0/$6H�Ɏ�!�I�)�eyQ�˞��>����!g���R��ؖ��݋)��UX��o�Jl~���E�#�9�w�8�kK�\�����"b��y�\���v���~IM= 5��5�
�lě�k������<s��4�Av/�7\���j�yKq,7ϡ}S�i�W���qɗ�����-^���hôNz�S�h�H޾�K�R�'�@�_aG�ohfP��r�<��m;޹ѽ��Ѻw��n���
�_Z5/EKp*G�0%a|<�y��oz�7X�`���ӝ�2\"�Ƅd�K1���&���N�� �B���2�ol-*c0R�8ϻ��U���eA���=��ʙoO^3$ȭ�´�Fڍ^yyq�'$)y�T{V����!S�G����1��n��X瓸'�$Q����P-�%(��/�W$bL�S$�=esv.?�(�����s���0@A�ٔ�v��}�I�s�j�8O<�i
4��m�WK�j�+h!��~�$�r^���i�Ѩ������	+���f�{�E?6��_Sxآ�i�"-!�K"��>MVt�peᙥ�j.�4`����h���;Y�S}�P֚��,lvE2��ψ��Cƌ��Ё�=��2�*	+�tZE7ҳ�����[�kc^**�P���D��\��ѓm��P0}����x�/I�;g�5��_ܧ
m ���"ǐ-s-G���u��!��K|����"]8(��+���I��l����_WMS���Mٟ�(yu}��!�P =ǽ6w��K��&2"~Q'\>w�q�?�\'��vr:��j{�Q�Y�C"�.�}ĳgXX�N$u���.`D�:��u��g�v!�H����s��:Q�#Z$�6B���Y�L�!�9_.�@�BG��T҇> �n%�Y&���U�zc��fUu��9S"?��QGM������0uB��#��-(�� y@�4z)���qG�(��p��3�^̅&���^N
2��
�=��:O}�4q�֑Y43Ba��f����1��8'*a���Ie7�mj3��0Yg�Q.O�c�펢M��:K�1Q�����Zv��i@W$��4?!�%ڦo+H�&�WW\{j��+�tg�� ���E ���Ջo�Sf�b�*��#�.Q��k6����]J�ʨ��H��Ε���_��r��P�)�T��/��/��A�|i��߂3ZEI�9_�~"��0�Ɂ�L+�\���}��~�Q��8(�<,��dPٷ$�p	=-�ַ��Z��*Ky��H=;��}���1�^��zӞ��Ȣ�����������oY4�p,�3G������3x�ޘ���'"V��ng^�с��2��k��DlxuA��O�;�pa�ߡ�.�ے�(����'HZ' "a�9� d��a��·�钗o)��T� �!앵V[W�8t� ���� �n��?��Ps�V8��	�f��A�2 ��@�p��Ѽz7�t�U�#D�zd�Bpm����^�a�6:�;�% p4�g�NE	u����&~-0^kۅ���S��X���|5_�L�fǝ�f�U���T��x��0�Q�E?������<�)���k�K���C��P�� �������^;w,Ò���ϗ�x��־���3�;��,���tb���Q\";H�@<.�I'�Yz|��~�������sU�}~y�zhpQj��g��޶9@�]K-��4��Jl.����]�'B*>�1���6Z ��	H���\����sX�gԕ]�"��
o�I��A�\t)�t��R��B����NO7�M	���D!pRP�#���<9�Q��?vC�U'�7(�qqv.h���Xn������O��U�.O������,�m5J^W�v�Z�ψ2����
b�3�YV�{�aN�
Cp�F�Ii���5K;�g�*�z�m�����|�G��Ӱݾ<U��њ8%��S�dI��#�[w�Y�X�	�3cdw�3=�EF� %�tP �5����|�2�M����!���$q�����3vV���u��_鰽�h/"�SV[����ƴc6#�)���:AW�U	�����8���ZU�����?B^���P5���ezN.\�0�z�n#�z�ϐL���娦;�7��.�Qҹe�	�;I8���_�%H�z�棂�^۸b���f0�&�����*�bq�Pc"��Yש�+F"$��͖ՁN���4*�Z���t2�u�-�����ٚkq]�B�B�-��6���HD�%��A?=�v�� ��\Y���9:E�
��s�[xR P��p�9��c�_rQA��S�$F�F'�*:�2����X�Ȼ�Tǻ2�⧚ kR~��Q~c���e���g�d�9al������^��Ȁ������o:�@�PC�u)ʋ|�(/����j�.��C�)�6])Y3���s�g��pZ��������E�b"v��=☠����U_n��d#?�<*� K+'pWm�;zG���V����X�0���L.[�����lZ�ĩE��5�H�n���ۍ&0ut� {F;��L�y�Ye����L>�$��P{������e�� �����k�����WM$C�u�S�A��E�֟(�$�<�`�W�6m��.	�B��S~ Z�L� :��������l.�%�1�1��O<k��ߺL��n��g����BproaJ�
450BȮ���3�5$h6 K��I���2>�?o� �k[�ح$d�cڑ��2����γ!�.��u4��P(�Wq���@�$�ã��cRA1�����6�I�[>)M�%@e��Y��
��_�#��A ���nt��#�Q�H��JnSߍ띶�;]�L�յ��i�-� =K��b��-�' ���o]��x�3C���`��EVU�bU|c������5X%��^Q
	��U��n��R�ywBti��"jYd��׾��s�E
Rd��w�*e���Uڄ�tE8&K�tH[5���
��� 8�g�Q��֪-��f���������D�"�0� B2B���B��R���G$Fz<.$Oou=ʭ�0ٶyc��ɛ�+9��y�,�[Bsn��`�o�Q�8�C
3�w��=?I��W|{�Ղu/��,�7G0hAS!��2
�Q�Tw4a6�a���zZf���DL���D�8K��U��T���#��ǘ�w