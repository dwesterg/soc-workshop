��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qj��o5x,���*Psl*7Bɜ`������(��ГW<����CA	ÝJ�ٿ�#����Nfⵑ`][A�9;T�Ii�{��Q�[�#&]�l-��9(�SQ�}m���N#nd/�k��r��+<B��?GQȚc���Z�ÿbXL�M�?r��h�S�K)�6��(��� ��5��|��
h�ʏF�Z����mB��_�����H�p�5��(�e���''�ls���z`0�	���P�ahB�b8:�F�b/H�{d�~���7�'@U�n�K���'���at
F������b��	)n.���e3L��9�H��=����^P��@`v\.G�0�~��X�A� ����JxkD�[�d��Z	�a*2��F$zD�y��5��!�n���YŒO���ک�.L�9����Q�c��KA�:W�� �>���غ>8���Ac���n3��0�@O�iM`R�?�Fl4zM�Ь�v�L=�=�A(�1���l�U]���v��W��/
�����]�ؐ:wT�C���|�(;�_��c���N���?�|llS�:j:�4i�s��D�J�PS�
l�,i��tF
�/d�h��֗L%�d}}�ӎ�xrlz��J^q�dUɍ"M���1�Z���@X�r3������@�XeD�,`�0>�c\#7擘����Q�p���W�A��0���롏�~$`*e�
�a��J��E�&�W��q��A@hu&�s�ѐtou����w�B��~#reү6�hs��KQ�f%c���Kr����?�|i��.� �}K�y�����qj=rKO��9�9>Ś�.�J��Cn�s��!tY
���i�X�����n�G�H�̫L���� ʓ�8{]��$�!? �.։CT
>���Mݖ���D-�a3f���JLN��Q�u���sE���C*�>�#
��&H�9�H�qD��7�d�;)q`��b�>!���&ӭ�沮KG˯Tg�LQ� �q��J3w/�5��#"��Re�Pv\����b�)��-�sI>L# �?E����ʦ�qxoSշN7�V!!'M�i����ͷ�49k��j�]�˻�y�E��R�%��g�&#��z�*�cO��q�Ѧ(�V��&���MT���!��3�~!��ڗK�|�q��mW���(O��[eI�@���C�k@�"�`�r��s�C�:����q�Q�SQ�G_�;�\�3����lE|`��T�ɗ����З^�@�v�HI���;l��\���?D)��~��d�F��ʶA���\c��5����{G��lT��#JWh�9������a��I?����<��~���`�w�щ$-�@�3�+�p�ꡣ�n�D�P�w��	��YZ�
a�\3&9���X��C~�oiçE>���(�@E���ÙN���Hf���V�_bFsS��QE<?jR<��56��iF�93�����K�:����b�	����r���Q��`�6ri�b�$�@9��|j�����l��<��j޳��:���a�U���s�3��*�0��0ω�f��{�,��z�N������ �k�Į�E�E�;�Eڼc��G�LE5M���P� �OV���gзV�����#ku�ݻ�8��e��,�輛�_���y<4v��e-7�����D�B8�'e{����t��:��z��P��& k�R�Y�r�7
�*�RT��5B��ph��m�]��bX&<�'��.�{�l���0}����l<�j�^@.�:Z��ë(��j���VJк���DsB\QT���5�2�vi:>�`����P���Ӛ�0��]�R�ٕ�L�g_��g"ȫt �����a�̬�3@b:�2T�������J�1�y���Z� fx%/�� �-�kX�ܒ%{ͤE'��y����B�`C<���&���J��~��OH��~%mÓ�bơ��wK�Wv���IT��v�W���q��̋>��<�Q���I������v��	����z����n��Y������H A�)y�x=�$�3�p~9��h�X�/�\(9��&� X"d�������u��;���M�|<J���.����}+�r3���egs�@a����Ճow01��|Iئ\������(�)�Uꬂ�h�6"0D>�����=����i�j�i}�^�B=�`
��T�/����sTw��*����/7RFB�B2C�:K��hO�����ޓ�O��������3��ؔ���`��4�1���U���	u
zKܭl^�Q��g?����Ⱥ��VN6t�ע�����e�v�%z!}=S,�Z�Tp�J���47�i���,2(����_- (Q�o��o��i-�S�Ηz�-/��,��wdȹs\��J��T����Āl��~��ۢ��i�x�
��6��eX`H�8ۉR(C��~���q��F�G��"���\�>1f���J;��5~�
n��������������ʦs��`B
r�D�����J��wD���{Wo�[,��HT��]�n,yI푲�ȇ��ʉ�t~:��e��B����j37��yS#I�h$� HF围E�Nh��48�B��q<��� �l~�jѓp`7���P�R(�E)�+���4||?H{ ���� 
��q㬁霱B�WEm��r���+F�����<mIs��������8|+��k�z���3���-Mߢ�Ԁ��ri8���c�>=4�Ip^$K��Al>_��i��LL�\�3�/�w[u�/��/�|	��,���z����i�7-5���-��ZY6Mʶ7�+��ym���$%_n�4�K���(
U]��	�d� �V蛞��,/�L><2� ����������ek���d�U0�\�f^˝ �H�n������KA1��`�t��h��o%����{��
x�7�q�V�����> v>�����ZQ{__i�Uc�B�2�9��,)��ݶRl�Z[:�~�$�z�%EH�Y`
��E�,%!�ͧ2*j(S���nM ���]{L,>���6�oJ������ϴ�~&��$AP����������Ao�XHl8M�b�4��s��Q� �%TN$�c��Q�@P�t�[ґ�+N<˼��������@$�y �Y��*��	�]JӱPP���\+�[IJE�a�{� �g�^� ��(K���ͯ���,���!rF���e����SD�l�H�����:�(�<
k���V�����}+�����F���<�h	�?&$��;	Ϗ����[�v�md�2���l0�� �f����b+=aT4��4���������B#5��G5D�5��d5�hM����"�*u�_�O��
nxQ{����^��6�xo���c�^<Fdjt	]��>�pђL�D�c�X73���c�&�����v�k��p+�?)��Ɇ� ���Q�`
����`j����,8DaH�r֑C�C ��)�{�T�37�Gv�7Q�Fھ�����9�oN/�`��B\w�*L{�K����{�y�1uF�jVFu�(?!�B���:/ ��`���l��B���c������f���s���Zݑe�h��B����`��|X��C`c'�nKk���MV��7�þ��P�<1��{)��V# 4%��Ғ�2o�S5'�����7}�;�!�F`ol�wH�
�|D;�F)��3�y`K�G������x����γ��P)α!E��l�U��8�#��0���9פ�Q�j���{5q&}�	��:q{�(�~�ss�9�!��[���}��76T�11]�
�u��i��s����!u~��L�C۩��^��ֺ2�Y]#�2D����SK�����6��3WRe���n�'�mن ��Fy0V�їp�i� ƋVhJa���|���અ�4��-�H ٳ��ۋ��@��6������\�ò�i��^�f!���o�b����@`ο�%�%O����ml�v�{��!*=fc���at�wd[#뵙!��J@����q�ƶ"0'�r�f��s�,Є>I�E�D^��}>i��k3���ׂK����-��,���e�78�4���2�`	��TD���7�7���٩���ު+z���t7Ds�yͭ9e�^�a�v��p��p���=���|[�	gy׈<����d��SJd�"zV��HZE�z;F�*P�>6���RB����a��6���)�*�O�b^�M^�ۂ���(&y�%�?ɼ#~w5`������7�F'`;����+0"�ܮ
��-]pГl]f����B�9�c͐�J�U��B$����t��Lyݶ^�5֍Y�$��B�~��C(J����i�Z��A&�sخc��u��9f~�
2K���@�ӏis=��P������@)�L��3��N��ѥ2����M@�w�@��v[z=��/� ��	�(�祙u�Fp_����ܹ�Ԓ��M�$k��R/���Y5H��������ϞG/X��w_�+$,�E��]�ֲ
I� e&�1�h�y�h}D1�����>:!of����v[�U�&T�6��6��N1�V�f��%z��Q�;�9^ �A�:E1����>>���G���2�+�Ł��]v$��f.>�>=#;��ړq3��-4����3��A��|�>!d��	S
�}�erT#�YQn�_"�▉�zw���~B�u��q�I��RP>.Ϙ�|��N�q7����Yx�D����g����k���(]�����9�"3G�&[�B+۫d~p�R�A	8��QHx/�k�%x8���A7������Nˇ_k�g�D�U�L�Z
�'FL����S���j`���F<�Y��`���Xv��QZ�M8�l/qT?4!�y���� j��������̉�6%Wm�Q��
�����;��ʓ}pN&�U�ϡ^��*(�&U1��@�(��|D΄�����=CΉ`��c|����Wꧺa(�tz;d�b,��v�o�w�>3���3:G�W�K�����9�Ac�L���X����ܜ${N�6N慄�G� �F&)�B�.�yB�
kݪ=_������Yw�I���K�	�l}�sL����N AF"��Af;5�&h��`4*�c��B+O�������6~�_���U��?yZ����)ɫ=�wF��$�d�}&Hxw�K�#�����BjHT#��]q�$ ~NVS숛!�).��y@���vx�M-D8<>F�y��]��L5<��&K���z�d��
��
@��lN�C����*b�đ��o+�c�_|E�G0�͞A�� �Rm�q]�L��p���?'�P�6�~Dہ�+Lͤ�� ��j�Daa���llh�� ���z�����s*�H�A�A"�f��t]�
�NBJ?҂�F���QV^N��){@�%6	&������l!�ݛ����6l��SXH�{��5L3%����~�vzC���	���'�ab���Fe�଴�ThƝ�!y�6�p.���X���F�����v���<�#�.�r�䚏� "�~37z�`t��h��x�sR���/ƅ?h�N��-��E��K!b�H�!��dP�^��sa���0��{�hiь�4��B�-��+�n�jW�
���ݪ�'܋�����^���5�"��c7r�I@�c1�(\|R->���^����	:Ծ���h�l��n����_�<����CXO�v]WJ�<�P]_��wk�&
����o·�=m�������T��p'FMqʰ���?�*�c�\A�m��.�h9R�U:�By�Xh����B}s��A~��D��4R��V�"���Z`��.G��}l��oLΆ%]����<�ސ�/g���^?��'��g�Vɵy�N�=.�J#Ш����i�o�6�����UU����X����\XE��/��<Ӆ�����Fw����~�r[A���Bx蛲I,�l`y,��\XD������i���᧳별��R��j�Z�	����������@"GV%�C��n�`Y�i�N�c��'-*ۢ(xt-�9�2s~�j�GjML^�9��e��Cb��Q1��8"�qa�EF��Fg	�z�����~h��qc-�2�6���6G38.�(zd�)ϼ;���ǌx��[%4d�x�p�^�o�K���d�g�l�{� a��yR��~�?C��Sa
@*P���Ϭ���X��7�Ԑ�I{�����!S�R-9;�,H��X�[�S��KKW^��c�=p^B'��5���M��
t�W�q{��w�������>u<��d��-OΆ�f�\��X(chk��K��C�z��G�s�̟�%�U>I�g��n�4^�y�VV�J���GZ?ytb�/),(|B{����Ppj��:6[��T �Cyj�'�L�Ȋ�ޣ�,�- �Q!C\믱+�Q���_�0��C	Y��}��ё��p5�GA��A0����b��rh} >���"�~�^13P/g?��]^`&t奬��z0�n#��jf0/��h*`�@V�/�f��/ ��ӘU��r\���^p&6=SF�ZH9���هKV���e���
n��r`B�a䃜����W�Ӛ�56O�+d�vK�Cl
Os���$J�3쯊ӯ��?G�2a}������^ηX�&��{5DԨ\�6\� a���i���,����:�a�a	)��e�����+T����nY�Ƀ��I|�x�k�E);�is���uԒn�f�43́D�V��yE�[m���!�Զ��p$%�����{���>_��}ezzK`�w�&�b"q ����q�b1�6�?�V�`u������)��U��
�S��G��ҪiҠ�A�I,���h�&I��MO��@K��[��z�X^���"�P����#G��;����riVZ�0�.��{~�K&��"�~��v�uG>7t�����ɬB�6�U*D�_��el�m�V�M��MAt�_��M��d3%��n���hR�Ǝs]�?b�E�O��W
_>m�;'��݀�Hڗ�k�l�l2v�D&
��A��Gi*9F��É��������΄\/�Z�l	]�!�z�R�����M��q#@e�uO�ExG�WQǋN;��*�-$�JflJg��1�A���]����~����B��z�Q�Ԩ�1ΐ�߫3�{���4%9*mN�mU��#tN�z���Ĳ�7�����G�� (�άY!�{���M�L���v��4|8^| ��Tv�t��3�F�&8��?��'���l/�G^ar��  ?�?ɓ���D�t�� �,9�2Co���/�#�Phe��9�@�]��VGc)!��L�[}Q9�O�R%mq83���*jB"��u��D�=�D��8:n���+Y`�z����l��Z9K����IVtNr�1�R|����D�p���� )�4~��O�l�z�	ӷ��yU�Ĺ�0X�B�R�M;m���p�� ��Y'��J�_�(�Hk�qp��n[�댗��5��G�u�( ��7eA��l��%����D��%e.S)��V�X����C�8I�ׅ�W2�J	��w���Hy��
BJ.�s�"�n��tp�ô9\�XS�E$t�q��s6����
������/4%)E��G�Ò5�.��?�ŕ�A��
	J��X�5���)x�P�;(z�b�	��~����zl���z�R�~P(���5 ��\�o������7�����sv�~0Y�|ڱw��u��/��rj?�<V��^�}p?;t�1>3����C`��r�9����:�����
M�y��w �3��.��l��kJƍ�E�-o��"��|g�mtn�A�n7sk3��
��]ܣs�gV�k��rK�B!�����랠]����Z�C���V\$�f?�H�8W��'��Y����S������V�Bc�D�8e��H#��W�æ��Hg�س���ɉ�E6c`H�q�$$ю��#ᩨ�Ag���a��)��,<&o:=���Լ�ob������2h�@k��,w��v��$���P�ᅛ�άDH �
��E�,Ӊ'_p����A������,��36�l�Q�F��mC���+��a����R��AC��mϺ��-��!�*�]��܂ŃȌ[tW�\�t��sĀ��cB���w-��Ad�_��v�
��9<v����5
�	5�'޹����Y��P�/+��Lr]��a)+}W
]^V@WƖ��ih�s�̽�B�eM�r���pR����3��"���6$O_-C$Bޢ~4^��\�b5�oY!�I��ɞ#I�ES��uH�|$4e�B�	�Z�l�FLvu�m�Ld&B�.���P<<�B2� 6(t�$�֞��j��#$�~�!&_?|�N���~�r2��`ؾ��;SP�M����<��E2��",��Ιc���G-7"�Ǭ�@�2H���j���Yt�E�xˁ�|b@��q_�
���9�ih]�h����ٷ5�Q�v�N�sU���{�τG�(m�>UA*�rK�M8�1dN���16��'z�t��K�O��]@� Pv3y�(A�GoI"�k׏�6

��^%9�4i���Q�|g�\�!�!;N�3�P�W�v����� �:�����uP��{gQ�*��]�Ʌ�@X,��;���?�3��xm�;w�1B�����X3e�m�\�~o%�iN���D�.{;#�?P����>��l����+�/m	o��(����"�p@��\�G��9z���3�B,��~���q�Ć�0���⸶�[���4�`�5��~��I�����c��:~Ƥ���NR���S�(H�7n�
?X@��S�Tԩ�2�����ީAЖ\�{0 �,�i�J{�*�)���v�9�sC\�#��7����&��wy.�An!	lA�U����٫�li3˪+5��jrq�gU�VA��~���ǣ|.(�v`���x�&�%C"���O,��G�`�"<�?�z����"`�}wDE������y��3n�n"W�&@�l/0&/y�&`6S�v�K_����j�k#���8��U,���bJU^˗����be�[Ђ�3�!:hu��ʘ�b��?��G��*�Gcz�U/��{�� �M��a]�JR+�R�X�J���vZ��~�g�2���9w���"�&`���� +�"������v��ڧ�}װ$�Bͪ��l���d-DY��*�n��e"y�"�3��{���@��4�-���K>s�����	��@)���f&��u�=ݦ�ݒ�g��6�<]�%w},��`7o�j����\x�� ��O20[FSQ��3�b��Dq�Y�3���?�����_�������O��D�ȋ��l������V�˨���b��#U���"^�j�;Ѷb:{�%6���׷�~��35�lԛ��*1uu�`�����|�yw����s-?{���'f�y�`L�*���gm;-���G6~�k~3�������D%��.��X�b��_�>���of�W-��X����<�l�Or��S���(m�.i�6���	����Aŷ�-*X�褉��Z���]=D#
t0�'�[��8�zKW9G�Qk��V͕��y��C����!y'�n�N"�y�i(oa<�8��gO�=ނ� }}�o�x,�ƺ�1����Ш&h�yA�?y�?��i�����뒷�����1�p�댜CW��}&QE▩jпU�q���{��ޫ����Y��C#z)?��q�U~���``�R�q����W��^"�Ӡ�8�{�v�"���/�m5����{ب�p�S��:�<���U��]X��*��AʽD�w`���w��W������/ ������b�H��2Z� ��ŕ$����.����5~ü��RF3:���)\}�c��@��
D��/�)p����^6w_w�:���F%���6�6G�3)�����7��i+�'.C���W���˙�����\�͝<�n`�ʻ��<���B��*��k�S�UMʡpM��4N��Q�7��0{�h����1bb<��]�.�#�tz�Ť)��E�7q�o�)װ`����kd	M*��G��_��Qd�	�ֲ���ev�eKx�hp܍��%"	:��
��*�ܭq������#��^dz�`�KW�A�"��[<��i��M4D���~|��\O�k`�k;k	uA���@f��£4����u�/I�1���T��ӻE:S�O
%/fJ������^�bJ����Fk�[��N��ؠ2Ȍ��h�R�[��H�G!��:s%=痉Q���r	M�#�$^�8Ŏ�&�EZ�+T6|H�[�KJȤs>?3v܂a�R���T���e��524�o���S%-���Ox���G��i��p�������}Q��w�s8�R�*��}��W`w$�59�{�G!�cUHLh\w*�Y�1��h[����7���k�٢(��1����+�D=Hg�%ڿ����t�L�D�.)w@�O�D(�C��$��qx�A��uA��h<�E��ES����i�̵�-���~Nq�|� �"��4��m-,yH�Х͡�����jw.c7�=l��Nd�t˚��re��"1���u��u}�z�"[=y�g��C�%y��*$�s�&��~��X�܃q��w�=����,�&?,w<�4;��w�"SM���&��Ժ�Fh�i�S�̄*��i��n"�5\�z�fD�����wE�<�e���������ne	q��,�a=S��R}j){����Ǖ^ƍ��j�}
Z�.E.�J�TtU^R)��=����v�E��F��e]o%���N��9N�>�~����On�N2��X��K�����"W�7a"M�>�1/���w��}��S=��~��a����'n~�\7P����wZ�l)$#\>Y�9��.ii�M�@���hO�F�oA�u��rc�(�<���I��'�\������s$1u�7�~ɕ�MLO<dR߳������<"������g�6�%~q0{b��*L�K�U&�Mk��9b�%u�	��n�@Bi
�ꂓ���6��=`�s_�^$�y�w~`���ψ�������p��ʱ	�?
|�f�Bvbu���s@3f��H*��'tX�bE�u�]$뭸���j⯨t��D�BF�lPv��υ���/��IK�5�SF��W�a�,0;h������#�ڵ���$�GK��-Db�f�b��"��:܏O�qQ+�f7V����D��;���C#lՙ\��dU���$?��Wʽ�m{��Ek���P��/ ���\k�� ��E|�/��ǟ������`�,������0=������݁�F�����2z�j�o�#uRN�ի�~��dS���58g{�b��E;�l�B�2~�YzT&k0G�SCr��i5��C���^�oi6&�T�1ZN�;�7����Y&2�:;F�z�!�㘜,1l*{�yK��h|�I�np��-h���K��#3��c�82��|�& �[/k	�An�GM=v���0)pf��Z2��ǑR�_��9o+4,�'|o�'��Jo��Yt�g1q�SZ0�U|:B.�O�>�S�j�Cs)�j��i ����יb���K�w=��x����l��ڍ"�k㘉'L������ bYj[�ǚ&�3��Ύm
��i�H���u�IA^��cw��*G=Qmp�״�Fa�Y�p������z�;s2ݕ^�?~�k���l�D���)�EH�Y*%�9K�p��Qɓ��X�N��1"F��pmZ�n6���Ni>��%,'��Y���Օ��&�yQ9�ꢷk�����h��o��H�3J�ܰ,[i�l>x'�c�����vk($u~�|"j�Q�;��|����J�8�b#�4�(A*���,/[wh�Vt��D��g�4�����=<�XG��^�|z*�]���W�BD�\�������󴬈�Ġ�k��S\���R�7=w<]�G�:����<0�_t�H����0������b_աN� =���+*�_��_�	<�s�d�����}���s��0��9;kdg�	id5	�	�Ӊ�O�'�	�T�Q�iO�hCI��V)0���GG��*.�"q0��xI�w� �j�0�̜�@�ش�o�r#m�xD!�[���U4���1v��Y�n�`�F4��X8>��%�VB8B`5v��X�! ��Z��ُ�n�`����G�}_$L��@R>�n�cr��(hd<q��3�~Ͷ�(��,IM}���jdd��Z�ޟ�CNJ���l�����k1���Oo�s�.��:$���5ŏ�B����W�8�s�\����Z�p�b|�>N�=3�D�PsR�R��(gp�����"Xa`�����#�o��s7��`I�Ͼw!\c�3Qt�'�W�f����#��]JZ�t�H44G>���?��e�Ұ?���?��7	y�:M_)� �H�� ��D�r��ے���t����vxN�P8�m��y�)����FG��`���F�fj��*���Y��b]�6��0LIE/�˵s�X��d�^K��aPt#}/$�P�P��O���^ʭb�[\C&ճ4���7��q9��j�Ds�,�>ӱ]��1@�1�lTr�0=�����vs��X-ޥ5�t��ng���������ϐ�����4�Sz�+��P��Q���5�[�
���:'0s�c~������-:Eg:���l�⮒k��xL��.�w���@Ł��P ��O]��)��.�"66F�-k�lP)�/`B��sy	!����"YGc��<.h��~��Js���@|��! ,�3L�������w�k�s܀Jh�|cһ�uR�.��`(Rj�.5M��'�Ę���� HG����Q�>C:�W����h���:�?LJ�L��^�[A�<�l �6��ᣟ�ޠ�)*�w#ރ�bF�߯R�z�-$���Mn��`�y��q��V���Z���>�p���Ujzc��o��šA6L�Е��H)x���1<w78����a�w ���s��%��:3�B4{��U�?ZR�%�v��q�~8�.+R�&�=�xNht� W�؈��ܥ���ym6'�I�T�x���y�>'�%"�!�\�]�V��&�J+�T�|~�L{��Y2أ_��Ԋvt���'�����uU��ì捯�G���ژ��^<}:��&��ټz:O���%�0w_���7�P$��r��=��"�;�Z�?=[�d ���*�<�����G_�}E{ˣ����ՠP��d���%��"C�[g.խݤ'�K�R7`�*�>.��i��!�1� ��͑�<��� g�RL��nt75�`�2�n$S;z0���/F<̎���#���e�����T���h��Ղy|�qJ�-�"in]M$�\P]a������2p{J,F�'�!�Y�q��`�%^�d#�;hM5�\���D����k.�mqG�u�p꾨1�ZS�\Rhy��bR������Q��j��YVӈ�x>��C��Y����ķ@,9���oK�n|�7��S���%�
���s�������Ԙ]�|�ӆ��	_���+�b���/\��iP�9�^З	�/�ԛ>��:hG"-�uk./&(�Z�U�QKf^LV�E���Σ^�C����I~w�j���)����Ɍ�����?�2_
ԕ
�C=�!��\�l���\�+9_�)���+,�����r���$H����h�gEc�Ę�/�Kɭb�Y�e���&"���+D�ߏ>��{ �Td6��q�B�㳄�LO��JY�k^7{h�'�.M$؋��D��-���
dǫSsin�Dd�7fy	A�}+r=�p��*��&�����pd�{��2�B�wM���+�\]������/OS����*�i�7a-���9��AE�'�x�T���A��l4R�&�{���0 N�e\�e��|$^���/���X�\���h�C��È�������::#W����P:n����t���w.�2�� Qt�mui���uk|� 6x�����φd�v��;�g\��ơ���$Au|����g���v�����z�+ r/9���4{�ܩr	�a��7��ϡ_��KGmY��g�4�R�7�3Vẞ=��n����s1����O���=��:x���@V��gi�%iq�
��	E'����˒��\�v�RgPc���H
��H����..��b�Q�)F�k��Jr}��Z�iu���-;Z�*�eNj��#�&P�Fg29��o���q���!I.+م/�@P���c� �m�d�tA>�*�f����� �R�[�jw��JʒA�WG6�}�l^�:jXe�ď�X��S�8�k'�(Cm��$w�o��"�8��g�)�,
k�<�}�2r��;ޏ��_�z�(M3H�?��������
���f��AĚ��@��2������ϡ�b�"�g���3>V9�?�W^,B�L[[��hU��|���/6xnf�C��:@!\�ș�jaFq���ҁ�q��O���i&F��t�����|�
.�˧s�'��1�����G�7YYt��A|0���V���L�߱�T�J��oȄϦWnL�cF�ђA,�
�1�j:-��dh����~W�E4\��2F�:m��eDKCyd���k�Y�-���3m\��b�}HB{@8a�����X{do��C�}q3�b�r�g�x}�-i�'����@�)�"�̮t�wD|���w."�k`���}\޴��\�.fJ�2-t���N�J��U���ǟ?��q��>8էTy�aP$��J����h�\v�g�5c�{�UԷw+{�W�ˋT��CԤ���:�S�l���/�!Nu�e.�)I�y�&�J��E+�k���������#c���腨�֠�>Xň��w2�	��͜�#8 �љ#�"I���5��rnn��uƁ�Ӛ{ð7��TX��փ��%�"�j��[V���Q5y��z/Ǫ�=�	�����j���M���1�Y�(�X�a�Kk�x|�j���h�d�#�Y�G����/S]cZC���(�b�p���7�(yL�i&��s&R��J)k=�b����ba�d������W���S�� 
Br2�kZz���t!b��Bv�����l\�����M�CUn6tKB/��}�
�l�k��c�u��3��?5��b�:�Q� ��D�\څ�_q�et���A�����CJ%mY �<�~P��s(�5�)7|��-��S��j�YAїI�*�$�0��C�p-�\W�V���H$dg��DmqVK�2����B�n�J�q�ĖK8QZ7]<�[!ń��ZL�%�ް�C;>Jk����u����\��R��>�gWؙYL�Nm�"��X15���m+-����ZDʁj�w��c��o�!���Օ�p�4���e�E�k�g�ˡ4��գ�q�,##n�]�@�R��6D/�h �$w�#��3�ji7��B#�Z !��\�,D���zP7�H��q7�D�s�N����3��cU�0$Z۲��,~��{��-��XH�J%�(�J�/R�W)�p�h%���%��~x���� Cp[1�b%�]T'���OAY�씩�\۱S����G9�X&�`l�����-����{���WfZ���ì�G���s��dL4�`�.����nv��\��Z��������t��X��<���40cN�rxi{}q[��.��<5�>��0A?	��9�	)�m��~+e$w�P����6D��z��<������io�]3���r��es��^��'�:��5�(!����撆ڟAK�����?��ߍ�,G>���V�Պ]ڋ\s���P*<��ϞI�VB��p�.GԸ���`9
%��*�)﹌�f���1�Ȇ��~\XE'��e����e���W@�����8���UP�#:� ���C�S�$2��γ�5I���Ϭ��hȲP����ԞT0_����$5Z�ݜ�υ}��fa�6��2o ��Z��"n������n:��n��]����*�'�S`ë����#	���n��2�V�ҿ�R��T��P�Wt'^�䐈�b;4��k������_�P���{�6#��O�6����/�f�Z�d�_bi��L�g�f�;�r*�!nxUh]�����i�7���iZ9^��y�q��I���GS��w_���JL�H���H��Q����X�A�(鱮̉����*i���e(i���Hu0��a�n��E����o
� ;���TT�Um��{��o4�2�\��5z�a��U��&���W�J�"�w����we���W����6�-ꅼj�#��+�`��M>E�?�#��Z{u �(Cl��dp�Zg��i�C�O��:�K(���r�@I7���j�$<�G?��+ɋ���9����~��W�}C�J�O�.�WՏt�_ҸTP���x��?yY�HP�l��W��L��K�G$��0�ػwg�f:��@T�<��l��r�~�Y@
��o(�E�GmƝ8'dP魆�אm�!��7Y�x���7brI�F�x!aҳ���n��;�Qٛ�J���Yoǚ9��E�����#��/}�'v$��Y���jI�q*�X�ax�v.�8�S.�3G����~���tm�s�_��c	٨���&-�� 7fL���⊔~;ݗLM.F�О!���U��J�p�3�A�o�S��R�9�ä�<���z�j2(��E-�'��%���_��Q�I$�$�YyN�M��j��z�wͫ���ThY6hC���hm~hz!����U�r�*�c�l�J�Է7\b#�`��i"}�~�A�R�(kY�x����?݃�h�2y���)��J6�X:�j���۱�r��Q�J���q�5\�ZoY��)�V�3���x������c[l]���(�*�j�C`�����x9�g�+�x]�M��F�I=���L��	��i�8,��10�5�$�+MV`������5��j/Õ��Ĵf�N�^'D����yP�g��h��Q�E6AN�u~��y44pc�{3��M�A~y�_�\O*��V������p�A��f��r�Ф�����ߢRT�S��,����I�-3k��<��tŇ\#&�b	XS�SI�t7|8ǻ��;-��1]F#�]�с�#������8
�u�ڽ��+v�}��g��%�H~C�Iʂ���3��y����Q�'A�P��],~�����-S����b5]���Џ3�P:�/d\�H��7��`ث̅C�6�'=����A���;^Jo? �����0�P��N�h���Y�Y�؏�㸸���f�Mf:G�x�HO�m��W�>�>,����x�4�9����2"ՄﴹG���z�;G���I�6��m�L7�gP���LڐF��o��>��埍���p�N�Ϭd�ފ�i:��/6��կH�.L�n�ai�1�󖽞Z��͌��c�������l���#�!����u�]�u���Z����]�d&�\����J�)��o�?�~�]�W��|,x�kaI��2a��V�p�uD�t[o����ܝ^���.r�H�߳l���Dǻk �y�,�w�z��;&�'���q-o����¾�u��4��F��luQ`ֽТ�T�<�Mv�;���N|o?�ڏa\�@Ā�t�r�d팹�1;�H�i�H�V<�/&j�W�`�
�~(��㭸�Z���#�p1:\1��ȵSoH�9Ax,3Y���1�^���C#�XIӮ9):�`H�� 6>��1�V;��� L�EQ�P�1�=�\E�v�D{|pĕ2�5rǹ���rt�_�
�`H����M�����Gٶ��&���M�{�N�$�S��n�
ڝӓ�3�ГK�#���Dؒ��eO��C1_󂌉�SJO�N��OX":�$����׀������%���Ą�,�aؼ!%2t-'�
��1�si+w"��,B�X(�C#>����F�:c!4u�"���j�>M��Iu��j3�n�~��k���
2m`?o�D�2lG~��e�?C�)�y�oSq�����l��(}�ݿ�jW�>nc4�^�(��`V��F�hT\��N2�W�&X�R��G_�i�d�1�QK�6ӻeV�Әi�݈�q�; ̓�D�E(ѹ�-8^@�j̖:`'�v���(
�:�2����G$����B@����h�jD��ʮq7x<Ag����x�}}��D�d�(���pU�)��Q���'Y��)�Ҷy�p����3�kS� �f�9���R��R������ 5��6���W
(-�f2�Lꑁ�72��`�\��@��.��]�V,h�;奮c����T���t��b�l�f������<�pf�Qr:	�K��K9��$sӴ�S�;�k-j-�X��މ1�h�k�N^���Z�$�u�47s�ӜdS�K�A�v��`���Є��@����䑅q��+p��fa_K�󴍙k����omG_�g Uq�'�%�wM� 7E��76dzg3|i��/	;S����=�4��O����RG���K���0�-�_ �ݨ>�>)!?=[J�]��W��뿄>%ʮ����k7锡 31�@@�8��7.�L��1$�ж�fĖ�GM�K�¾RA���K������G��.���R	��)�p����O#�Mĳ����r9
i�J@EcS"���;��$�b�"/��ǁ1m1|�<���Y`�O@=��P��Ϸͩ��y0}3qF
2�8�X� ���F��t���B�:ϯ٘���Gl�������o����
7BQ��a�A_�	jL&��>Ú��]�j$D8q4�ظ��ʷ$k�?��ө��\�G���X���u}�_�P)��H*��ú^�/�@�F(���ҵ{P`5�_PS��o3��k���x�v�>����M?��F�`�65��)�p�j�;m��,�����}������)rP��Q
k��:�1�	�Z��_�6��+x�S
�����$mmϬ+6�.�qe��]h��	��[�����.��Uݞ��`����3cw�-����>��%냁��q�V�)[>$(��m���Z�1x�{x�D��� ܇�~�:�G�--�6����˹�0��vJ�x��.vf��m�l+���72�O�-� ��W�e���VГk!���	T�=��⑳���8�m!$l+�?v6�m�,��-��k�o�`�#׎�C^�])�`|�e٦����u��鰴'�����%Y��g1QzEXeRQ�q�?64��I绮s��y{t�K�N�|g�5ԿxޓI}9�+_w�2���)�^Q�iLS<� כ14gٚ?t󞾶���dYi���;��<{�+��?���M�XAP
�%�X&�w\�f ����i9�M�3H7�ьl�5����[�kz�� J�ʽwiE�'���B��fK���o���r<��ae��yB���S�>Tb�Y�4{���@mdg?�Oy�
+ .���=[����La�կ�ue�]���`9�ۗW��,B囬���TŹR3�������$��e�W���M
����$��H+�A��*����ܷcW�A���0�~!�C1j�A���tv���cgԒ-n+c��0��P	�kB_�X�\�k��*�mC`�ڇCĵ�N�y��I?E�%�X֕ˏ��p�m܎���^�%& M�%�$�Жm�Xo|X��+$��|�[O�$���r���=^{��`�BwV�~��6��.�1�Ix�qY46�)�3�(|h�7S���n~9��L�v0��/7'i������?�LE���t �R;k���T��"��3��7$N��:0�:^.q��Ze)�`��1�ٯ�7���~�_R��<|�K��2���)���^��B��}K�3��O4ԫ1�یl.9���2����wF���Q�b��ϛS�ʡ�窤];����9�8�m���?��߳q���.��X�a��v	��N���yW�.~�h�E@����\��ӆ��t�"�:����P��w�@�7H�G��u�B"�E�D�Aj �T��]�R�)�_�k�Ly�D�}d�����:QVMCWV�(�|6�x�'���'jd��$6w�8jo�g		Ԋ��R0�$u�:zE7�p��ϲ��p�!>l�����<��^\�cS7�_����hޖ�V�?��őoV���,l��a`�QEĘ�D�rv�I��BtҒ�R��c& �q��??ey�{QA%����H!n��~D_������,���i۩q��-iǰ�{���8j�S�ҊFN8���?6(@�i%�x��@�u�%�����L}-F�И���A)��l%�����͑L��%%�Dg��ț�h��#�쬲�B���P���]ޔ?d�45泎�""H����|�o���ܺ�o�6��f����[*���H�����\���r��$tU;�R�|�b@���*��vw��&�p���vVt��NԲ]��%rR�f^@!�O�,_��1�۪3�&R;(D8�e4uJ+��R*i��t�[��5�~7�ҧ�����`Jy�,�9ˉ%]�} ��y���j��R�a5�8�^�g�H)$V�+�0\k%�ț-E�
g� 	!H��F�]	�0
%���_.��<=�<���_yx��*ѣ�{�o6A���Ys箅7. ���
F�wٕ��ޒ�Z���ަX��Qil?{uā���������1I+b�'��P���wBP�q�\���GT-�B�k�a+;c�my�M�5�
)G�FH[S��p�R�Gm��c�b��fvjK4'�3�{���F��JK���;�3>�iD[�/��J�Z�'�x�O��3H=[ؤ�5mod��1x�[U��i����f�z��L��3�bϓ��B�7�}o��� Y,h�<�#�j���\������;(~'C��V�<����}���;d��͡�҇�d��D�\%o$_z[����=����t!A�����<u�p%L*��k��ڛ��gh���g&������4��|�+
(ȪD���S�C]�mӶn�]�������W�&�����S�R�J8Ol��'9n�K<(t|��ś�oM32p�w�]=�c�'X�{}�A~(��B�~r:F��8�}QiG�C�P��J���d�X#Y��]�)��K�����iu�B�f�~v!N/�9��H��O�TS��u��x�>���$�����H�S��8;����iz��./��8��4O�d�f���a�6�G0*�����i25q#�{-Z׎�����J�X�dk�j(���i�Y��I��_;KM[���_(�b�Z�^D},F�9ʧm�).��x>�_
�RQ�X�h汪+!~�S%$�U{��74��Wv�|^�X�cۈ��b��z�1Z�{��9�����I]˔z0�=��nǜ�#Z�wb���9���� �'���X�eu156���Ҁi9jD���< �ʞn��_�J���.Φ��>T5�$޹��$f���~Q����a�b,��J%�Y|aF�+�?t?�n�	[�A�����S�}l�Z�N�t��?��J�<��PD*�N���D�7��#�p�""a��sՓ�D��8�=a���躐�6:��ߓ�p&ѩ��jwF1�V��\�J�W`%�]:/1?���c��/5��p
������-%�q��P���`4ǹ��=K���Ɖ��;�U�����s1I9���/\Y�c���gH�g2A����]�������Pϳk8[N��]qa}��t�`�����;Ev��R
a�^|y�O_����a��]�?$���u���c9>��_�E���2aP>>OU��Y���#.W��e��T�`�Ł���5�)�r�+o�vm[��YsZ:$6��(Am�1�a��C��C������$���
��C5��[m3-ϴ'Hi�Y���Kg�N)�IX��C���KZ[ }���z���c�4���\Lt3$34W7���\���Kn(�H�M��)�̎��2?;�M}��5>3_��F��ը�9Wn$-���.{	����p�����L2�B2u=-ۓ�l%��Dy7���ޤ����(���(��4%&�γD���%�7د��]��7n%&�S桞|��aN��[\)d��S�B���Y�~�+HK���k�\;�Bz�g��x ��%j�e���P5������k)[�)������s�%��>���|h�S��ߨ�Tk�8�4m�6H�u�^I-z\	$���\]$V���V����^����dَ�,E�8�\��>}��������9Ī���wIՎ�s�?�(�-��а2K���q�U�fL dꠠ�<S`��V�|~F�.鴲B��L���q3��A;h$ǳ���G����[�(6�L������+Cc�c�#���O��1^��Ct����*�0�M�i����#�V���q�b�����}���mL�������ZX�}���jF$O%)Q�y1crR!Sb��~��)��fD(4b�Q�¼���Q34�%"\��U�wőK=�i���[��SO�1�\@"Fc����َ6�jjѬlv���i�0�%{w�\Z-��f�u,(/���X��rL��ꪨZP�"�|	Mq�.��W�0�08��'�j���]=@��#��u�A�?(-�R�����D�*�3�B�����k�޶���Ez�8�,M!��$M$��|L0�nr�W?Wl�S�&aY��r�����ۂe7��rQ��90���HY�US�b�3E�@9���ˣ�s�P�|�n�&���=�ü��~��� �xP0��C(����&�u��SR���7���w��<:���:8��>��3�H��K9�Y
�9@�n�d�S����9_弈�� ��%fE}gi�b�����C]`�����F��R�][Bۆ:,�).��fvo1:��R��(0&N�/ 9���'�Z�(��Jn���S0%_˨���I��pzp͡�����a�"����ҠU�����]kV�[��)�Y0i��Lj53L�H;[M�x�Ը�E65�BK��5�C�A�W�65��_^21ŷW"���"�J�N� Te)Öt�V*���p�V1b��_wuD�8"�����]��)ϨzI��Rw� ��Hl�߬Kz~K#��.yo�!��Gp�
B��že�3<lm>W~�h##��@�(��X;m
����[(�	�|]�o�����s2��L�CӤ�T��|h�B������ �<|�Ш�4[�gt� �eT,�]F_�o^~̉/e"E��O\���C�T������~�S1�gI>$HKp���c8PQ]B��l-{A���n����V��*@������ c��s�L��M����V��3{>��O��l�d������=�@f���9!�(�l���[Ǎ�A���݂� :�ed�ѐx� ���
���g<{�x谾�]��([�=얜ڰi�v�;9���R��vx�����Um��Pm�iP��Ԍ�Ȉn~�˛�?0�Pt�V� �_��hi��%�O_��4��; �?�z��h�������Ox(�f˅��gw�5RA�r(�5I�̐��A"�i�뛡{���>W�Q�q�S����_̥�V֝*g��4R�<5B�R|�`6�|[��O8H4�FM�s
�Fȭ;F)�h���ҟH|(v7`�ԃ>C�/<�8�'��+�cܶ;R����C��j���#A��A������j�H\W�㘴8#��產���z� Y���tY���8w�-�$a9$�D�
�
!��Ϭۺz����򭶓�k6��g������^p��شH�=��+Ő����r/�\�@#3/8�`<Tڿp��:�p*)黍l3$G?j՛L���r�b8��Z��Â��?��4�ͫ��|�{{^��ʊ�ܱ"{u�&r�	E���:�����h�5��[j6�Us�/9�x7k�FD��%��y������j�#]0t�l�,�0�~�w�;�z�Ģ��w�s��Nϳs�0Ėp��5��h��Q=Me~�[�;1�����ؤ��{�2� ���\i�!Ǘ y���lCj���n���À?�$+����b��x�����.�wOz
[_���m���&�� �iZ��Uj��#S�T��֜�4��Qq��U�k��Q��S+�~�=�+�kY��nB+�6$h_����I^F��U�o0�R��˪����КSJ z�G��M�dO����L��;��l)7��=0,g�L��D���R��؞@Fȭ�(����`0H�+CHw3ȟ�xA$����93����\ՠ����|fL��/�|{���.���aZ7IQ�5����í���ZB��pz4m2�I� B��Y�Q>��y͓���ܒ��L�@��Nv��o�ۅ�
����+a�T���N�7�F�C��S k᠌6gO�K��|Y4x�'�o=-8Rl��'&�����馇n���%RT�C��- "�Zc��\��V����:jXTY�2zq�� 2�������Y���X2��WHj	L}mQ�f�c5�*i4���߽��Z�ʶ����3X��Gɯ�m�(�g7���ׁ~�mʽN]I	�U�����W�����Ul�;	����R�z	� n@@@�`g2��V�g� ���?n<���f���CJ�%���?<��L�M�P�yf�B!C�����q��ӶL\=ػ��BS[�`��|1S�{w{z���@-+a��J�@��;@�،|��a �%HJ���/���	%�M�_�IrY�h��F�ȓm�� �`�-�
�o��ª�
���`6���E��u5&=ȶ�e��6�Ɣv����l���U�>)�=�ds���w�l	9�2�h��)��FJ��3�퓛PT{��r�"�ŷD�"�)$5o&q@�[���񯇍��?�s-�/�el��%h�G�@��7�3Քl=r�v_�"�V��^N� ��mz�;:��!�oÄUc���+��5��獬y�y'G��%!���Ș�^����{�N`"o~L��uS��4/h5z�JFS]��O�e)���۪}<)j
~����w7���p�p5���n�e��a�ױ_S��ݖY�����*���*_Q-����)r��A6�Q��] �t+(fܛ�<���|�4�9�x�y��;�{sIh�˻O�`��,A�WhiL�'����g�rXD���S�@�E/�O������:ۄ���մx3�:Y�ү�2Tr�ܽ]üsQ���>X����|����음$�v/޳P����wPZ�S&`��gy#^���Y��ȑ/.jQa{��bv�@�����t 8N�QΤddΫ^3^�Tf��'hR:��\#��K�K�)q�ZU��ň�O���H�a��$���D�O�������`���\�y�@��䅽���#r4k�Ks��t��=ĵ:�?5�u��dg�~_9&��{����뒙����Nѝ�(e�)�2��cw�K� ��
���Ҹ	��~�E�<d%]�N�HۀN�z =��w^���g�'2�@K:+?����#�j0>����V�b8,d�>
.��Od��a|u�h���E��IQg��y�,���L�R��|���Z�Dv��Pv<�	e�1X���EYʂ�-�N e�P��7nt�H�xkHJ����tgݣ�wWH��a�bMOg  �]��1p^q:�0k�)���4\p��~�Ǆf�"D���3-��0���`����+NT�с�Ē̡Ε��X
d����] z�
e_��Ѣ��R�b<���܁�۹�f���V�D�>�l]t9+e��⦧�
o���)|Y�����F`�+��YY%���+�w�r�H�h�!���5$��k��)�W�Q�� U��E�Nwm�.R���v�-pl{:ls��-� m����dm���Ns"㎏��5���M�P�g�oLS@ [���١,1���8���0�O׏�������ի��9RQ��{����Z�O����ѯ�+��lR�!$?���Ue聧�L0y�@ԯ�p��}9fY,yb�D;+83�ĵ7���.�������="����Ht}����b��ӗF���]khg����y�#-��qn��
�F���w�%��`EDM�P�x�Իv�<NQ ���:����}N�b�X�3D��������A?�_7F��݅.�(��)��{��X�4*-7lF��A��������L��yi��@���0oM��ΞL)`�'�ԭy��;�e0���
@�C���Q��n���f #��ǎ���U��:�q/N����r1?���"��J��|��%H�(Inɷ'�9�߭By,��E9����6�i� �@p����o�]�~~��M���(|�� ���Jri_8�:_Hå[��L7�6db[Gz�C��"�%nG�4b.;k��u����ũ�H�e�|�!I>!��׼fs�嚶;�Qӈ�C��X�����n](붢���ֈ�w/���F�x�xyf �N��4���f-����<BJ6v��iàqF᳣ɻ�����O�d�<y�@�
0���ޚ�s9�Q��ve�������f������4���������ƗLxz�S��p��ʏ�:B���[��|qSi��;R9a��@����Y��_��l(�Q�Ϗk���x�u��>M���[ ϶8b���&N��r,{�R<������W���I�&�"������w
Oݳ~M�7@������y89˞ xQ;��B�p-��̨_-DohƑcEb������߾ٻG�!�.>�b	��sg��H��n{4`�����}����Q:�J�+�*�߷q�����l�a:Ѹ�I/���j�C%�/���@�����0��Jf�űQo&D���},�V���C�����dQK	ZʺB�Qq �b���'�0���`,$�XjGz�wNmƇkU���+9��'�ɰ?�E�S
�<�Z�&���sH�䗚;�4��ή������>'JO
'��q�[�׵�!�n8Y�L���?]�RSϚ������P��Ldbc��M�(�>L}����g��a���~����A� �=y�Q��T����؇y>@�*��/z��>Z��bb�T�����I��lO�(?~�#��2A?sY�ߔ�{BA��f`��@|�Z�޴Z�/���=o�$����f����@��q�7��\�"2����q<�"�K�T��FX���5��N����4�^%O��ϭp��FUy(������(�.���GS�^�d9�Ϳi����\���ů٣=�,�_��漡 ���X�m��ek�5��c���T��n���nnt�ِ�cM"K��O�]��]���r/���i�#����@c;��,�/����<����Iv�-|n�(I�<�ү�fc��,�e)x���|?�a��!�#~C�!P50��6�H�y�M��mQ�9=_QH�1����
}�׹����l��W0|u��t����X���X�-�($��j9��F*�B��s�9s2� ߜ��#S��4������
���F��y7�$��_`�h�8; �{X�9���w��,X��m��0�ae�Yļ�({����2��>c��W͆�=��\Bj�{�ÒN�M�>�J�`��fY�P�y?��B�,��W۶�x�R�T����#H)�y�ɐY�����tm{�j�l�0<$�Z�O�a	�`����IO��F?.��T�� }+�O�;���> �#����W�M�$��+@yWs]|O�3��RF%9�ߊSt^�k�B2 M7~,	�g��-�E=�
aS��u�2����;�Tz��I;����ߩ��M�yy^ �cI
�)$��9^�Y�X���Ɍ -��b�y��Q��
�`��O"~��6Z��m�H��xK��,{��y�iny��y���BjKB+��i�K�$wa	�v�_�Aw|Y {�pN�c��w�\'X}a*�Rw���縬�E]hm �Qǧ�Ώ>�"<���r�dр���h�AKǲ��S,��{	�c�&[瘻P��cT]�P���X����r�/�����W�iX)^a@"��Q���� �1�D��M�����o-�K������a�I����cB�o"�^d�mF�2wq�̈�0v����s࣐y���J�/����h��1�[�w� ���k���qA�E���{~�G����NՐ}����b�K�g��
�M߆�vs��b��ʍ2#�\�i�I��	�o*0��u�`�>�
���E�<���r;��h��Is'����ƠU��T��|fa��	o%p�u�Q�A%Ҝ׸i?�H���SA��������xyr~�0D�sY}"#u4���<��{���5Ͽ>j����\��f��f���z�ҹyı�Vi��0���Vc����]8��j~�X�T��=VVs����aM���:@$�RTj���S�E�F���F��<����z�.�K�����#�t65+��|rW龰 �a1�Qq�_ٖ��R)UӬ�p�|33�}�.�#�AV��;���
�����T��ER[�Y�7� ��W�ŋ�&�Bk��q*���>%>�0)�.��^��b�h�X` �.�G���ZS`��lҙ�|N�I��8B&9d���ׅ�M�q$;�ң>D��;|���(��N䌌�jQP�P!9�582��Q݆?��_F��1��d�F����̧�Q\��L�'a� T$Y[[��y�(�`�B�����@TCb��O�X�5̨FtrM�M/���-ӗ�o��@�)��l/d���wi��;�F4�b�v]R��9�'��~�T���=��>v,2��hJFF����;�m�'C�N'�a��mCG��sǄ�fG�y,퀅R��<�}�.�9�t�0-n�8s�q]�ඩ��C�Y�ҿMZ�C�d�������Y.$�Lc7S�=:���S�DK��j�47��Fm8瀤��x�Ҳ���9G��<f�����}��`EE�X|Y]"�ز�I�2���>��i?8��n]p߾�:pz�g�돹j�h�<i��=A��馵A�B��z#*�>f�}����_6cU�-�R�L�_�<���ﻕ�����iv-T��S090k�UN��Evc�����jq�����1�^��vזؑ�
F'<�n�e�&_i����wX�b0�ή?R\e$��,Z�ʑ��L�	Ѱ(:�u2��>Wg��y����q<;��pU<�߶���B�^o-����i�P��1���o�6zZ�����K o�!�g�2��D�ݶ{?������a��p����~�}�5:�o��e6t��z�&�&h�����K뻺/�bE��l�}ϧ?g$���G��l���Y������ca� �����R����7]ɣ�S�P���͚C��Z�jRt�2LbI�]�t�n���������ް��Ku����/�%�D災��#���ԏ�g�w�	^�j	�g{ ?'�or�߃[���+Ji(��~�#��/E����y>f:�����< �T��gG	qZ&{}��K�,�@��s�i��/�Ր���F�#\ӟ0�ޘy�HsՓs{���������n]��%�5������~	
k鴉_J�^4��a��ܮI�jF�Tt��"�hv�b��N�1Xk��[�<����
g�xKJj�v���Fr� V�����`S�l|��H����r���*W�)B��B'��H�#E )�u�e��{��ѪjM�����`?ن���>�
�$�f~xNo�h��<CEX�ٟB�H�x�� �غ>��`�0d�蚻;>y�b,��ŴU	7&MW z��3������I�a�m�W��\��>A����?�8'Nd-�����z�����Y�����.*��|w��ӊ;�-�XTNH=(=Oa�T0ֶ*R5��������������� "ހH��Ԓa_H��
/!=5V��w����<��nL|�/h�9�X�#�8����PQz1�\k��QxW��0É�E!Xэ=��lN��'�\bH^�*_D����9��C�]�W�,Ddl����!��ߌl�����O�t�r���;�*o5e#MU�m=R��s}i��� �,��0F0
�~�΍?6x��7ۣ��Y�D���%b��ހ�to��
f��s��Ug�� �����q��sq��������+um*?�~�R��$����,*RY+%<�t�ҌZ�A����9�_�@�2�\d&�	�E8�D9���x\�#��/�c���1���b�SA����
Gؘa<*��,G��M�f)��k�(;� �"W�4
��c6;A������� REh�9�g�5K�#�2��w��a��Z��������Zf�-�uUI��~&u�����z����$�M��v��@bn���e}��tǽ�z�`��S�l	���Z�a�Cdd���1�A�> �h���B��p�Y	E5zc۷"��D�bIV$&cvk�-��I�vT���.sA�1�v���L��ā^rz��U�) ��v���D��:�x"�~L��kvU�Yク]t��rP�x�Qu���B0.�_���Y�j5o%&�	��ݝ�)�o�jF�v�f��7U?��o�l�eU��������!/�Fs�G��؜24�l�Y��@d �t���S/���謙�HG���U!]|D�ykcj�%W-Ǽw�#���|�ǃD���,�O��p����<Zm�ߎ����8P6�SC�d�+�������U��B�{�s�m�k�W��|���i�L��Oɢ�m�r��&����^r��*�e<��lUC:�D�v��`/H�&�Mm����^E�"aG��N��;����0�C
W_r���if�����
XpFP��W���&��JE��!�BeC{��u�:]���|��Zqj2��%Z'K=ʐ�.z)�?PZb�TE�AeT���|u�`�WNN�mm��Q����~�E[t^���V
��6�~���<bW�GK^\����������3x�������fT X��Y�qy��o��QW�9$���fK��%�LTjHԤ�j/�6�����V>Fy�Y�j�����J����b~�<":���?Sd��<���"�cgY�3e���5��Gd����N�x�������R������t^
�o6�[����#f���2"��e�~߇o�h�7\t
�e��mieQ�B�[���.���*>z��v>�k��6vZl��z�,p���2�"aZ�8��7��~��_��x��L*vcO<ْ��:���k���(����#���`�nEuY�(Y[����Iw��'66q|<�|K�D�=��H�@������ZB�`T�"7�N�q��*�(�AX֢����"x����>�*��*2?���O~�.�/d������ ��K��D5� �f������q{h�K�&b�2Y����2��[�`���
���|b��5�,o~��yv�X�l�u����9y[�(��,���F��&��|�����8��O+����Id������ai���L@��͗4��f5�>.�7q��f��A�أ�8g��	�+�� ����7=#��Nr���aȫ�e%���㕧Ɖ�xތ�h�5b`�/"+0��kug)��T�&A:�\K@���F�UN�IZq#mB0\�8�ֲ�]<���S����j��N�������>M��*FtY�P� B �5㥉�%�T;4R���o������������n(�T ���v���BN^����^��¤"��7g�!��g[=�o�ĤV��؆o	ԽK�"˺J�-���Y����p������n/ߊ,A�M9�۳����������e#��R����il�;0����qIdä��ؘ�t���$�q��<��@,ׂRጊ�G�W��jMW�˞O��	��+"4)�C,Ds�/�����;H�{�P�ݸ�*���.�q�����*{S/��o_�+�G:r|�8ο^����٢���+)��"���$2�]��@AI�3.��~{�5�����a8Sl��*n��o�5Q�v����i��yW��hJ�6�d~>Mt���W�����6V �� =F3bރ��^1�� �l�N��<�ނE0/W~˒K�����d�6j-E&�k fj.���z"�$4��|��_V������� <<��?
�Q�J������@�x�4�0�����Z���&&�\���F����rJY�G0V�Ju��6�J���)�׷��C�2�[5�*�v��<%�8vE�:���2�e�hV~	J�M�� ;Fє���@��\&����;gc�{�T?�*֝G
qw�~�r]�����D�.4XF�!iӍ*"ݡ����qg� =*eG��η��K~HSͪ�ТV�]	��h�����\�h�W�����7
�c����Μ�>ܓ��ao�)d�P痗�"G��r�������#������HPj�c9p}� &T+�V7�\��/ah��Zu]>E~P��?B����9p�Ҟ�]�px���&�`��p��%^��&+Ήw��LVB���;-��_i����@���!6o�^7K���Z_��
��"'�d,����z��Y\�g�����$a�������X*SEY�nÙ6���ގpK���Y�6w_�Tv�>�F)�+��a�A�[��8�g�M���ܬ@���Y0��K�Vw��G�� ��$��șbRP�*��Lr3F�v'no�g�e�?JOf~�Et��M+u�K�XU� n"�x� m��p 2�����J@�I�3�7��!�P=IK��;+���w"�>�z��ϵE~E��󲲭�0�6�_�|�ŕ1�I�ifP8`&&��4C�=�3��s���H���Ϣ�^�Q`�����ȡU�(�!�����0uB�����{��������GEF�쪡
�׬'��/�5��O�����)�����!?��p5G��q����7�D`WW�tu��}s����=]+����&�ь�;����7Jڂ�1S'���v�'aĔ��h����5�Y��£̚��Y&&'vn������;K��r�]�*���|4*��E���8r'�$�/�ڡ
۟�ft����/�����A#F�/_=�����b�,��9���͙�EElA#�d�l�?XH�$U��W,��`���o=�i�l)/�f2�D_�s��7�������L/gX{a�%75����x����㻂��YŗL%K=�T�7��i���F�$q��t/��&*~$�/���7+���kH�pz�hL��}JI3.�]�¦��ϵu�6�?��"-]��gF!�T"%���CG����Ɵ�ȅ���F�zx~g��0�u"{S���'�`�*�kx(B�S��Ri�gG�/�&��_��Y^��m�N��4Q�V�*��z!�34sۑ�A��P��6��j�#���u�o[�T�u��cԪ��M�)��Ur�� �1���~03't��{���Ql(FJ�Q�y�cn�fw��wo9���j=apy�D8��:�{U� ��m��Z��|H�|.�����<������h����6��G�㨒}�.�Q!D�hMoف�%�H1x��@�����>�	�5)��=�.b���c�P�^0��{�-o)�z�|�V�e��B
�)N�7g�p�Q�T�aݮ'HR�t<��Nh���-�Ʀ�A!:�X���v���֚ZH7����I��`��_�-��Y�ȸ�A��#M�he�-B�D����:"S<?ۺ�]k|�2A��z�ل!�tf��q�/�䱹R�8�a����v�#ڄ����c��˾��������{��8L��i�֪��*	.]�ศ�ʓ�6>[��ܰ�ƻ�7.���JNN�r��-�!G	0B��������E��6��B�đ�,j���l� ��E�Q�����|�R����$ �Y�x&a}䚟4�j�^��>�m�?�U��	�n��ɉ4�u4��>��q����W=����w�h%���^0!�\G��p�|�9�.�X=�ǫ^�`dj�8�<�`^&t#�7ҽ�N����VI]=+zY��w�0 #�,f�0�T"f�fn��i����k���@c]� �b�Qk����r�?Gy!vٍ'\��#�H9�Y��ѡ%sٶjb��51�?$IJ��E���S���"dL�#�����5`*�=+0zc���s��ף>TN�7����?�@@j$|�+΢����*��ڸT�;��G�ȑ�1���~�s�8g�����1E�b_���!)��`z�JG����t*a{�e4"q�'<�?蘲�ɿ��k$C�w��i�	���-���	�#�I8/q��9��C����uh�	޿�E\�*'�q	���k�1�&��^3�%Ύ�`��g�n���,�X�(��Bc����ߡ�f��)��%QC{m�7�u��4΍�Q	 �ݝ^�&�.����'3nұk��#'����#�� �-xSQP�����CԹ�hb �����7J��Y
��i}����gN�;�6�g=��yHj���=w,U�f���Jb��Fm�|�H��ڀt^��Auy�J�����_=W��t7�-��/������d\ԃ�#M����|b�gF*��՗��{��VU!�~}�fIj����%&�%��C�<�S�kPbˎ�2��޿�'��,<��,����HpygG �}9��Z"���ED���baд,8�@l ��(�7����A"3�(*T���f{�J�+�*�!@����؍��������qdm��ȓB|/��>�/�b�z1_�+���|�Q���v�c��0Z�Lؤ�H��OMF|��j���ܦ���ЊK�	nj�P��?�r��
�H�Epv��y������1��	g@q�I�/|�X��>�3������ӎL,6��T���"�Q�,�._ݣ�XY6���@+��Q�g�Wt(�+��8�QI��ފ7U_k)J����fݭ��Ć��q�f�����F5�:	���������d�Y�)����B��1���uV��t]'��'�\C�Y�]26�!�͙DP�ޜP�$�J��۫�nplǽ�Q��tjk���$
_�9C3�Z�ˑo�,���RG�M�����*�A��c�g�A��%;��I���Wk^��K�OV*(h�T��e�?���@�o�����H�hi�Z�my/�V��m���](���iH����7���6@��� ]����Ipa��ou��"1ċ���Cmu�K��:�u�B�Q� @�b|D&P<����~�q~���"t\XG�f9�ӱ�O������=���ɨ9�F)DW�0�eͿr`�w�jVl���@��7=��V|�����Hw�B�/�{ e��zE���sf����j�crY'�v���U��>��6#�|�.�w|BI{�9P	c��0������]�]���˸n��>%_P��"��7�	���V"2/5��*���4��P%9a׮nb����쾃\>^�32�����F���݄���V�'�<FfsY�!�n�vՎ�Q�h�I(�L��-1��x��p��#��>�i>U��O2��w���v�|�Vs��X�u���η���O�ǹ7c�S��X�Xp�"� 2�p���1��-�R�)\���*���=��kԐH��%���u��ڙ�TX3?���t &B<��A����)�����l���W;��_�&Y|m"���J�&e>d^�����=}kR>v��/>�`1��B�6̄�ք��c�|H��8!L{����/�駤�hC/6�tӫ��<���y5o�̐�4m^*'S�;��Cw����z�Ҡ��4��!,��z���� ة����$*l��$!�%�O�<�I�#F;~��a�N=��!��T�捠/◟�.�~]��ɗ�0�����Q'�>Ѳ�gJ$[`ofmx�^cݯR�ce�*[��{�4�T/��8��pm�;����������tS_+��SlܢN�f��x�X�\緊z^E��y�M�{@vD���: |�=���o��a��VG)�4�xӷ������b�/�#`�AR��Ě�g�5�t @ X�#�V�3�QR��N7�AEtM�v��תs�Sa>���%+HL��g,x���1�	�9��Q~�+U�C)��W�s�*�QR��G9�f���s�}͒Z��^Yy��:y6�յ���`Wk��<Z�)�VE0��y�������*r	%@x9��-����bNA(Fp..d��,tX�6~�w��+'���x�u�.n���W�̄8�5�m)���M�E�&>��Z֣�~�ic�k>Q�z�,tE��̢w�.��0"��iQ(�O�6��B�0�/u����������:��h���O��4;�M'����y6
^�I����w�d�rf�`�=#�x�/Iw�3f�l/�h+w��*���[��'�ca�%(��T^0��U�V���;�IR�
,������\��.%.��偤���|���%�������+�7-bkv��<�;�9�k������R��DO[�~ڔU� p��Y������k�$�B\7�X��4�������k�/IQk�5"�W\���nPb5�����>���wU�z��aR��&Ȧ��('(\��w@'��[��tA$"ӂ��}� �y��Li~6*( _:p�̕ڍn\jz�9�.�gj4�3�̈^�����ψ��6Š�ZM~�ʤw�]3�*~�_o��T5�8��<Ӑ���r�����X|J�%�e}H��D1As1�i�%C�T�C�1�^� "AFSqb�����Ã��m:=w@q��D����k�.�D�?�3N��Ҋ�]�O�P�������9y��7����Ȼ�]��igǍh9o��WMZO�<K2����$��zj��G�b6W�.i�sƔ�N�ϯ���U68 <p������Z-S�	�����w�Pp�����ޑ��<��k�l���Zn[y��v~YW�>�ȧ�Kbũ�۟�E������e<�$��g�sŭv#͉{iqbW���V}B%��u:S�?�)�H�n_�a)\D#����,k��θp��W����s� ~�(�]~DJ��E�a�QO'��fx}�Z��|�j,�@�-d�sO��X7�!�&�%�ok�v�c�����$L��r����M��9��%
�z��݃�A�Yj�]T�>�m�[��æ��Ej�v�����s$F���{��[��E����l^e���mE�8��+/�Ro{�ݹ>C���C�]�9D�jni��d�hU6|��ۥ�l� &�i���Ho��?���'!%"��IX����䤽���(�h`�-0!�e������4��/2�{�v��7�u�����%���h��<�K�^��ó�� �\*�w0����o��M�޶�5Z���ܚ׈}ԝ����'��#T3:wD�r6��p��%0��]�MW�5���`���qc�L%�x������l@��IhM ��C>�A��"C?�+��W؜����X|�Fz0"-qP\u��&&=@E�H�!(�0����]��8��F�#ɡ.���M]�D<N� ��e�G�(9㲒G$�+u�ۡ���J��S3�U��!٩�<޽ #�Mh��w��u�IҀ���G��C�P*���e]R�dC��|m��&�O5=UˁI�����{ꓙY5�~K���<,&�O�S�P��i�f�ā����P$xOa�za� g�L}܌9���/��bErڈ�s�'��Q�S񎀽H��b6��g�,w�.*�Kwq����U�O�T�%�J�/ME�$M|p��X� ����-�V�T�����{�W4�_���Vm��2�x�;�j��/�1�+��k)���ȐuZ�ȿ��t\i�tӨD����nI����$���r�ْ'E�c�Ք��{V�W����F���aXj���+�ń���k贵E+�����J�U�6H�(�"��ӿc��Z�����|��F�(�9������B��̊��ψO.t ��ײ�������$p�˭�������Isbd݀3�]�zs=�@~�4��]�N�u��
�%�>�_ǡB�V�=��Ս�t�^��l�H@��;"H`$X�~�cw��+3�:��s�V4+��@�!T�zם��9���������="\����`�4�q�����rȟ��g-Fy�,~R?����Z���*�*8=]��1Ѓ-�*ׇ^[��m`&l]]jz��� ^.��N2�뜃�e�1��I]���	��2���d�������nJ#�sPwN�r
���#,�6�������o���DFI������q$iM-P�S���G�w^uG`%MXx�%QX�?�W*��9�N�rt����/��L���9<q��`r!����G�\�m����O�.�g�f���.V �IR|���'d~4q4a	�h� _������YIDBF�����]j�«�!Sǐ*b��{c���*��Y@��V����}�:�8�N�5��;U��fO7ϋa�V�bȏ%4W�s5zUΗT�����qɁ�e� ��	�X�*�Ye�$H����ȟ)�pB�AyA4���D�-���ɉ޻�X��K<�}�6�5s�o	Dv����]�Qm<Tyv>���ٿ\W,���A�g�����y"�>��'v�xGc�I��'#�&0r��������kJ����NO�2ڛmX��D��)$�k3�p�. ؇Y6g	!�����A�Vnޖ8�}RsD�Kم��D^�q����-i;ȤI���'�����.Y���J�t<%��d��b%�D�&7�d��[�lVx�@�k+CA��q�@���y]�fc�3'x���DF~��u=���#835��wyP8T��U3ް)��ӯrPղ�!�E7�pN�,\������g n�<��Y]�c��OZ��T&���ߟ_�Pq�-U|�����)E>��-}́�?F�?��Fn%+�����<N�s  �M@ �(�|c)\��l�6�S�K��=G����~~;���h�\TQ����X��	ͣ�<EW%�#� ���-�;D�)AXӯ��5�qb��zjn�!�..� q6P+W0G; !�������#R��)��f�
X
���t���������ݛN��c}�j�Z��O��}���l"��8�A�F��h?xű���̚|�d�J8�(��a_>���/q^۲s�]K��(N�9X}X{�䁭0�I�t/�F��q�\�!<e
Ո)��à�q|UsT:6��O�w�i��La}z�C=(�?�K���-T^�t�Z�K�*���<�A�_�A��1�!��ݝ7ۡ��r�9�1��D F:V��T�Sw�m�*�GF����`� 1�vf"�p)M�y��b�QhN� [h��f�Ur��6g	x�T�ײYZ�w�ǲ���W@`|n1u0N�s��Lrs{?�PP4-r���C�X��wF�3# &J��I�{Y7r
�z��+q�Ҧ��;9_�iG\} �g^&5���(H��[�%�s���-5$�R3�k� u��u���Ɋ\'�8͜����~��{aD������_с ��b�G�v��|q��u��x�t��&nS��l)Fg�E�1�ܭᬘ+�[ؾ�`��;�R{娥}��L��˦�pa��$�ݨ��<���&�o���5�rƨ�ְp[��߇պm��N?9��n���惶E�ᠽ_�"����T,MN:��?0�tP7�E�:�b�װ)R��ވ򓵗E�<��6Ė
��O3�C�|R��tI>���l�	���u*ⶸ�gRw���i�p�:�'�����"�K��zBK�\Qa�&��hB�;#�٘J���?ry��J�}�1pm�\�0��B�*)�b^�$_3��o��̩��-�/3�Z�ǝo�z�p+4}�IXRZF�Y�����<Ђ��G��Q/�*"Fh�<�(>�tƭӚ�Ed�.t�}��8��߄v ~`��+?��*���Y6�i�7:�������T�E��:о`$�'�*p`4�� #����'�Čo�p\�d�O�����B�5 )�����Ko��Þܰ����0p�tK9*��`Ү�s���U��l��\y��ݡ%�d��b_�$#����S���ʙ�_�=�HUe�i,y'� �Cw�DL�Z`�j�,|��C�\��9]#G�	@ �x�a��A������ϥ09�g����q�������|pv~��H8�W��]������8�n�N�GR'H4�����Sl�uG�K��4�?f1`���F`a�F�t%�:�/���n���
"]h�T���¤06�)k����o�/"<��#A�gHJQ��3><�c��^k�+}�`�<��]�fO��B`����C��_@�C�*�Ϝ�g��r��^��	�oe�d@�k�(TN��TT��+m85e!���3�Jg��K����)��-��sŃ�F�E;:��qQ9,P�r�i�WӖ�4�Td�?h���c�6�r	1�U���a�j�+���˕Dq@X}k�㘫�P=+p�ޙ_IyӟP�Z*�z�u��B��������pN�������~��p+~��X���y��a�r��W|�\0[�Xoj}�#��7[��/7D��4�(�$øt��.��d��AF�g���ڞ���&��4�%��Zq(3+wS۱1�hv�7��P�[.2�����ʁ�y�PvHsƹ�x��3���_����	�p��ܾ���x� ��tA�=��3��O<��]Ȏd,�������^�(w�9�V�n�kȱ%
N�X?��'K�M��+��5�$�HTx(T���a:>�ɑv������@��H��0���N�Ø�x��0�N%YM��8T*Y��F8��Tcs��"�<*;;��ϥ����P痏D\��?|�8�	�u�B�]T������n����On��f�i��Wx@����7�
B����8ңZ������â�����Xb���U5�df�o�~ȲہAjHi%�l�nů��M��lۋ�q��./3�x[��lGw�L�!s�>B����.�3B�ތ���h�$����W��P�x.�	��|�C`�N�}m!E7!���&��/�É��?y�}�4���Zn\a�
�P�}Ύ��3��g�"6+H��(Ҩ���&�4)V��g��~���Z w���,	q������͵��97E/��xR;��8�{m�75\�&�b�0�!G��zj֤����5�.2�������nWzB�ԑ1���2��+d~������Iņ�%#�f9a�\��H�(��3J.�pGjsT���em!���Mf˅�+V�'����,U?g.�/�^i��Ƈr��씼ńXc��j�b�y����9d?����Ok��ĪxUy_�m�g��C�F���N�w�p6%I%gS����.Q�6y�R��dꚒ)���)#���:�������tr��� ��U���ʫ���|��&�#�RF���e���$�/�8���.��b�l�BpR����r�	-�㮨G��Bt�"����.�����6X54K���@�Oj�P,��H��������B��d�R�Y�~�&�4t���(���t�LT�=D%�8ZWeMo�ѱ\*�	E����31��㷴��@ �k'��s���Wsͮ�ڒN�rޑ�*�mVl����A���0��VHV�$u��Ӏ��	��i$��Ȉªcn��E/��v����a�X��r��>/ws�\Y[;�ɳ+	|φ����6i�:Z���eR��S�fq��v}#�:�v]g�V���q���f_jFM<9�L�׻�F�S��;�Ɇ�@�J�(@���߽��LMg$ �]�G�T6]@��F��1<$-�R|[�.�S��#OUä���F�����*� �����������A��6����Ds̱QF~4�*��a����S\4^_eӗkib0� �M�>������0�إ���jM]V����BS�?�Q\n�P�M���\��l%Uf��[݃V����MV �ݔ4��]��l�YaQ+w�B��4���Lضz������X7ㆫC��+<kR�H���X�q��;H��8��z����l?=�r�����o�p����R,C�Og�U�� J�k�O�f$�t}���R$��v�I�h��µ����}�28?w�\�sm��L�&F��nS�@*�f����/�=��y�g%�;�6;u�1�Y��,ʚJ��X?����[p-6�L;�Ch�?��:p�o-���Q�SyL~��Ŷ�d7��`�xf��G��������͒��>�d������GR{1Ty�R��8L��r�������I\�y�F]o�
ʃ�8[7�4R��#8~g�n/�<���K
�(��?e�sJƴi�O��j� �>���գ4��J��¦��3f�t��9�" Rѷ�X2��&���g���o{]0��|�Z�K؉�<[��A ��2���������v�O~�GF8m@r+k>�G�7�ۘI{D��,z�V�4H�q'���մ6�H=�^�J�}���:���`d�����S]ք��ο�w΢"B���M�!��\��eF'�$3�.^��P+!YB�Rk�Ӭ d��e�e���5v8a�,���j�m�/ή�D�?;������0��aҬh�[����u���x�a�(��up^��cl���.��l�#�� ���������`���I�Y+iuJ�Ј���7��_����~M�G�l-"��LX��2W�����˦	5w�J>��ܸ�1(��t��_�U���)>6�t9���"07�}��=f�G�|�C�#�E� ze�I+뮡�т*�
���/ؠo����f�.r�I�@Q��^������vKZ�`�h���p�1�d�UnO~�'U��s%����C1��$MV���8�&��cũ����_�3����D�\I�9�}���o�!˜�������K�L�X�G��ό�F�b�*T(����g߇[���',�K��F�{�t(#@BK��#�Q��Z�ժ��\��n��>ǆ=��Y@$*�d,����^�˕�5i�Ț@��mb�]&Y4��&���Z~�߄|Б;n|l��\��T>�-�����g�)�V���2EY.�@�?>� ��xc~�"����`X>�r�}��r$U��JO�+B����y���=�i�]2�P�y��m��Ȭ�-��v�d��K���쟬��}��\BYd1�)�A��'����!�z��u�z��!�f�\���n����ٶ�vP/X's��#���J���c͌�����͓H�UO���q  ~��3V�5
c7V���	3�NK��8��~4�� �	_0aa���euۘ+�$����r%�5O��ǟ%�~��|�"i1�v�m�G3�D�K�{(���sܵEp��b<8� �#Ǹ��nσ�z#F���>HB��KB*�w���.���@+]jVVY/��qQ�N9��(n��iUR����kp��Z���-\������dQ^1�����	D��%��T-����KfxǦL�ďgS�۞[��`��M�>���cv_���if:�v#��'��u�&���:J7��&V}���>�(#)~VG0�Ɍ��G�ZO��̺(f������ �	�L�E�Ej ��'#�+VS�e���g	fk�۠L��c��$�谶Ҿ�]JO#���� ��r�W���۫�V>O�)��&1���K�	(
��m�8�T�����&Q( ��+׶� �U5l���ֆo� �������ۂ�L�J��G�69`gψ��S_K*�.	��k���ão�w�y1|�!Yr}Ǳ�ܜ8ן9-�;��C��#,)~G�.Y��o�K��*�]�E���������+�4��E���ϩ��jB����6M�P;C�&���P[��Ǐ�?��G>����|f)�qڃ�B�7{X���2�I��^)/ٱ'N�����x ���	zHd�	Fg��$�n�t�睅Zh�Q��2~��`V�u��?�И����q}UW}R����iÒTf����)b%Y:�>̯Q�#>~�Y��F�i;��\���E���tZV�EwM"~�0!�&/dbm��l�ͺ�cqر����ny2�
CC	��,I�����g��|��_&�i�C>H��&�DdV蜙|Fg)T��r��%}V��=+����T��܎(����H�!��9�/�--�<�b�S�נ)9�н�d��"D!���c��lc �=H7�[Zr��pA�.h�{����jL3�����s���f�*��a�;D�@�H�(HcYS����s�uCW뉳�x�rv�@��Hb{�bNA�����ܓw7�Z8ޟg�Gp7э讵��!� ]m�^�h����J����m��ck��q�b����Pq7��6Q�kEV����4� *ĭ���"[�k�aI�\�=+�_�`l25}��6�Q	W�����o!��+sO:��(���^T\��)�Uc�dP��< �!:���:�l�L2'��?DF.l�>^���sUq�f�6���0ɏnQ�`EwC��oy����˽T4�;��� �A*53�Hu��"0-Mⷘ\k
�mB�΁�r(<)�$�t��7h�i��ԜHQ��+�[�E�{����z����+9�Ic��Q��6k68ΌViQ0�r{
+������[�9��+,!B�8�b2G�$��Ap��Kܤ����>���HJ:�. �0�ِo�2��g0�s��᳿�p��eI��s��k�䝠�/��C�5L.(UYc�����S��G�G�=�d�l��mv՝Ly&��sE�*�!�ƣ�On|�<s/�b�h;l=�+��a��`
G�l���&&��a�8D���> &4�a~���	vWZ���fyx'Nbx$��K�I(;3i�V�#���a�a���N+�D�
�9	���.�V����W�����(4N(=E�Ƣ�YG�{G����V����O}���sX�����Sn3���ﴴ�h͉5��'�l�W}������=�u�T��<PA������X�����c����Y�?~���T���tᄬ�)�f���
�)��=>#C��x���ĠN��{��%c����V*X2F�ʝzѫ8���ž������d��5�(���Ȗ�O-�wB���Q�!�Ў�Lʍ�F1,�����ȖA,��!,����u�R��
��0E���^$ğ2�֙�e�5���/����GN
|�|VH~v��Y���uڄ�vT�p�hs�߱1w��=k-�5�����;��`CW~�[����qwdc/_��e^3U%0��84�����"��x�Dl�YՆx0�!n#����^J9���i�f-%Ѹq���,k�c��&7�;�"R8*�.x��E�S��p&�%�&2�-�j���q���P�@�v߃?0�c!��XuL�e]wA�(��U(Y��v����ו���8��8Q[Q�@)��� ��⫼��9���1%k��k;w��<��f��Q��i8�xt0-V��Z^�2�� �a 
�� �o:U��R���~��PQl�L�s%���q,*�L���DT�����9�CΕFqoE� ��P�4��b	�yq.q:W0&�y��WȢ_>YH������7���5p,lul��
�i�r��ܒ'�Eedr'U~�z3&��*~�m�h,���"�����	�=5{)�u��!;�:�Ş�=�'��E�B�2�p*��sj�2���9���X]`x�Fz/�\�\1��Kl�Ji@B���I��B짥N9)i\�|uS#����E)�h�c�^��\,�@C[n�+����� A{����W}�.�qԩ�+�$�j�D@����a��ˉV��&�����w��h�#A=u�>�B�|uA����m�(5Q�;B� Z�����y�}T�^��!I��zh��t���)����P:��F��9���Vz:A���EB(��h�Om���*$1!���2ta>�� %�N�<��`�߮�@��7�p������� {5�1�'�\�j4���2��&[]k��cۋd��Yڧ�#�L�6lvSj���ѭy��b1��=���3?��aS�C�Tp0�^��@\�)��4��3�'P��r\ۧ�N}%���������!!v�H�G*Q��������l'-�y�I��Z�b�^1fm�5*zյ�ڦ�k���*��:� s�Y3��3B$�%��XF� lJ?ܜ�+HG�w�;�>��g�Laǈ*s��A�d��6�o�G�oR<��I�����^gV���<ՖNL5��s���7��(u�W���Zv/�<>6x��.��ܷ���.�d�6�\~ԏ%�o U����m[pI�@���٧�1aL�%!5�>d$Ӿ�^��|.k	���'c|������7����ġ�O����w��c�����T
��ڮ�B�j.�-S�&�E�F}�`�!�=�Ȁ��u�J_g����'���V;�0-�f���b!���ES���hhl�� ����V���6��^Vw���L��Xr"�ޢ
����ǯ�����QH�]�)z��Đ�.T�@_;���=>����ԫxL�l ��WIX϶�K�I\_t���7;㈪S�F�O�l�/��Mra����I�q�Qe�J�8�0���g�F 젘�>ߒ��);�q
]�;蜫3����
߅c�(�6శSou���q���Fg��&^�*�[E��P\	��?��|����I���a�k��g�"�٧��Yi��O=��|o��ܫ̚l�`���xy=Y�@>�������T:�P�� ���Z �0[�F�fCj1\n���r��qYI|Ȼ��qs\�Bl��P�!�?Q�>mN������Wbf,�H���(bf�]��p%��M�D�n�ج1��X�@�	�Lx�VpBS�)��
��q�dԟ�.���,w��F�� �L��[�%5fy�~.3����\At��Ó)>+r���Aa<�^݇=���@g���������f�0F����l����ݩU�n�B�_l IZ����:����^�����X"�|��D��杦gS�Y5�I�.���O�z�I��S��1m�z͕?5�(�*e�)�)�o��h��8�<Ci�b�F��fxR�1=2q�"g,�O�`!�زf=�޺�U�k&��;��,��Xh��&�[Ԇ�"���6i�	���Ms��"�<n��5w-j�$a y�����Y-
t�d^>~5gt=d�o�+��6�6�2VS�%��O����BZ[���0eȿ�+!�h�W;�&�8�E{�z�wQ�"E��=Z،���Rs�8��g��^B��3�Q®	b2�k��Yoi`(��Թ��<���(��0n�s�;����u6�z��ݜ��rA���z� ���0��Pv5��GT��[r�2����zMWL���p,�6��e=���KHv�w���l-z;����Y�4r�ݴ'Lgsc&��)���T|tx��M����,2.�����	�����&�!á���l�]���6��z��:�sW���9d�ڒH�8ndh��
M,t������靓����5�;�-/��KR�x�Vg�hbm��VK��ZXs� [��-Rqs�����b�=RV(I~}閒
~p<����9�`�����,�`��`�m���m���p�^8�� U�fuO��y䢮Hy��~,�
9���oaD�x{�����<�H���O�0�qoxWӥ��0��4�u���9�*`��պ�Ky�D��_�2���5�S�$������z�a�?���D�d���/��X"a9	۱�2�F+��
�?^I�gz�M�b�,�s;�o�bi�(z;9h�����s���+�?�+�p�Q�#-3�9�cX%���[�Í2+��aӄ'D8ta�LP�%z�Wߕ�'Ù��=�]΋B���Ҋ̷.f���)�� @��|*|z�k��]x��(~�� ���v�͉؏o�C�,�|�����'g�zh׀<�M�p�K��
�z �<��^,���y����R0��+�)gC�:��W��(��e���+a�h�nr�)n�5��W�2�
�R218�T������X}z����8��Oڭ��9Q�N�&3��vq�* }�:�؜�[��TdH+0��O�:3�u��DޤJ��6���X�2�J�{տ|�S��`�AL)a۬��=۾�v鱻� ���ZgnOm���ߢHl���Ǭ����k6v�D�_�o���<��]H֛n�`�0Q�X�Z��y��(yFR�����*���:p����ȝJ�!bYs9b�^x���d���	ڌ�
ՑҐ��9]48$�IC����J�(6FK���8�`�S8I(�.����2x�
�V�8�*�A�<����&��)1c%���EӮ�Jq�����+�G:��gփZ���0#B)�>��8u���%"���[��m��U��«�D�nb�m��e�D�l���� +��t���ڻ��k��Bz��2�����F�K�z=p��n7��R�Cȁڭ����w�c����:CO�,��z �YlK��v��যH���e��@)3�I�-�/v�$>��W��ӂ'���*���1�b�=�N��mztm��|�#���N�ER�	[�\�Rg��؏4Uo��ɶ҆♌+��}�;F&�?�w*���0쀌��P�}{-�G�?���\�m+�ӂ4A�[�Ui�Q[7��:�Y)��>*����Y�Ra��3HV�d������EM��*'a�|��V9h?��K�S�L,���x���/��ܬR�������Е��!���H�ǀ�A(�:^�N�:�"|��O33U�g�Tn����$�rR���h:�s�b<������=�5�Ja�/*O�����OoW�M~�"Pz�����7�����
5�?{�m#ݤ���^�al��|�B����H�D���l3�̘��b��}e>#,}et�2��mc��E�	I%��?���KOH�#P/B�wf)|mPC,}Ǚ,�'e�~7�-�$6ɿ/���k�A��¥^�C�C\ܸ�"|2�`T��v�u�IN�[�D�F��E�eb���!1������0ծm-/�\����j�,�\�1b??Z�y��(oy��+}�� </���'$�ai�3�Q��+�18����
�H�"@�^��[n�C��j7n����y�FGa��0������/�$5��÷���ȉ����3P���,J��F��~����l��c��p)���~��ߑ�g�N�2y��������p��n��8��]�G����F&���³����Ű�9``+t��lO�C����E��y���x���������p" �Z�mKBp���8X�����B�:4���NH�C��D��sb2w�w���!��}U�w�Ix'�����.=�8�U�G��е�CM���.T'q��#*��A�������(��v�^.��蚅ٗQ��b�Z�W?_��>�	�����m�4 ���L�y�~}�=v��LE�<I�����=~�!�&�Y��7��p��Y��7�׍ ɰHȯ+��$w�:t�=A���	f�܋RN�ׂ���֞ ����ھ���0�����TÁyCu��P�k�e�,��Vt]T��4A��������n����q�m�y�\\N�)��/g~�J�h<�5$ū��cS?6ǩA��#��<Q
�o|�繣�N=^~��Gˬ��0��fJ�*L�Ka7: 2цR\�+��K�� � ��M(��V�.��������T��<��r=�Q���TYog�	*��톢����(u"�Q��X!�p���jl'-�wxO"��R�Tϟ�f_d��re�')��J�vL�\, o�e�1�|_&�ZE�~�r$������W�Ղ
���5k�Ni��`	4���md����kR Xy|*�l �RA�lJ�c����L]�>h�[H9T��[�&U<�"�9=��JS����Y,.n��^C&��E�^B�*%�j�bJ��O*f�Q�8`f\Y��]Q�G�9��!o��ejp�v�&�Z��2GOJ�5�:��@4#вUx4�`g�'m+��{�%��o�A��i�ύ?grޠ9��Ǚ_t�(�n���b܌�.#0�d��Z��L��2`s�bt�a�-'����x�HHW�XZ�z�~�Z��-�R�W!�M ����Ξ�hg�X
�SP����dr^�b��I���xJ'rVk�GܾJ_5�ނ�b��b;�C���ǆ������S�	Sn��4Ω��T����]X 2|��PQ7������d(l~1����D�hCԷN�s
��Ċ� ��T��(g0�jDv��1`�9�z�S�¢�U3\E攜��4���v�k�n p$k�KC ���#Ѥ�{7�3�_�����;|����]�<x�m��`��W-��qi;�Q����}�0��Bh'���-�i���n�t���fWxJ�.,OMb�j��K-�nu!�],~��R/}/��0�#��:�l?V���:`����h�'g��i}���S������I%����@���N:�-.� я@ϒ:8�1��-�al�=����PTY4��&�P/��W����=�X��r�*>ʎL��K��:bz�l�m��s��m�
b]uB�'I��'���դ��)�G7HNh��@�2�xMݙ�n%[�qk��`�A��S/N�!k�n���c=��Vt���ׇ�H��3�%���⢥!�a�"E�~���Qܥab��C"Ʒ�L��HA)�'כ^-�aW�(�r���6G����c��mn��z�i�J:7M�S�U�p�w0��+n�g��Z��^:VUR'������揑UZ��)��Q�5��Y�a�d��Ar�����o���()J�T��%m�f�����Bo���>�4_㠀IWgwxsX�hO��U&QA!�9�dÕ�D�uϡ��V�����$�cX��~��o���r��5NAe̜c_��: ���v���|�� 9&Y�� �X��s�HO$R&�{"��\����kH��ɾ4����f��x���
!ێ$���*Il>y��)D����i��B���|TH��"�L }�ۙ �A"�-��g�[�ɦiﰂ�Ƽ��Z��i7�������q�����砏�/��y��k���0�ހ٦�@�V��*�<�S/,����}(5���ZQ8�|y�'���u�=Q�?���:�U��� b����������z #�Ѝ�d�5�祿�VeppÝa9�LMd��{&�� ��!l���<��X��Ր�4�,�ީmN�4�3���ב߾����Ů$A�13�$Zn����Z[b�x�/`�4�Ǔ]74�(ї�,Ll�9sr�ў���Id[A}ίZѭ91q{
]�p��9F�I�MI�������4����hH�=�;�Mbf���y��SC�r��b�![�7�Y��
�l[�u(WyS'	�N>��4u}��9VD��v�l�+�T�C�?rNן�� ��a8=�I6���~���=ԅ��14�$��ؙȶ�Z9Ib�6�Υ1�o�1=_]�ޚ|0�"�,�n�Yr�#~�WM!����+V�����,�.,�H���ppe(�b3�r]Ǚ��0~"�w�����!�\/�� L��b ��9�߁4q���QG�|ڔ�>��A����S�+�=n�q֯!�47~���o�b.��7Wȵ�}nmx��B���h��h*u������~@ŕ$	z��� 1PKp���S|���r�$=�0,h�� ��Y
�9���m��!|��;�N6�\���E�dܫ�T�!�Q*�h:bҚ�cJ���4�
AnۥΟ��g���m��(���v������`f��Q �w�!Qt
c�+tfTph2� � ����%'�i�0�:��˓�����Z��m�������E'@ ��F�NM�۹|�֨h�.Еawv�ު��eo�몥��>o~�W:pA�+_fQ������6kiʪ �H�G�Au ��i���Rv�dw�C89������,�Gc�a?�ޤ�~�.\�w7@W�r�g�P1��S��6���9�
W�M����2��9����o�DY�jF�T�����KU׏�D�]@�b��F1��
�`�q*${B;P���	Z� �S����т���gkٙ0G�w~�O-(�YhN}g�n<b�b�����"���1A�L�V�^���A��)ȹ�֞���>���^���;�<����q/��!��-�h�ɍC��ꕑs����z7o��Nd�	��Td�*�xO��Z�Z�����3IY:�§��ܨ��i�'1�;-�����iEבך�N����`�o=3i�'�iH逖�bl{to�Q����sڔ�W����T����:���~�X��&�/���+?��r�N[���{6Hb�n��h�=L,e�9tΰ��"w��x>�����~����cǞcK�ąX�i�,�%�N�߇�0��cxe'�f�oJ=�k��Lu�3���H9D�00�~.�/����T& ;"�1��e�\ר�P�/�Y⽑J��VZt,��SK-U�����y�)����*5�.��������n���7g�� �@A�8�L�IE�J_NG[�᪀_��0GQ.,�oW�!��5u��޽e=��=� �{Y������S�􌨵[ ��Z�--WBc�e��d���\sO�=.� �mH�
�?I ����Ȥ7=d��&�o7�K���
-T�PC�V�Hq��M4޻����Y	�zX��������� )���C�#A ��rCC�FL��geV*��'т�^�Lת��'@��jg��FD��N=+I:�/�HX���] ݂K��tQ���W��ޞ6�`̪Y�x&/i�t��}�"�p����(�(��pA���rh�?�����ͨ�,p�y�5�-��*������{�uX����>�4x&,@6n���zw�mz)E�U�E�$�,��x4~�$�d<�_��}����XLT�%�j��zE��ٸ{��Đ�����b2�~Z�ݗE=��;D���yN���k~��z
o������I�g{J�!{ c��<�}�`��O
����Q�R��U��}���&���0�\�c��A��r'�[ f�c��aɆ�!>F��=��dNU���]�I��
��H�ť���9�U�%��`�3V��*�ɲ\!�1)ә���AM�a��D��ľ�2�3�����%�E��	�`��u�^�S0���5�tD�$��n��|I��F\Ư)(��QD�Q�H�m:xf�B�9'�s0�����C�|�hlS�|S���#���z}���ꏋ��d��sV�V���ZN,�#��n��`"�M\��{-�Y1��*�7�Q�ߥ]�V��D��^HL��&^�;P7���Cr���U%N�)��޶�˙<�V�.�-���k��Wv`�n��m�_��#A��b���<O3Ҳ�+ˑ��k\Q���[�28���9���D�ε�}���S�(�@��砫e�%g�_�����*�6P��R�.��b��D�����L��K�c�e�pde.�J�o��\� �9��Vˍ��`�?�p?��I!���-�ߴ	4��R�N�U���T���,]�>�\%�R���R��NF��6r
�޵��WS{G�P���dt�/jBmP.���*Gy03�$nkmA�^,�Q��D}��$���nYD�
T�w��1j����G8�c�T�5�{��1�_N��k����M_��S��æ]_�z8ֲ��ۂ���9WJ�0V��Q��kot�u8�-^���
�-9�vB�Q͂�MH��00����*�"6pw���w�fT[�:)���Q:h��!� ����L���&�.�����7)`�v�h�0�B6�ܺojs�C*
�RI�`v�ѡ��0���~��`�b?+����"��ъq(�7#G������@'&R��</q�j�@�g���RӰz� jI��;D9�?*�|��n�}ZXa���!M���2P�j �0N�xH	0\Fz
� ߈��?�<�7���q����ڽ����<��oSBF̗+����R�����ۙ�.�}�@���ᐚ�6�;�e��*���o�9���;��,�9�1Ь.2ʷ3�4����� a��?�(����TT�c�<���C�Ϡ��;��2V`��|�/`��n�j㉡zQj)c�l���O�!w��h�Fc?�9|qw��,���]�=��9�K���E�L�B)���FD��"|����	��1)���Ȯ�s�eY�R����
�X���y��Cj$���NE:Iw�a�X�u���^�NsN}�t�t��&��җ����a��fi={�V��ކ<�l4�23OPa���#�5�yŭ�o����w��\�p��F�3�3���:��<l!3�9�!�Um9��G�iv�=o�\?jZ�l��i%'<kq-�O�M���Yo��p+-eQ'hӎ��%" u�}~�2��q�K�X�"��%�w '?_��L�.��������T���Lv�������⦬eK�9��9?&
������~�!Va2������Ni{�,%w8f��l�s��7�c���>����}B~���A�_�P��i���)�BV���6@���m��������g�߬��-��͛��x?L&*�r��+w:M���mt��QA7�q�������q��-0���%��'vɢ���&??[�����¢J��\���G|���""��yH0>�����G3�>�mt������>�"�:��Pjj^39�_���W�������G7��A��`cv���9'?�SezA��l�6�0����I�+RR���v��?}铠�1l�4�BG�@۵�Y����j�����7���J�/� Gm�Y�����v�K?�ĕ<��Z���6����~�n��p��`�-�<�j�:��2 �^k�5v_�2�O@)�����k��ٳ��*��9�iAv�o���>����^HU!�Vh墕K�%4[��GQ�(�?KBK/���!��7N;[�{�o�*��oK�Č~�c�(A��m�BWZ<0Ha�Z>f꥖v�|ˇ�&ѫ����[Y�`�~ ?d�g���rʑV,�^��X�JUPgW����U�;���)\��c��ɞ��F� F���a�}sV�g0P�x+у��3EN�Mm��Yij���&ο�r��0+��D�+H�o~�,�>� �����!��{t?���;��oa�׃�;ޛ�n�g�K^���r��״jAGݞ�[y�݀9�����F�����2t�/(��I>����Cb�E�)�DD�ﹺN��r�����E��!X#I��Z�� oU��"d�t���!��|�ȫzOq�^;
>aٱ�eC(ti� �'m����u����<��'K�͑|�$�<�; ����a�]�:2c���J�o�&�}u`N� ���}Gf47�ۉc?Ӈ.X��˴
ӧ<?�Gǔps�O�x�����Ã�r=��h)�����,>�r�Ff4o�X	��1���H�ȯ�x��[	�����5Y8��=��i��m���G�ӕà�O�i��k"3&!0�l�aF^�d�6���*�i�md#���%r���h* 	7ǒ�M�P$�Y,�Ő��TL�8�y�`����m^�^���`e�繨a�!l�k+фtm�[0x"�{�Ms�8կ�0gb�mi��Z��E\����\�M�y� �1�L�G]�G>ٲ^�C��4�f�-�m����LqϽ&��s
� i^�.W���F"#�A��3%���]C�/g��تi�sRH��1�0I�����=$����(;;k�3Vs�B'��a��9^�������w�����ɔH�y�7���2VBܻ���o�)kH	�/w+�ԎT������/��b 'i��UP=����0O$��6}���K;�$�TtX�?E|ԚG�H
e6�nn&��8Կf��6Fy��O`�g�;��0hz���1�"��)9�Wi��GZ�N�U9s� >�J~ٍ.��}J�>f�����."�8�"J��#��x_���(2Q��4��R�pvm$��� 1�����0���-w2��v���>��p_�]N<��'��2��L'(�0���
$[������$��'��f^��˹w�Gh,0 �t�i&���H4ݔ\HY�4������KPh�.���+".��|8d�8J�r��	�#F��{�L -��<�^�#W6���YL�A��p� ��\	MJЄ��\5(�Q��A"��}}�7џ���B�(]?�3�v���X�:Ȅ�m�i�&��q�ɘk<3U����L"�����b��r�h�v��va�j ������&�e�g�I2�2֟-c	�X�'d�2A&L8l:�V�D&I�o��f��nnEB=�s�������XL�}�������3q|N
4!��)"��U��@�g�A����a�/�Y�H�[��w�p
0��Xx2A���ٙ��Yi���g�e����[�m[Ip��,���TlÅB��t�Y��(������5.��w�Âz�S�3�w��� F�{j�8�j3Sx��Mq2狵G&_KU��wM���ͣ���ć_)�l3�A:�ho�;%�kg�h���T�/fP���,ŏa?��9G=�1�c2&ϤE��_j7g4P#?w�Ń� ��Ӧ5��ԦGl����f��j���L��K���93�7�qC`G��2,M���n���R��>�;��e�������<ym��M��.'w��.1��i
��B��}ԛ�v���U8�������L%����刦��m�\2��U����+�.��ʧ��H�NK�hI��Ծ)prD5�*:�sN���~�|�6vEysy��J�����m�-�MCK�}�L?��\c�֢V�7�cX_�A��-�.�3�F:ڌ�୽�U�ʊ�3L��4�q�b��N�0�	�t�f�w�NQj�"�� ��������Y{#�U��ZO��'@���d˄�e�m�[�Z��kO��J���T��j���H�*+��T��e"-�e����`Y`�9��@�n���>�h�Ձ�\��/ɹ�1����BƁH��Z�Gx���?��Г��7)�"P�� �5 ��b���<��Qim�	�ӥ�9�3U��s����U�Ӂ!г,K�쥤��QS���t*S�f��ط�;-��|���= ���Ne�F�\�������(�T�<V({%���5�\PD�w���X�y�c߬S��)4����Z���{�/&4�'��,K��N��^5���K.GZ7�JOg��Z�h+�o��l��f���d�qN��M��&b�`HK}��5k���>z=�R������f�珽,�!{xDV���c3{
�[���ʋ��As����bA��HWy^�п�]bo|i}����Rm�"�(�ÛQ��{����3F˺�u�Gu��еXԆ���E[�=�j��k�n2���>~x�yq��D�|
��+����7�A ,-�o�=HV��6mpO��ۯ��8C��5 �_�6�H�ވX��bnʹ�֯N����IDф��5�G{��Dm�E��A�^��>D��b�z�Q���$�o\�R]D9��Y$��eG �;�7Q��e�-�h�53��ז#{�)t���q}�E�Q������ �a3Z��A&Z�/��
��i����i(PV�1e�lW�J]i|J(I,�(��~h�A����p��T:�����%-3�^�s-LdM�Y��Ѷ�`��zf[� �}�^1�z=�mH����@�Q ����3Jཛྷ���7�����_�C܀JP@��O��I��:&�P����'�]�Z��J'���P�f�� �V#�mcdZ�Qw��)u`��jp�T����������q�b�K������`�}���%����FZte>��C"�.RS�D��|�]�Q6�g��l�p����|D��x����d~����&w��9p<�(�*���0�]�d��H�t����!V�ҪT�:��?2d�`$G�E�)9B�8LV�H�c#���US��T�wk��M�8V�~�����du�s�޳�՛'2�+�i���a��q�/խE�;���<9>M�����3�� L����0�?w�$�Ա��*}���	�L�R�QIע�v�@�:�v��v5M>�:��D�������f�w_|b�W�©mbXc+HNk�6�%_ty;�2��x��3�v�����W
�r��/+V*�D۫�Lm]+���Y�s�z1���L�0]u���F#=L[�h����\��.���GO��N�[�5�����|��	S0�[��(o�'�q�
���:J݉��{t'��ׄ�G���qh�Sn�?4�yH�x�q��q��h�v�1Q��#��@�D����e����*��c+B'T�%T~b/7<��v��	�zG�%'�	xn��<�wx��a����GԱW�E��ɯ�r�5�������s)��8��Ml nD�*ݐrU0���pAFu+6��q��A)n�EN+x�%���n�A���0XiI��P5#w�» ,��{� Y,�K'���R��=9ʹ��M��V
{p$ܑ��%�y�^���|In��������ևiY��S��X��Н��*��u��
ڏ25~Dtäڀ>��Ce*XȈ����S�~xY1�sW�;&��G��v_æ��t��'E�R�b>�5�tN���i�,`���:�(�N�/�A��#����878���5EО���G�ʤ�|��Lݽ9]/!��H(%��
t=�ٝ_'@��<6�ɵo���w��9wW�`ظ�J����H�7��O ˗X�Fj��a�c�)�|¡�����?p�8V�~L�qa�7�܃��b!��8��V}H8��$�����,��bT��Q�q�L��?I>X�M��78�b`e'm�!=�_M(��@Y��З,r�8�jC5�pS|��.�*(@����+�LmƬ+^�����*\��o�f(,�Hrv� �&�}�a���tё��a�L������XC~['%�o>�f�7�a#�ݎP=�2_7�{)I��݊�m���<�(���TZ���4TJ8v�`��wG8q��ﱭosO���i���'g�öၞ�Z$���48��U�0�wK��F��U��=�*,���yK�~��Ŋ�)��J�k~��ġ��Ц�ڡ��˘��&h,$k��%�퇋.꽒�c����iA��D�3���,����;�,�P�[���c�<�h+�� U�L�E���a�W�[��z��7��L�a�2q4��<�F����Y7�f+�j����<��S�c 4��V���kD��>~��l^��8�䙀���:_�����pr��z�q35�����s�kw�Qo���*�:�W~X�ܥ�\&R�^*E�}���T=��@n��V$R�4e�l�V����%�puqR-���1^>� �W�)fS�Ux;�L�v����3�bЫ;Vf�|S�}��	�m�����o7C��%�ug��@�K�:���juX���$S�aȋ���wN��a`!>1n.���f�f�V��_Ifq!O;�o�..g_���25I�ۤ���4�t�1C���D����]�o��	M�6W�J������Qwc��G3I�Q�3W�
#G�H������O^yW'F��k\��"I�/���ޡ�5�_���s���8b�\mF�l�]-m��;����{���bjـ�IO�U�,}��2&��H��ڕ�͓����84��
�j[��3���p(�D���XKZ�> �aăz����y2�I�@?���j*&����~��|�U������D�R�8����_�%H�r�B�Ϡe0!��a�7�+��!w�Ļ����*'H�G���$ra�77P��6��愊���R�Q���Tx����
+Ŕ��)J���p͞'�F�\_f�0�h���i�O�=�@��S�zwv:��C	V�!�gOx���Wg��'�>�P��ID�I�pl5K�#C��]�v~�%�����.�ks�&nP��7� Y~�G5ʨ��I��E��Fg��/8%�⁾{��J�:k2�}���)���ȷ��~~x �o�Q
'3{��C�9e���]�{�`�	�n�3VI�����޺����K:���÷]]�����]r��6�Z�W��/>�!ܝS�+뀦?�`M?��I�X	�+�)k������cq2xW2�
I>�ު9�����jY3<�p58����}���u����Q&1i��o�ۥ�S� �1Xǝ
>W}�����ok�6�]����6���=*_�7�*	ӕ�YFE�MEB�1�,�������gC�<i�joY=�1���t��o/FLO)��T~��7�"��C�+���%���1�� C.�l�O�k�R��"�E����s��/�p"��^��C|�Z�㔤d�A[�ʡ����� U���i��5Iw�Mo���Z:�o>[�5- "zɥWj�m�[]��Ό�9�<�;��=�Ͽ�j�����0˴�f��U$��(�9X9��B��oAxj�@�n��i� NM&G���5J5�^��n{{ېYso�,}�;�^嬛Ԝ��A7��{�A��פֿF~P&���JF���V��3
�5�s?!gE�CE��MO���k�$!c\���Ļ�Z�]D+��.�W����s[�<{��z��{B���Ș�ʰ����[�Z&��6SI����>�������Qz{���M�!���оu��uQ�]�!�X��6I�&4��]��\��
1�������Ğ��0-�k�7]�郎��EV	{��gˡ��:�0M����V'k*ʦ*�����x�qЧf"k��@��q��þA�)� �u�0�x����j;�`�]�C!e�o)��6��w�E�����Er��1���d�,���ީߩ<�TW�#���H#��v��%eB�V�a���܀�pZ7|�_��O�U�;����'z/�O�g�k���Y�]��lƠv*��%Q_�=�y��"t�\�m�_W�s�b��[���NK^4|^1�c���_��s��.̡��ԭ�/��8`�:���fʸ/�XXtZ�`�qg0{�B�'�ڡ�eoHq�x~�L`�F}>���N�0���~ޑ��b7�b�d{���(�ii�g����Я�Oa��3�d�?�N~D
�`�	�6�wD3ӿ���]�{@2�H�����;DX2�!bi��@��l�>��&*C4���B]�\b?\�9�Y;(w�~\�SW�LJh�Ғ0�)�i*�S5�.���Ի�������1�)�2��è�͘��V_�6r�˘�?��~�2Tf��R�Λ�'X�8�&(�6����u����Kp�<qu�v)�4ٍ���o��@O�4ǁ���Z�9��T۾1���0�8���Y�]�Y�[Ht�b�R�
@��:���|-�#�,N-1�&��v����;؀�(���BonƆi��+q��W�Yw���v�2'��DV�^�i5=�28I��Q���IfJ�oVN��Đk_ ��?��A�]N�e
p�J��`�>�	t1H`R��.x�6�?麑��t��uz����}���)��m�A�����m����E���`�9$N�U�g9=���`܇&ۗJ }�퐠sZ>��
OO|4v��J-x����.�I
�X3�c=%�9�n6~ |n�c!�u�~oI��4E1�U��)��mX
��'�W�����jm�qc�n��^�n��@1DJ~i\�����+�yqt�6_b7��;��ځ�T�[��#�	Ac���$�-�na���N�����x���|�n����ʾ�ښ%|XX
�o�Nk���P������)ut9� >�D�`�PFdҔY2��l�t"h�R�y�>f�&-�����b}�|�:S�G�5�c��Ȩ�D�jm}K����4�{��I�ؖW�,�*�5����2э�� N~������i�F��G�V��/B�:ON���D�!�_GZ�_d���R��C��Ɖ�[j��(�h�E�{CL�cF:�]Zt�w��=;	0"i��.��M��'!���	WA��X�~i�i�$�"�#�)]���}B6�J�C����j�͏8^�ִn$�z����qs%���uY��,�7p�Y%�ЯzgHo�B��2⡆ �j���k����0e2b���ȳ6��xQ�quգ݅�����[q�2�|�&UzО�&��WSdO�w�לͼ�z�}�/	�t�r:J/6�K����q���e�Y���S+ю�",���4a�ñ��h:�E[l�1�˜��]�w,��z�| ~�� �����BDj(�R��8��7unJ66ZG �������E�����}��=�^@L�!S1p���`rt��t�����bt�=HP��L��ڹZF3QŅ�ཐ4�a�.�,�G~�����"^�y�w��K�&˨��7�"�
��!U��)���o�o�{f�V��tfD���{H#��V����[6�ژm0��w�D����LI�1���cvԀ��t��V�SD�B�X�?&�S������0P���X��&#X�����˂��	)��~"+Phr��h��t��ĽU�Lt��q� �l��Cj�nR�����_dYI�6h�����L���VɎ����u��ח�M֋��|�4�؅U+��Qo�bh�U�&�W��Yj+��ad������	]<O��߄�y��7������vgo�@NE��bi��6d��S'�B�/&�h2���4�!J2`"RUA�NDMZ���Fp� ��W�*�]x��v�@\91B����#�H�AM׃u�m_3����ql*�J��0r>���:�����'�|�dU7��R���Jw`QY�~%�$ʦǾG.��E��\ϐ��T�1VM0g����z�| �}�����j��,��� (	ǋ�O���'�����Y��aLsĪ�wb����]lO1X�WZA��Vno�
�爑����:�����\,�?]��%�jU���H�s�)ق�O"OuD�H�w��A)�p��b�Z��9��y:3��^?���N��2w،R�/�� ��y���'����������p�I����*�jD���Sr�����'X�#�%6u�N4�%蚀j�})�m��Ud.�z�Q��JV��4�<���^C��p
㘨��=��c��Ԅ'���?����	j�a�	�1����F�_�4H�N.�|@�����
wA� ��j�x��ߙ�ѽN��;����Y{��S���WH��D�2n���G��^σ5�8>�
`R����U"�&�e`h���+�}u��&� ,\ж��#gZ6"��$������dͷPHFK~��-�lޫ��R�D|�ӻ�NBK�V��ʊ<ָ26䡕b4l��O����ۤ��1t��ج&94q�L�r�x�#)Ց*_�H���cl�ڷ�d1$m}�t��w��� �#7Q\γV4�2[��}xg���-D5��T�����	�A�<�nK!��SG��L q�>�PpVΥq]�YN�b^U�{����`�H`rYN���ER;Ay��!�?,Q�c�Pw������xH=��r��?b�vH���7�ek�Ύ%D7�F��a�d�̘�S]�f�D:5����iU'U�R�迸��S�Zo�捽?m�{9�lo�9��{��G���[�	b�b�"�΁|�h��3$x񳹪{|$�����m&z%�d� �������?!�U�6��6h1���b�9
_�+�j1P%�'�#���'�m=*բ������|IF|�QLZ������Sb���f後Vs)'��5
�[�:�!��j���f�����O̞�D���O�u@�T(� 
?��-0���`����&t���c���,�+���33�+&�ؙ����b	����x��: �Z�0��M�F�A�:����t=����7�5Qd���}%�Z����S M��M�4É��I������Tjx,s3nG�U�D��o�q�� ���Y���PJ=~���	�	���c����,iQ2Ő�BM)��sUg�7�q��K��6���B}���\b�K�7.��QC�w%\:JY)����86�׊��F�:�y5�����k8��qⲟ�ڨ�L��=s�=����1Av�ъ�X#�~��z�.}y�˾d�!���^&Cm�N ���Q�ic��c�k�hL�(y�u-*�H�r3�D�BP�y�c�� �-�zP/�>��WV�[�����>"�Y���X�̻F<�i�o�(JO�1%���`�V��E;d�b��1�؏���d!�roxfcI7�L˱��90U���
�N)�P�s�n���!��&�u\�L��h�޼���^�Ѻ�A.(O���(5E
G"�X����K\�����
����(ĩf�C.�_D\�g|X��\O����Ê]�������p��
��*l�n�A���2i��F��+3����&rp��On~�ơ�'{���ÐC��TFa�D����������{��T��K�Q*��w��^�.M ��N��N�:q7V�!�17\���Z�m��j2:�����U���׬��S�Ӡ[�%���wJG��A\a��,�_��2i܄�5dژРX	��O>���4o.!X�0�j鉫��վ��I?m����z���Sm�:Լ�'F�0�� �!)$6P�f�p�j�h?�;���[�L�!U�~f��֙�Y�C�v�V��a�pŴ,�`�)�)b!Mo���f�	7��2 ��5���i�4��j�蚂�B'͵�������<b�ik��b����]D���d-2ޓ_���t�{jGc8k�������ؚ�Q,�*�����]4`䰾D��E[�����~�>N�d��BҾ�$����ʷMo���A�R�������I�!���Ke���T/�^y�J�5%�+*@=�ض.0�С]i����\�� a�F��`�rP��g6�������-��E"��X���Î��|t�Vʁ�%�٨�7(H�k�w�a�I��wpKOZOPR�?{n���0;q��Xs���Ԝ�5j�ݸ[Z��3Y#k	�߳��Y�k�܂�bIO �2��%I�>�9z�u�S��i����b�J�女����Q}V�O`�f_q�:$e'n�����2�q;�ey�����l��?�M]��Hن?ٳU���j��ݬ�B��rU�����n&�a�g���<&�3y����չ=�r�П�8���_�u�Ȇ�s�1O��۴��o�������'ؾ�
,���~�(�0M�e��1��S�n.��8>����Z�a��-.\^>�X�Ł�[3�|ۄ)��oV�CʷA"�'�lsG���F���~6"�:铠�} 	�'�m0��q`�p<�ho*fz��� ���Al����J>?�P�G1�A��
HV}�Nn��us^�f`4h�\�U���M�LZ��t{�x���&���Yދ��"��y���~`�]U�-�O�Ï�Z|Uu�$��Qv��0/�H+h�"�T�  ��W��GS�x��9�ϱ{���������9���)Yc��E�^��'�ˠ�mi���B`�Q+w��n��ܐ��i�p��HL��)��X ў���H���{�#�Dݫ_�]72Q痺�1
�?b���A���M�;k��/��9JP��p��4�j�5dcucv�5 ������hg�N�3�l>o)�6L�I�v$�5�7=�#��JH�\4�
�qf:8�;�)�~h��UQH ��^f�,����D�^3^��8ϔ�T�$��T������
�ذ��9e�t!�;��<X	Ê�(��]�p*�S���+�_�6���tlk��|��H�\H>qAV��؏i&u�m�=�x��%棯�i^x�P���#���)��yH�ʵ��L>�f׮ha_��@:1^�;��c_h�3����.���� h��>��֬�9�&���;�QO�ѭ!"�D�+����=���b<��G�Z��ߩ"�w0��;����C����\^��E-��C�y#�`���@�h����\C�@��}k�[�g�@�r|�ن������G����yL2�e�P���@&��?[C����~˒�9!^�%���a��6 �P�.N#�\Ls�^}VwU� ��E�Ӈ����.J,a��3>!ji�(ӈ	ߊ=�m���0/���?j�,�w�'ev�nG��[B�\y�*���bY�d!, b�L0��Eh@���e	d�r���Z��:o��ӓN�d/)������L�(��'�f��W)��bC�A5�D�*�֥��13�P_?���
�Uc�E���u̷5�&��k]���F���Z9��-�a�{��ɫ��m�j�LI�Zr�U�q䶇�:�%����lߏ���o�I�5����R.O��L��M������P���		��@w� �K�7�#c3%���l�;UH}�*ܯ��ɢ�W�^
��k�β-'��#X8��d_I��m6G��B�b���'�)�-�/b}�͙ S��0H&�v���\��h�鿋�
��+G�X�����N�w"-���p��x�cf���D}���?���q�������w[��"��pE��s쬜3� ����:�yv��*���+�.��q�mkW-����B˛���Cb�[��LM��	�/�,��L��NP�G����Y�����@�ts�A�wlCQ��T)^�DK�N���v�'z�"9�2��+)�WΧ��y�A�Q`�W�1�z!�#5$�m�x��D֭ )�6����B�_�HB::Z�f��ՎK�L&,n����-�miu(r���Xx՜�D߾�-W
"���̋\�HN;�/}!n�u-	,ڷr�.�O
%LX���)�~���X&�w\�מ���w��M�"䑆�cQ,4��O�h��sP�t�� ���,���O($�ogt��]�$ɖa���FR�9�a��$��4wf3"�n��"^��K���˕@l�m��6����4l���Y��]>|��uW\�'�Z>_UU�e�햒����{�m	��\P��nV15�G�!όg��V����|�,E�</+�iP&"��|86&b0k��
ʤ:��@i�t�-܇��~A!	qZIi��<�	�0x�30I6qFETϢ�#����a��R*EO(�Q�
	��ʳ� �O�`��+B/�ωؚ�ɶHqD�Z��G{�������9GkD��X�Ѓ��#��Q��{�]\JY���2�m�E��x�"̋v��gE����n��[���J3<|��"jR*?��[@���W�L�2z�+�IFo	1�g`����eK��ߋމE�@1Ѫ�ŉa��)��+�W���l�� {Z|���U	[x(�q3���ZS,R��e>�`��`�$�(���,Q�����5Nm�x�q�1+�M�Xyj?�C.#/f��j���N�EO���O:2X���Wpg	��71f�V��\�w��	�|�"�ur�3����!���KBf5����n#c>���DJG�R�]+���J����L��p;ئ�Ȑu���U�^� �zdH��Z\p��<(`�R�4{bj����X��R�t2}@9��$t��؎�N��9���$>q�^��!�!s/�蠅
N�+S0D-�`�4��S�Y�2���K3o�e����y:K����E%wլ�C�� �\S�Q�"|��kn��f��K��e;O����\�9cC�&VL`�_Ǉ��˦R�!�����?�Њ��=�c�������C�Υ�[�k3����c0�:`=0h:�e��_��6��7���a��B/�e*���k��BU\Z��)�W~2����?P�,1T��Y�5��\<�1��e������"����&��4�-�- 8�a�rܔb��;�6P�1�M-�F¯Ȕ�=6�����~���rd#�)�Yk���������(�^)��w���A[\d9�n/
�Rfיޚ���pM�����Գw�2 %��TPtdf^t@!�����K����裏��X���Xzs����Ԓj|K=���j'z8��VKs��G��?�5]��JI���/�J'���3�v��nN�Da6�B� ��'mg�H����D�Dq�Yx���@��l.�^/��i�Z�>���_d}[�n0�gO��*;��|�z�3��s2�T���EMKn�k��o�M=��b̻��m,�9W�i����2�qѶ%�|^.���^�EךѠ
r�iZ��2.�S�X����̂��k��	Ydc�����L}K<(	$�O�PJ�:���z4Qd0Q���qڵ3ܝ1��'xJ�4�7�Nx�Ki�V���	j��� L����w�Bz��ae��V����13Xߎİc�y���Y]Vƀ:��q�x���_���K�Rܲ�*m��p��$�;a4���B��I���;����,Û�S��$\��pr��nQkp�`���X�<�T�Jf�'.S&`WP�R�4"��"�O����y�����Ȼ{��q ��I��g'��Ƽ+�f'�����k�Qh.�b�Y*��	˩�q��:�)��	��������9�Li�+���EAA���ڑ�#3�Ô�YX����S��X����o$��q4'1��I��u�ж÷F�螶w�q�}4ٕ����z����K��}�o.W�i��3� �OH����=���	r������1m�6���Ģe{�}��Id��aQR���[uI�Ѽ�(����� ?�����w}%M9�B��+뮰4� .�iMC�*M����w��~M���t�١J�r����@w��鼍��V�y'k����oE	�F})c�	vL6���VG�CVv���z�8��1c쀩y��ϑ~��JQ�����q�fe��L�nA��qh�e����m����XU�Px���9r��Z��?�-�s$k��J����8�b��Vm���n���#Q�:�WY�S�����O/�r^��K����pM�����0E��v�)��	.�������U����Nz�X�C��������	�`��0ʉ��$�l�#;�_�R�����H���Z�Ⱦ#��
����%����h�7S�׸Ѭ�vc� �\|�� $H��`� ���xˇ����&�Q1��R�� >rN�)C���%�`���y�U��&���e-������^#�*ns^SO>�)B~�j,�(LI��$[C�P~�s!x��)-�A/�-�&�`q�3�~�fV�/��C�bs;̖~��"���yܥ��B����U�HE��'1�A�Ѝ�̜�Y�͞�d��CT7�3i�q2��ƒ�sM2z�%�_[~�%Q��R	px�K�JLe��@&kxo�x(�GmHi*���s�����y�L�=�O}/�Yo�U+��Y�K0(<�E�g�V�E�Ä�x|��9�&;��m��"��x��7�C]7o͔�P�2�w�@k���}`I��'�tqZ��w�o<,-[�E;5`Ǳ�)U�G�~�� �(�w�)84Q������^����G�6�}��'����\In]�[ǟ�Pr�M���R���z��ٶV��+3�M�Y���t��M�o�u���t���>�_�����RG���2.Q��̅�A�#��R�Q���������a���~�߇��S0�<!h͹f:�������XFl��l�f۹o!��R�LԻ��`�G�*(���x
'�΄cX�n�eg�>�E`�BQ�KŽ�S���wz���"�����#�ߍ���&��Qx��!��pp	��n�1PP�M���6b&^]�qQbH�J,�6��QE`���̄.i�H�W&�6����|��r�;�
�ػl�4x�
�rA�s����\�Gt�l��\�B7۪gV-�F+��,E4R���gWq>5ܝ���?����g&;%�B{R_����z:����o��_h|;#����	I��7Z�*zy ,X>6|$��Kd�/5=���.Q<�=t⁴�+�e���ǃwӷ`����Ż��Kg׽���r��7%G+H~���4�e�55�7�J�qV\��O�_�$6cEw/N'�[���DW���q�%��E��������}��G<K�)@B��������|3nQ�����8�q��Pf4%�O3�#�}�m��̒<��{�,�`巍�G�	����H��RmS���I�k5@�f���9C{�J�+�i�xʢJ/��q-�:��zb���U�@�j ��>[�j�R�MĲ\)��sm��Fܑy��.꒪�?���4�'�ޔ����A0��U!��n>d"�P�U`�Z�(nZ�r=���E|���:,�������� ����������_��4�5�-�Bڛ��Ji8�'�>"S��6/��J�+JZ 6���M�i��"ݑ�be���r;��Ib�}`��L�����LO��G�dM��������>	{M'ѧ�*)eNo�����B��Ufd��iK���T]:�S�5����:�A�F:R�S2;��/ӣv��w8�=��u�n������	������2Vil�EjJ;���Of���@��dl�׬� �P�b�l�5��c2����,�4�s�S��ղ-84�f�H`P����0
���<Ig�<�V�+y.a�j�u9��R��g���B�]"���YN��OG<�"O�?8-r ��(jur�$S¨F]x3��:����øDf�;��ʖ=(A�N%۝:�����C�.�J���!��^)��P�7�)L������{n������C��
^�ebA�c"�;1G�6��љe�G�gN-����=�o�+��'�{`h����ږށ���<�=gl�S��M���T3��Q�M��]��ү��;���2Z�8c	�F
�D�g���2�wvin�oL���A�i���`~hVb4Y�h���#���v=��.XJ��W����KKm�X��sK�5��|�[]X0���l6���+����[�/s�
�fT7������T�'#sH�>��L+���p.XG %��B3�6�R���S��\6|�
@��&(œ���x�2Ǎ{e�e��yϋJ��z��g���L@��'`�Չ�*bϲܱ0�����e�e9����@���ܰ�`_��
�R�l��p���V��,Ak�Z/���A�0�rr;�Ö���M}�*�W&��(ñ9���b��i�:�+�H�$�Gх��;�D���c67Ar��
��^�CAZ�M&(Q�z�/��i5���S�l߮�75���l4��g ��.�"k�F�Eº-���&p�h���@�d6� �?j�t!n*=���g��d̛ ��o�<�.�%�wmB`�VTd�[���Y�:��US���D-�D�ؙ���.����;S���\��R�@غ���
��~8�!J��0�	�>�#8ߒ�M��x@�
�z�ϫYR�Pf�V//�)B�� weW����/EZ(�� uյzt=�o��el�/+��F�jq�Y/�8%@KB�x{^�Y�(�}�������}0�-�E>O�A��kh�l��DE)�whh(A}�z]�!�#�5��e�E�kט��c?��/���y������I[s�Yd�@>�m:t:�&=9F{�g��A����+:jGC�wΎ�7S$$\ ������H�}��}C���ЮWX���X8��X�J6�O����W��<
zؘ��+X�m�?� �{��t�I��ƑZ��_�`0;�#e6Z��B@2º���Ϣ|�A	w����i"�v�O��Y؍��	��z�5�ɇ�@��ڏ�`���{М��s�ӥ~�<�5T��]��I3�#?U����c?C�i	G��<�����7��z��.���D;��[��YA���xqJ6�π^�Sn͡$�@3��������<�?<v�R��d͍D��/��R)�L���a����N�FI��qG��Rl�6�U�� $��a^`���=��� ��W������a� ]O�5�j�^'"lQ;�F�O�{z�]��f���H�4���qh]5.�W�:��2�����mry!g�U�S(�v�!R�/?MB�<��h��q��ڪ��0%���t�X=WNwp.,��X���6��i"�����k��
w��o����6�TI���)��*R��"��i#��Z9�?�:�Kw+S0n1�B+5Qt�S�!���������TɄ=�dÙ���9�)5�ʯ4^C>��[�8(�1G�^�j�0Ɏ3u�� �A��xvZ����d�!�i�X?���9i�)�T��Ś�V�Cn�1.D,M������I��U*���@,�w�(`T��J��og-I���7����U.lu�K�y��]H]�U��r�r��6�<��<1@0~[��n�JNe�֌.�u�X�%x1D�����V0Lx�b(�@N�k�&��Ԕ+�>PY�(Wq�o�/���@K͒������Ba���%� � �wۙ$�T1*��Iǥ���������(���:�H�>�_~������������ȭ�gL�v�+�y�s���E�F���Pd:�H'��c�����R�|+H�R�<�@�J��UN��9�8Q\o�8�׵س�4C��dZ�D^�Z�Ҫ���t^���`n�b�P�(Ez�kRz��Μ�c#���R��멱��0l�HvJ�ƖT����=�w��2x�˙*V%T�	'��E�CSx�_ޯͨ�������ў���c�f��Τ���?����,�/m?�j�?$ׅ�M�����v_ 5����ꋺ��@}�E����u�`S�P��x���<Ⱥ���۫ v�:<2�r�Q[,巇�:��q	�WV>P7��:nR���[�.:�6�1Z|}���,L��˶�d{L�>
1m����_��6��U/��ʢM-du�G�o�Ϳp�v9U��]�p+�9Br!�ad�ok�'�k�Gh�scڎ���ߋ���[)�����AgM:Ұmdd��\�H`�ܜ�-h�����^&�Y��(WL+өSx�jȆ4[Ik�fF��
� �{��`���ϟ��O֕UaMI�?�]�!����zNj�:$<
R0��y˫[�IAQ�2�=z�'5#N?g��,�'���R����$l���%
�os���S��>�Cָ���F(~��F���n���"$��׃>����>B��'js|k=�I����r��N��TTk�!��eQρw;'=εY|�m�,�X����h�[k�W�ӆ���Q��kP��æ�8*�x����]�)�������1�~�77<���^�ۤ9 N����������{�)Ow�C��n������a42
��<*J?��[|���+��K&��p���X��PK�#�$U��5O��;�PoE��k�7u�2�
����;��w�M.�4��t�7���4����Y��(KA��t�=x��Me�30ʶ]�Z��d�����W$�������������>�F����p���*ݶC��P�Ңt=D`S[Qmΐ��HWU?�;��@�����Z[�۪����qj���"F?V���B��m7��y�q1���EǊ9 /����2�[���h�I�o��6���l�N���;��Ŀh˚֒;fog~����/Y5�s���F��Q���$�����t���e����+HB�I�aHt05�}U�Zu�xÃ�-�_=j��c�U�j(��c�!ˋ�x�*��J>~�#}Z��mVSݻM-Z���-mt��3.��ne;g㖒+]�Ly���]\Z�%�;�&�}�3 �T�D��Үa�Q��os��I)T|���e-��܇P4a4�ﴀ	�3c��#�q��<�R��� b�=��g�"���Q�5y˩lU��
��L���bgt�[�}��Y8_��W�U��8���?���4ƅ2�r�Bg���ϲw��f,}&���)H�vc��B�����H�RR1���j�w�RA5誡1�Pe�x2Ӂ9n��D<�n��_ r�ӱJ��>@��U��w�uoJ�.���Զh����Dàb#8��S�����l�	ڲ�^�-��@tq�$a-;�ר]�H��S�=zV��S\^�SҀ ���v�+l�;��#�;s�s�I�c��d	��+
�i7в��G�s� ��t�u������m�P�5_18@l 2� S��wg�6�nj'�اb�[���V��w�Jd��#H_e}���e�<yϦ��H������	��dX���X�+��r�|4��+�1�,{�ZϢ��a�C��sw��~~�V�cŴeP�tc�T�5|�q;�R��m�;�.�Һ��.UHD��F�9����d�|�,��Xn֡�9WB�J;�p��c
L��hHӑ	\�8�S�U2uW���/-qfl�M�|�����]�8��KC��$u"!fR(Ca�$�.��)�4�뺺<UfM>�O�E�Cq�
��{b8���wc 6jq�*P� �#V`W� ��D�UqQ+�*.E)O7L����	��y��pm���glV&O�LL1y�Ա�Z��<~��{��}�Q~��^��p'��.'�ݰ��N�6�'*0_ׄ�˨W���Kn� ^9g>�Z��01��T����Z��=��:-q  �4�Q�H��-���MogyJ�C��a�}����s���F�i�W��Ii���Ԅf�H�޲>��M��X&S��8a-)O�~&RQQ"nfGp��v�"^�l�9\�rQ8/���� �Q�(D8�r��׮=r�ya"1"�dO���m�/]
x���Q���������>�1`����B�� �D�ۢyݗ2_��3���y�ӳ�`�Z$]B@ �^��v�1��[՝W�Bw�+|���yi�D~���sM�����%]<���H����(x�*ˁ8k��@_�6��l��pN��lR�A��Sim�S��%2BT�5��[g��nB$�'�'�%�CK���+`�ʹ��2T�� ��O[Y5;@PJ?�:nW1H7^vN��AQ#R����{�������aa���-n�P��,���7##�`S�]���}�h��\�Ut��q`���۹���33���BW$wM����Kp���k�59~�pNp�:g�7	0�%Ǒ���̎��-�`˗�mnV��d�:�'ߝ����e���Ν�"��@⻚��)��<���݄l�r�����@�cś٦oppp+���Ɯ}F;�S*����8���� rm�Nh�a��N��g�)���ʕܽ�Y&J���-֡�;��WmҸ� ��� ����4$W��=��ScՓ2E�Y4(���h�E�SZ�u��Lgn����aQ]�wA�&I㎽����\���[�6R�6�ژ�ZǦĎ��S�a�
Q��ڼ��V�	��hXe�V����E���+�U$R����չ�&c�6S/��W~�I����~�\��a�k^]�5X�+��i
c-)��/�Bְ'�Y+�|u�8���j��<�oeJ����w:ԹCJ�4�2�� nԸt�A�A��@�r5jb �;�u�	ACqSQ5!��'��6p����㒴+���r~���诮��E�2���M%��=��(�W�(��4�<���k��X&?K��'h�5���9��^!ԖT��K�j�ip�����lb%���m(���ǽ m�S����P<�k���	�+�@�k����u�=���E����Y�$[��D}I�S����U�ڈ�y��y�3�6s��mF[��������b?�+_�S�.���}k-�����n��e��VOV��?��ׄ��@/Z�Xr���������6��ճc?&rw�?�(L�5j��!F��Ӯ��ڪw���
k�W�_2�Q� -x��9�+/v�xk�q����ƀ7s�U�<_EZg_�Ta�׏+��ŷTQ��#��`�4����&Ѣ����E�,?�l��T4dʸ�����"�o��K�ʄK���_k�t���Aۋ��G�~��$��Nq�%[˪z��D�� д~�X�1�N�/_kU~:Gѷ�k�UA-����1�NtY��4���6?�UDab8��PTdY��Ih��������͕.�%�H��Fj�bo�{%�I�F�I��S�O��*K�ʠ��}���;�Zx^��)(˅�|�\-A<�X����҆*��o���m��.���&��F��"F�wN&{l!�u�$?�\R����5>N��7��2b�����3���#w�.�6�SƂM��r��*`���j9ʗ�0L��*x~ao���5WR�uRM`_㨈�G�H��/d\��2��P�����q�׎:`|H��[����Ap �E�ܟ�V�8��j�0�qfNz]VM%�l`��<sT9#޺�tF���S�BL_���� �m����?��c���)��:���	�DZ+���0:<k֩�g��6��O�,��/��ՔP}Pԫ�V���1w�c�a�SR#��C5|`Q3����㡾B�cY)t��K��֗��xu�`���{�U�ꮯ6E�aM=��9C5�C,��\��R���69������v���W����#��d�d�}y_=f^����j�-�{�9�\2!B�L���evI�EJ��ca�褶�Z����T� @A)h̵��.�)t���Fp&q�?amڈ�bRr�[�04�fP�wx�e�=Ɣ�%���g<�;�Cn`+�Df���n%�y�(���Dܟ0ǁכ�ie�K)	]c[7>S^���tkQ�c<���ԅD@4��3��˅�]3�e;�~�H�U���C���a���bɒ���t�p.����)�ǺJyO��a(�v!�c��,������V���}� ��^�Y���Dk���v�EiAރT1̳� S�T�7'MG�я���[�?DJ's��ҿ�W�멼6����k�����$��֛z�?\���Q�h���>�������~��Y�QZ����J�W�S�N����Tc�b���-ʄ��D���9�>�7��Kma����?���;���Ğ�Y�,���v�I<U*74�7����$�oK:Mf��.�� ��jZ?�5�$�A�jljC�Q�-MW�a�~���apF��g�X3jj��ky����n���=49�Z�0����w�N��2��D`m���ߞ+�K<�){}X��V����,����(���X��2�.+o��
a��l~=�:������;%$K��X�J-�K��U�Y�;l���9d�ljڊp���ڭ\p�r�Ynm�3�� �ݝ�R�;h|ҭ��8�cG�$,�q�\��K�uTJ�ou<hK����5Sf����	$y���hQ#ސ�t������㹒j}�h�{̬\���n���M%�y9p�zt��L�D�:�D`�Y�V�����n:N��m/�Y'�MO�a��gŷ���3_�e���s��옠y�2H�~��ݕ�U�Ď�-�%)��)���#��N��S.�R���V`1�������
���!ķv�����_�O�T?r&����X�v^\�]iD�\��lw�Q�<��SC��܁�����!H4!)�� ���ІÉ���:����cSk�4��Vc�bE�{.3�[.�L�dJ��/�.�a���G�a��mk��e!l-��.���T��p�|���k��Qy��.�P���d*Y��[���_�{M0�,����@������`���c�.�3��S��P�į�$���3|�Au"4vR�A�e���Ƙ>GUO x�(�����XA�����;�**�ee�	�����|);eKC��� ���:������{h@<��xI�;hv%/�ȱK�?݂��^'��SpY+%�p\�Ӿ���0��ƀH/�H�Sʖ��,W���h`�����G�P����bҧ#��q�L���b�����6����m6m�t�*+�ӡ�0>��|���e�R�4�]Z�m�qm�я�q~3ꈙ0�,Y$7�����JR^��Z~)v�g�6�]!��d�xx9\upC���@��Y�11�g=�y��~�!��ߞ&&�/�G%��;�A��=> ex�>:������q�2p1�峋�J���=�{��9~G@5{�ݼqC���|gB���9s�}&��;c����lM����1�j��:'?R�9a�/׽�i�>�u�?��3p
��ɨ�/�;:q6F^_���h��F�)T!���1YBU��J��K��x�i��p|z��P�zh�W��˷�	@`�qܽ�6���j|>��2�sB#CP���'�kj׊jmJBǍ�v���1Ԧ����?�J�!�;'w� ����]D *��pӄ\1�g��rs�K�R(���R^ayx=�<,wX�i��iY�ʓ50J��']���{|4#�кwXI�9Ԍ W���i$��� ���d{l��4�I+�yuf��MTS ����=��!��roH~3:�Ts,G�yڃV���'�7e,���l~%ezY���b�"Ɇ��ċm%L]#�J��k�����\q�QF(݌B]?���%�_��t��?PX�$rҖ���6�H?�N@��h�,w��T���/�<�Ʒ/7��%�xG]�1u��iTîjle�j��V����Tʎ�� ��:��8� �sl��c�q��/̭�����~�s�aj��t3���{�
x}����{�8��>��	E������p�������3�r��\n�	�/l9r�D�����%�������H����9~�/mL�.�0m� �ɱ��L�U#�G.��X�2�x��S�c���dz���*��@�//&fQ
:P�����v*��ܓz>P���x���AS/�t�ᄡv��7c9���g���� ��"Q�oac>�f���ʳ���"��I��d���t����́R��,ZD��"$9n͜�"�O���J�!�`N��K�K]��ԟ�/Zp�R�ʢ���bJްF̳�����?��,D-F	�g�B࿩32���#�Z���rA �_�塓���_�����t�J���,Ѯ��� �� No[�d�yd]��&F�w�{�پf38۶lT[R�.x��M+
�ئ�߄.����߄�����p8�@_o$2��K�m�{��ǻ��H�DmϷ��2J	=��L,g���u��w�'U74o
=N� (���ѢLx�[�y�	͊�w���d��������¬DpQ�N��F�%�\��+A�|OS���G�}SȎ!L������	!o���α��X�\��]��(ϘM-� �fN�8y����oE�S��3�M!��ױ���zP�2-�M�v�k����7@��'<�l���^dcQ藖b�ف��W.�cgH��`p��w�A6���nJB/�车(᧳���'�ʕ��nZ�~��.d��D.�:.b3x&p	�p�>��Jw��ۨ�=E��ϐ�Bɿ���t���bF"���bG��X{z������[t� W��,$!��>!a]�L�=���k>=�\�M(��
<mΟ�a/�CF�֦� ��ɫw�9�L %t��g2�vF�������.hC� �^���ށ���J�	b��d�����E��<��g��xa��O��I��T��g�Ϋs�d��{�>�F6�?-�d��e��a(�����e�XT���U�8J�p/=��vV�n��\���A�H����	�t*�Q}�T���z��v�e�-�&�"�n�0׼�K
� n�[UL��%	݅���w��ӫD'\8�����nD�}��:��[�'6��jD�Z�{R�xɨ��[�p���@���]��F��Co�,%/]O�q�AML�����㬌�3羦�X��[�
Kp$#��/������ټ4d��Ϧhk(yI��
�r塊�,�&=����	:�5�mւ�m�Q�H����v����W��cd�;KѶ?��ȽW��bk����{@���)���\J��Crb��&n���ޜ���I�n�d!{xs��?�R܌w�}6i�2��\�;I�GX@��3e}"Q�Hƭ=�cR�y�7"#�� ��k��_�k��6z�c���MS:�
�J��h�'�X�����-=��3P��ۅ�~�8=�U̍��i;�Z7�3��j`�*��f���!�6����Z�הb���9�#3	|�%
]��m���[���7x��Sʹ��.�~��+��q˕��v2z�RѠyMl��a���MY%�5"��m\ޏ��ڜA�<�{��$��|�>�l�	�.��"G�v �~�f�Y]�?g��#'�����d7I�y@�d��ыg�v1^�zp�H&�Y[��n��#�4����A{��U?��,���z'�� r��m�E�ƧQ�1��"r��s�]Y�d��6�S���уi�����]h�[Pb�l���ߘ�M�B���F��Nl<��m�'s��Cr�d�ڤ7����.�fu�U�j�b�~z��!���
Ⱥ�n���
1af�X[�A��iR���l��iwGc>xv��&������Ѱ�1�X+2Gu@�|Sу tA�͚А�++- s��j�~�R�amU�)p�,�ZfhU�>���m�s�XO��n x����1��}�+lqo�}�E5%U�x����U8�����nu���Ũt��ĩ��"�f��N2c����T��6M~�����ATS���
��T��wW3d1Ucr�eU��f*��4.,�HBN�3�p�����o�Ō���p��T��� ��R��o�Ql�Ь��h4}�ɬ� \lQ{(�uQ}D�a
�]6���P����H5+�C*�����-��>nHnY���KF��D�_zΌ�$@S��؃s#N�,�d�JY���{�quJ��	P�K_r��LjV�T�-����t��A��8�X�(v�WM���Ƽ�Lo�K@�r���2'߯1�^`z7��m�����K����?Lo�ꄨ|f4S�e��P,�����5���������?�9'��_l����d]tڡ<�7;�:�9F�^Tl&�1�uJ�7�`>��^�[���+�8��S��؍[Q�^X�25�:>�/�|H��nAS�=Ҧ�<XL%<��w��
�/�*5)ƾeA�t֐��y���g�<�p@���9�єf���S1_�f�ң[e�OW����~F�Fk�f]���$�G��'�I?���)�w�E�2�k��K�W����f��+�%�C���'u�FtM<.�V+D$L���ö,�7=z�s��L-�kw ��N7��V�p)��Ų,%��_F�����̣%2��A$��q�d��6����兮y�E����1pNDu�r�������ހ�Ȍrf��ިM���Im!t���&���~���&�' ^���Z<�<]����N�V_f2T�D�<�|ܿ���tf�G0����Ӣ�p��sZ]�=C$�H�:/�RaV��ג�9Y�@��E��>��l_����[�N�G��Ʈ����X~8]t��J���U>O(5��ǝ�a@1��w��7��Q�ix;�jn�>#�v���sYҼ�DQ�?��qr��{�h����p�ޝc����J*Ny�]��J
T����C�*q��˾~+n�h�q�\����y���'R�p��FxL��A1�rl��5�=�6��|��Ǔ����I9͗��P}v�<3V�>��0ʽj�l�hN��|݋ C�EyJ1x�֗f�|������)w�'j��I��O�Ҹ:ר���R��pN��	"*���=���jlR���I�whL
�w�@9��;"�y{d
��u5�/�fP��L1��A����qc�&�7�L(ض������>ͅ����'����� ?#@m'�g�`t]d���/�L.;�'���zy3-�9���yvd�[�ե��js�ڍ��#������ۖ�p��~��e�m Un��Nבuk��z�!_k@^-�8�~�UUr4�~��K�W�rP�*�%<�Aހ��F`�S�+���R"���2��&�u�5.��V����9����U���Ȥ�W�]M�ο��SZ��3�� ^X���/��i��������\�Nz���*���+Í\��?�~�>m������4k�^4�^q�G�_~��������z���e"��W�\W�����!�H��=�.���ԯ֐��t� 3�s��B�t����H!g���0E41r��rn8��E"ﱋ�R�������~`_�DUbp(��;E��D�9��}��&�R���`�fRK���
�h��=���ť�JK�h��p��N�~��lG>u3�Pr���VNARy	5�۔m.n��p�.K��S�x%6Ƨ撻���b� �B';@ȹa8�h�3SLP�ե��t�Å=p�^?BUrI�C�;F�q	Ҏ �|�i�bA`�դ�3��Eh$�����z4�Us��,�c�' ���?��D�%�� F@`	��<�)���>��u��ҙq_ٽ}�^Hf��2i�M����T�W�݂]QK�j�%��,:3�A��`�%tV�����N��6����f�Q�p�AE��b�]vS�"*��I`'�� �.j���!���=��ܣ~�+�	V7�h��2~����N.+O��:U��%B�@ȶB,�ʑ�a7�U�ly�O�xF��%zDDq�)5�������X���h���r�K�,�:<u��7�HZ��:����`�G������f��)�.�4`j�'�����]����%�aL��Z9��%�k��0Ȟi��Z�+�XI��)���﨣Z��2�zi�1���e.Ӱ"�FSJ���i�����l���l��Ҝ't�v%%���㼑'���ϸ�^���*/;^���x�����/7�Bo�a��i��F��H�KV�^̙^a�90qM�&7$?#8ǚ�+���GAy�k/�Rj����q�-ny�62�nm�C�r��!������dx�z�&�H%%���|�`���*����T��Yh���N�ӄ���pEN6�X��[����<�4F~�v��O�PWM���WI=6v�y������?�0�Y� �יִ��^��j�X��8A_�>%WR�A�k����̫e�׮�\��"�%�3��U����A\%���7�U��t�e�C����Y4�]F(^T����F��#��)�)����%��0�$VP��<e�������^'`YMP��X ����7 ��c#����}��;�`�<�D���r]�I�NK��oA�a��rz��L���1[�� �Q���  <h9���kx�q�!`��]�"XN��щ�RG;�"�&���pU/w3N�q{��"����`���6?B�bBT���~W~�ߢ4�.5�I�8)9J�J�"��OS(,B�sK��m��M�'>�=�R6,r��)����G��w�',�?|H�G�k��n��k��e�|�a��1D��*�k�>
ν�̿F��n��=ǡ@%+i+C���yN�$����7z�F����~Q|�P�3�E�������3�F���DZ}^�����J������v_)p,4�H��ON9R��"���$0g���/��l�m�u^O��gI���D��ѹ�̥�[��\�H4恃T��ݵO8�Ie�}���Yt�4!��5���3}�@��Fs=;`3Ǝ��T�(�8�͏5nj1���Z&	}�VZQn!�Ċ3��:��-��ؙE�����`��.��U�������.����!�N2���H�3}/�E.��E���V�X_�<�(��6	/\t,�H���8 I7�r���˳�����w9dClkE�^�PF�'��W��w
��w��W�ؤM������5���r� v�Uܩ	�!?V�T�b�Dp�	(cK���������.n�V�h$k�"����
wHi閁�����r��b�.��$�M���3�,��|��T^b0�e�E��e�F=�Y�Ϥ�=&|����� }�T�Al��ޖ���X/N��r+�s�7�`�P'���Kw@�s�Yn��:�O��;)��Ȁ�I�ԕ�p{#��Wv�1纕X��
kT���
��~)CzK�ЂO�T�<X��"\\�~�Q�Ne�� ����b�1Ͱ�ƌr�Q=�#�	h��jYu�h��,�`Rǝ|�V'�۪n� �Ɂ�����~C�8o���ς�q�PiT�I��;:�(�%ʕI�vF!$�=��oQ/�o�쳈J�ޙt��7�ݗ���.I����i:Ma�ԥ��փ6�ʊ}+�N�-���8b߮/J����ft���pj�<_�+C�A���Z>;&�P%��P|��Mm�+zZ+�̽2��I�Id �q��v�����J?��)��%�p���d��w��!H��m������ަHJ!i.[����S��h�*��&r�����-�'����*�n�غf�� (�ep�?���͑�0���e߼�zT���������	�zv�n�\|��3��|U���<��
`²����a�����^C ���&]L��A��;���G? ���J60TfoW�)F\�n�'4� !:������@�D�B�3�+���Jr:*�F
���L�S�?|�T�l��4������~u��[����Y�*�̫@�̴f�z�u��l����������k��߯:�y��ʰ���g�Ίz~���/V�! �3��u������"8��s{j�x��`��t����fW���uT�)��LA�M�xS0�om;bS-���A/\��HkX�'k̵���0����Jx���
���aꦾ��=��őq���r��f�J�	Ȼ�O�mG�"���ExZHv�-u�Bw��1bYM�R�L�v�]Q�	�����3�7M����:�ŃD
l��:���� �io���H�+����c�@���-�p��n���4��< �z'PA��:�7;nG�u���Ŭ����8��e�O��b�txX�h�wo��G�B!�y��l�qx�&�L���i�.M �N�*3���A%�:��8����V�,�k5���X�wNQە� ���Z�eX�!4Z��ۆ�ԡ����&���2\E�x1rmR%�α��ɠf�(��zT�0#��R�Ux��㰅UK��	��1����Ր`���*�����?�X�0���Y��v�Q��~��t���zc��{�����u{�Ǵ����"B��J��lG��gbƹ`pU7�cv!$�sR���o\�;�*O ���J��L9�6sj��O���Rv����N됻s| >���+��-
��e,�Ӊ���)����t�E<��(����:	�?���}�[����^�芻����ȋ�'�d�<��=����5jTCe��� �DVss��vW��̴���#��Z��a�^�+�r�0
��p���Q�M�#�T�58���-�޹y�h����zu�-˓>5�%I ��Z5h��Ӵ��!b�g��W2�pt%��{
!�(�ۘ�����!�[�]2V��A�&4P��)1��:�i��R�����J���<n�*���Nyp�S?%�8�fI�x���Z�������-҉���#b�rr�͎?�Yv������c%���-?�d����
�U"�,��>qs�u^{��1�9����*�i��|KI-8���D��_y5o]$a�V�r���(t��"(P@�7wkf9_���S�F��ۉ'�)��sߗ9��@BZx�ip���3�3�뤦���ǣ�8{�w�*�FԺ��0�vSÇ�p�!d'}mbv(�#c�l�bYEӀ�>�s�}��9Ɲg4K@��P#��4�k`����Q|�Q6�)s1ZӤy���2f�_������çh�Z�{��?���B�J���Bz%X��o��v�A�,����� �[Tq�'��"_-̓W]����&�M$�,I�����jn��@O.�Z풖Ԡw����h�6�%��m����h�v��vEj
����:t�䈏F��	�p�\�k����L��q��6C�Z��e�e�k3G7���%��E��b�o؅��g�|e��qx����3יP\{}\���[aq�{�"�п1ܟ���e�A����W��-��q�Em!��$ȋ�&����HA\���)��c��pr˽�C�
��+�̙U����'�K���z�`;��-�Zp��m�=.��{U��]��|4���@��[���+ iS�նpw�����F�i_+iJ�fI������I����48�5k�.��x�����k�D�}�L�6o㝊�O)q�G�B��hǠ��(���f��ʗk�_܅�����lA�pF<G�`��O����Ft�?Gھ�T��f=�Q	"�D#��!����ti�fj�{қ�=L�Dh�����"kZ�V�
�X94�kv,��e�3Ys���h+u9��&�Kǹ ��a$̴�z���ص�T:76%���O\=gFtM��d���)��(����e��!z�(�L�O֋�s���5@�����j�Ğ.;</qe��{�/h��G��m�+�k�@[�����vȄNe��|C�n��яW�s�Q�?�?�d��n���o���>rצ�����&am<����fR�(����k�� K5�V���(f�4�w/���Œ�+�_�A!+��oR4�Ԫ��L��S����ͣ��]�H��;�}c���g�<S��*5Q�y��ya#�ٹ��Q�`�nG�I��Ӷ��	��_@����n�^�M�D�ʭ��[��́w�]2\�*!Z4�	�'���H���o7N'��NJ{��
�A�'��%�0d&8l�a��j�l���9i�"{�ˇ