��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>��p�������~��7�G�����`�.�6�	?�D����VI+�)B�{;��������ii�j�Ke��t��2ߠ�q躤!0Z�� 7�q�������$w=f��Z��oH���#6e��re W�E���ı������F�A�7,�	d�'%|X���I��!Z��g��gyգ7\��Y�ư[c?��k%3C��T��̵Өfnk��FS]B�З,]d��O��E7��'����2�=�r��yq��p"�5<���X�q_�?/���YΑ��M�\N;�/0[��X5L���s��&I08	|�\�վ�|�U$p�~���?Bva��(�E�H���n�-(�$U7��<����KZ�pE#���{G�
�G�e�;��Eh��]�j-�h�(���i�^�ƿrh���ɴ�pÿQ�^�z���@��h`��d��V?>l�8�K�'&iҺ��Q`�g�x����&��9.�hϜ����l���
M�Dv7d|�V�j����/�;Pu3T<,I4���6?C+^P�tG)��b� u2��b���3Ȫ�O�NNJ�2�!ohíK򥩠K�]���pMV� L�=~���+�����ڬ=w�Xn�Ć��
S�f�
�w4�l�L�W�E9���,����r�E��g=�U߫Ç�n\�l`>Fll���}���n+}ނ_p%�8t��,���ڼ��B�:�(#2^C0�lC��ʞ+�ŧCdl��{�h���.<Ё���}� �C�,�tR�X���J$ߗ��^��w�gg�	�PN8gU<a��ԎC2�࿿^bJ��6yL�
�lY���\�����\̮nw�fp�S\��m�[��׼m����t!/���ΟQ���A	&��i�JsdO³	��}0��
��K��Cu�0�W���8�ӗ��m|��*��KN"?��Z���f��A���i��[�5er�BU=��V %/�P��#��ڔ3P�w��\���mI�8�1��k������$[��� �!���0j�JRsbC����M�Z�}��6\�ٯ�XUܤ��օ�-��L�~<>�V�QLY�g������鎍>���9�'A,����7˿R��o1Gu�1{Ȣ�8}*�o9����m��p�#1���rDW����S���?N��/�Ў���^o	�gz��O�>�P����g�OH�]�Λ�֪��@	4��.b7yK���Nν����G��1Y�bl�E�m�0�!�e�3��C�[Q���K��%pG�b�-%y����X;�V���N:��e!����ELZ.���u�����y1�O�[��Y5D�o���|��ʗs���St@����-(\�12��<�_{���۪�C��q:���~���n���E�T6��D���	��T[E%�i�YE���/����I�o-pFR��Y���8���|�$]IH^�#�6�ƙIS�&g1�0[nt���~�6<�{��nm����\���b� �� �)#zTK/�X�VL�7��;���Bm�s��I�ř�����o�� ��J�PLxm�(�T]��߉7�%n�eC�z�xgӂF��i|�����+�=p��^�D��X�B�¼�Bu���&�̼�S�$����,�(��#��E��LmB�G`��k`߫�|]���~�*���]De' [�}c����|U3�
��l�ߕ�3�"��3� ���S��]���e����'�<V�Rv����>5Mv���B�:�	�pI��V���m�֜�=�n�}q�S���Z�F~$�#^��UƽQ���M�`�[���<����!�h���Iv��
�/)��<a~Km�7�?s�CN������5�@�І��L�N�4�U�f+�8X\<%�Z���͘$d~G��4�of�Mn	�57�aG%
�Z�E�)��@�Nᢔ����� Q���pPd��9��t�{�3�^X<?N9�����o��=��`��Ҟ3��F���\�� ^����0W+����W�_8��Y�a膝2?�e�n����j: {�yA���R�O�z���px毁#A5d�T��bJ�0W���l�A�A��)]�,��L�}�y�M-�B��G�nYP
�N��N/�dեs$� 	 ��JࡹM���xF��Wభ�m�7MI�����{�F	ڄ;%��J.��D�j�\{�`��XlO)�>J�}m�C�=h�Y4��vS���KMe�����9�P��t_�5U�r.��Cw_�����1*yp�Vd@�������[r~*ҳ%�K� Vqo;��b���(�n�HU&�U��O�K87��gug�T����FU�P�X�*�d���&WW)�� ��8����ڛ�J����L�d�V1����,��@�A2VN�������	y�P@� �2�M�L�9@vв�����B=;}:'Q;�|��E�E�O��i�s�p�r�ܬ>{J��$�4.�e����a�gs=��2�8���2�i@���!/���'��nG�8޷�Gs� ���ϫvA�<�T��t��q?i�:0۰��VK���n��.��%�R�M/&2���Lz���&3�~�h��lY�-�]:t�l��S]�.���4S�d�ج@�{�\<��~�sZ��0쑫|C����E�aH�������|����k�N�a*0L�l�x�������*�c�WRB�iMt)͘״�z쬷˜�|F? (��?���F�5u��O�X��Fɮ�
��;�L�+}��F)�ud,�!��H��5�+b��`
1�چ��wP����l�݀�g�Vm&spk� /���[u�}������0R��
�~zK2L��G@��J�?-y���ǆ�\��ȥ��R?]<��N0L�EK��-K�'7���)0���s#������m{^kȒB�<}�=�5wxPe���J�K_��PH�h���v<�����96;˻R�c���[�_�=�p�ѢӬ�cq�2"�N�wv�5�g���!��4��2gz�wz����Juj�M;�ka��*�i~��~/��B�x(�u�a��C�v��<)h�h�.�XO��Aiq{��H����X�� �X��BQ'�c����X5M����Ȗ�5�ӵ�%��1HS��i����_6+�䕆K� �WUA�o�B��'�¶h7>��?��F���@ƥ�ܚ����<�9W޵��8��8����;k�$.�� ����(�Sb���}Zlk�џ��G�+1	�����)�&.9|ف�5�j�W���,z�]������&��3�Z���zk���n�z�Nj/�t����Y�>,0UX�#3E0�&(̃��(y%-��+��O!�d֠��0.J�~�YXZN�7G3bZ+�,�����'Q`��l=)��X�İ��Ϛ�Y{5���+�t�5(�P9$�Γ��Qd��X����FQ��ј��Շҝkc��(��C ��^����� �����6�0�[D�q�������A�����TD���j�h$ї=��}^��m?|*p�XKhW�u�� Cd�x�?�6��g�w?�@�6�f���=@��Z������`������\M٤fDƼ��`����<��ֆ�p��Y��HWw��^@\:щ�J��:��CjB�t��yI%ms�,GL�v�M@I�#��֦rYt��oԙ��Kt�áwSIW}�"!�3Z�Bb�߿����r9z5{���{ws:U{�b�a�`��|��6�Q8��xK����Txo,�� gP���0c}�A�Mn��R���: �q��am����c��2Pt;�i��\�ׅ�jU�X�N�BRKR�*��o����