��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��˲�|U�eu2���P�1����J�2�@y=܆��X�n��t���+-1#Հ�B�H�b�~"�{����;GH��Y9�QR��c��ׯ�b�i�j��Ñ"(Y y�AG��) lW;#��2��rn n�c��n����dӻ��4q���狙e};�e�h����ήr���[�̉���Y~
�-�ʙ�d`�d�Y��8���N����j�B��M��tI na��#B�`��f�v����+�~X�<�V���~�����p��ӕ�i�:[�<!n$
��� �.a�5���tVm)���ݾ�[���M!V|' �����h�Vb-���+Q�,��i�}z�[A~���Ⳬ::��Q$��8}M�ׁ����fh��W'�$�CV����Ԭ�\Z�UeU��Fk}�BY�k���v���˿��E%�
�-��5������s�ȸ�nF�?8���勠-���>�Q���-M���t��nZ�L�!�7y�j����Dj�`�0�l(=�]�}�bE
���,���Xȏ���꺠��B�w,��|��N������NzԴ��=�_�ߖ�%�&�I�f�:b��)bc��f���wv+,bg�yw���'Sqi��W+�xM^̻��r_$�;R� T�F�]/�k�/_�[�}�؃ן[��X���;�
K2�	�ևA��-xR�7����I_����q��X0�G�}-Q��0�KN�e!?����n� �`�'�o�)y��9b��T��3;��#��Tm\� T�?�X�����e��y'N����ێ�g��h�h4��:�����:����{V��p�A�q2��Y1|�0>nR�����F 2��/�j��G�mJ�Z�9�}Y�39�$NhC�MJ�<�.@M�@4��N��3�c��/9M�,�m V��n�������)W%���Ɂ{�ۄ��.�`	�w�P٫Mg�R�w>��� �LW� U��z��o�Q���'���@�� ����~�O�~ཀྵv�@:!Z�������߅wXj,˦94j�6i^|z���P0_S#�-�����{��J;��W�E�g�%n��8�y���)Gݷ�p�=����}��Z��v���a.�k�w�O�a�TW�s����/p�c��%o�" 1~�[��t	���[��^�fA[�������Y�N�v�$���br��~�/؋M�P�i���O\�$+{SL�z0;��uu�A�*~4�����H��_�!
�E�D��J.�Ĺ���؆�4��;���YVD�#5��!�w9���A� ,Vv^׬L �T�c�Q��X2MR l@C)��~G�f|T�ᚢ��#�Z�=gQ�����f/ac�����҄�\I��&�Q�W1Z�U`Z�_\���#�@�/W��4�����IB����N޲��T����4�0����
�'�-�YA!lJ�+E��`���<��ng�^;G���_�S�iK ����h�d��_ ���a��V7yPvFd�k������Q���B��.�U����j��
�uc]>���8���rj�Be�uD�-P��*AK���i�yIOr}V�-C���܏���;��w���`�8�l��Կ��R���7=H��w�4�ࣚ�F���q���w��g�f���Jތ���M��d��В�t�2Z��1t1���GvS!�L���bSi!�=͊8ld��1���"e,���
�����+WjjȖ�� 
|�Ԭw&%��4����R7:��p� �~��[�#���4��oKA�֏�N]ǗG'\���e�t�����@q
so��� V/6,��A��yd�@f��z�����0�&'�bT�e�WLu-gf�EZIB�:�Qm�\��mx��+k06s���6
2B�J{�C�ҼrD[�;����;4_�
�>v!FT��>�@�����Ψ�e��l��u�mw@O�S�	O;�ɚ�s�m��{���R6窻�EH�o�2�{/qF���� �Ė�]�:��ƒ�O�2S`�V흷�R �&�Ca�����Z��`QH�1^M���E�y����¸���m�	ǡ%*fRُ��m����0;!˅�
dH!g��Z9�|�7����$C�{ Y��&X����7[�1���|E�86�:������n������X-�[mäS)lD�Ì�"� ��ᇿ�3~mU�2���:Ð.,E]��f�H�����Y���l!���<(%�Y<�@�������>���K� y��.�:�֯Fc�*��60h���K���h�Yj�D�E��/�y�iḘ����2�3E�HTXg��ƺ���aH�s�-�ث�W�Gr�& *� vXN����\���:�w��Hc�Xq�Z���N�G0n��H�~.� �2�y"ɝJJ&!%�}ȱ׫����)B�|?��e�kV�t�x�e�UB��@�("PTdv�Om�v�f���k�T��P�q'OA�L~s�!��܇S�#�_�ls��9I�_�>i$�7��4�<�`���5�|����ph'���;�s�j���%=wh4�z{j�jJ�C�8{)�h\<�d#����.b��it �8�%я��/9b�΍����m�(͊	'��Z�  RQ���kВ�J��p�S!��X��(��A�K�.-�SgI����<��n!uwiaﴭ��b>����U\�HYʏ�ҏ>n��P࠿d
�xn�Ƶ�N�J��Z�T&� �Ue�d���g�>R!$|�7����x�Ǹ��X�Yڙn4�زm4C��r�;�whu�ð]�W}�V=t5IC�m�]��VCU�6�G~�C����8��:�d)����kmHMC8`����p,%�2���*6,�m�$��!u|5�.[��l�Gh¡�ڀ�h\T�#y�C�Cuh���JҙɖL�W���uT��S�i�W�}���S#:~;�y�I�w1GKa��*/���]f�q}#q��d�J���j$:����P�!U�TsN߉���@��t�,�Ki��?P�4}�@�[5ZB�!�`i!���l�ͭ�H�����D:�k����X>�~��Q�_ǩ�}eJ���&�兟ߒҭ��P5�����
�ڀ)c��J��q3j��.ن��䄒��B�R�tjN�%o�r+G7��_�Φ�G�<����`(�7���&|i��k.��p�.S��2;-x�z��`���ZQ��ڣ�*s��h�1 �&18\�v^J~�n{35�|t�V0�:*����~a�a��|�5!�c��{�	��!O�VT�y>Gɶ�j�6��,b-r�hEkN�
 I�k�Si���,m���#&B�5+���K!��,�%��Q�G)��We������p����H���/�:�Bu�dp�E��e�-�&��4�C�m�`&�O�\�\Tcq�G���g(�	O�/H�C�����A~�59�$���T���q`ș���}�ㆣ�z����m��i�a8��<R�m� �c/
� �"U�N�;���H�R(�`>��k��J�+��a'X��X`g�,�z���F����G&$�y�^_��A��_��CW�U6��'O:�SW�-�<��;S9��N�=�(e�<Y޿ �
M�Y�#�:��ܣ�X��
n/w.w�q3�,l {~-mn�*P9Z#�<�	ĩ���.��j�gҰ�j�bz7x�|��<��'��t�����Ѝ��V�H�}�Н��EbK�Ɓ)�솀�f�iB3]J�r��̀�N�X�m�y�IH�����䗐�H�P��bO�h�F#�.|g_�_ײQ�A�<[��4�t�D��x�X���x4M��N+ҏ
�+�P�|�>-�c{/LK�!k�ގ�i���ZEʷ�8��&h	w�i�R���f�ITP\�
	�T1��0ږt�2��diR��zf�M|�E/�j_���.�<a��9ܰ���� h|�M��:�mR��|�d_�C��VNk�v���#��j|��j�3a��6�!!M���yȤ^�?���V��h��ܖ�}�pvAQ ����T�*�UV��Ng<��ht`m�t��2��:[�D�D��#��\͵5P @@���\�P��_��:Y��d�7��"'��SUv�)(�6�Kq;S�����7�3H�B9��kMT��� @�߁dJO°H����R��4�iJ��ş�;�' �xd�i�����F7�ٳ��(�#Oz�׺i!������4n���[B���EZ9���]�9N�7m�Z�;2��GU8<����� +n�e	��� ��K��Q3�u~)17��<*�v:;��]�m�b���=�>��_ki�ɰ_�5E��~�o���tzf��o�H�~,�	�7�\�I�� 僈��1�w�X8����2��xH���e(e�������7��4��<a�v㧧��b�i<�Bzh��q{��"�fjl�%4#���R���A������7���GB@H��RF��?�TFy�h�@(���V�A�M2sF�p�2����Q������Bw[���aI��nMT���Z #����O���E5��z����۞�ZTTg�+�d��i��N���@&�4/za������Y���l�J��A��ǻ�&>.,f+���$�	o&}����h\3k/0*Q�����eZ3G��sʶ�ߑ��sM�7+�D�w�ɠ5fea�Iv΂t�-�(X����A�Z�\��8Ժ��T����ޑ�X:��C<���}6z
`�y�W'�i�6�w<EH�(����ԙ3�vK)��e�u�V%G��<�cS��w�r`���aS���J�-������B-BN9������@����{�%.v:z�!09��2�u$`%i�K2f���Ú!��Ku t#��"��U<������ �.Y;l_���45�y�׊��5CƎi����I�H�֥1ŀ�^��w��|������7D�~������ V����`����O̭+����l �;��s�լ�9w7&F���N5k��{#\�"��C*n"S�78Q,�����4�L��;^l�L�ˏw^ fqn·���Ql�Ɋd��B���H� �
d�	���OvM�	c�i0p��6��ma��� C�~�,��(Y<�A(��Aotw��4��@����!���$�h�1���-��U���d�>~1�eWYq<�a�)Rh��.����;�����"~Z�TU�A��Tϑ�O܈�1v�{r��P*�]�^��X�S݆��1zm�����O��-�����v�N�n�;̞�Yo�\a`��|n��fr�����\���T�G�l�\:|��6;Q�k��a������"����¾���E�%&�N��My�����&ɖ���0��2��
��%�Lk@b�K�Am�tg��7q�K��3Z�u�&��+��*���Fh��6sS��\����Mzw�o�����H�u�R~N�����ߔk��.�����wV?>��AF)��fL��Ɵ�m!���4���������8R�H��c�ڝ�Ѳ��+N�X�"B恬[
nix�K�N���Jxb�M�dp?�,78����\�eJ�o�y����9,��$/���`�m�R:��M����3}�6z�?��4��6��kqK�t?��Y����1�I�q^T+wя�M���*��
:�'�Pٸ�f�]����с�寗0�<PHV�!c����uy��(���ҹeqJ����HA\�C���*~�/��S�����aם5V�oH��e��-�����q0�$|Q8t��ΞnA��gH<�cMQ�3�]o��<)6�8}Oq��.s=�>��S�=E���]�R�'��w��!�ܴ�T��0Nr��� ��;��Y����R������R���!<9���S4��BN�q�EZ�#Zkۘ�ue���f����cBԛ���M�����3y�^�Zpż�*�J���,y/�'\0�y�o��;]�E5:啳�KDM�k�=P����צK{bɽ{Ee�\~OO���-�y�u��p�7�is������
Kj~|�a��W�T>n&I��]��b�F���+�"Z�������z��&v@��̬K��K��|��"�gg8�f���.ju�l����M�y����+����c�-��H�T^u�k��r����)70+Ź��F�e?e�Lj M+���/g�O?��3�?�F���8�yp���p4+�8`j�꣱i�x�����l��ݳjN���21�(�[#��X$��ʖ�	T4CWgS���	q��0M�>RLE����M~T����x`�j�̐^��.�p�=�#�Õ���B�c��lf��sp�[�:�ͥ��u�
pk$���1�B�b�C���e.	# B�&]��/[T|���(����G�W�M��������x��q5��p;�� �D�2��I���&퉐�R�L���?F	������Q%z��ESb�^�I�k�#�ت�/B���z#��ׅ~���
��(ff�ٚ����W���Φ�:�W�y�a���FG��1e�Hey����,�N�n���䂗�[�����?��op͛(��S��-�'��#@ �y�M�m�I���T2$-�#~��>���Ye�&�^���[h��vD�3��2c�!�dط�i�f;��?��*~�c�]��@#�&��)�r�a�ҡ�QܺR�ظCS:�wt��rf�̟�2�2t/����[$�6��J_�b6^m&�#O��� �N�O�9q����J�����}]6
���8�=z�'��h1<H;���*�)�~��Qs��Ѹ��^�%6��4p��2z^k��y�΀<y�o�R[�4�$c��4��+�ۨ�ք�{�:��)E�R�/��� ��ܽI�K+�9�v�;\�����'�89�m��%�'Ȯe��e�" }�sXL��T6n�`Wk8�p���:})zq@�����,���=`k��rV#�4��`�h�13�N2��
;E����Zr7{��*�0��q�����b�����8��:�|I�O��w�#�� �"�
�2?���#��nI!T�/|�L]�,�uoc	��s��³���٨)����񯔘���!����*�U�?j�쵝���9Xu�`���Z_,��.��L1v ;3�0�KW1�5D�\�|rGh���\e�>��܂��dFm�¢,���KB��V����umeO�.�B��`Co�D��Y���mR,�W�;~��E�~*l�cD����]H�_�	"���p_w�0L��;?"�������+��T�p�*i�;-����G���ME��>���L�������݇D'h����2(0�5���;>�H:�F�cf,E�07]�!�l�J��Va�	���A}'8w>S����lro������`��J֠����*��>�B�'����+F�1����M���:9��HU^X�D��hքd�E	�p��m�1d��4:�T�,�fX]<�\,�D���^�#�f���xh̛֥m��ޗŮ���:�y�O���sZ͆(�N�"����kc��Y�%궟f/�̜�!����8q���gA}f��Cg/�?+?h�7��^@[�������O-�)��AM?�o� �seM4I��m���B�q�ԣ�TF����F!>Gh�o��q�����(�xX��j:k���"@�x�
q��`�AI-iF~�%O!���Ey4�d������+���a޿G=�4*@n2�M�7���NmS+�t����V��#��1��f`����G��lʶ*�&�͓��z��٣��c�=�)����B5q�������>�/ˎ�;�0wB��1��"f�'��f�@�ݪ���Z�M��:+�Cg�H�I�t�kGT��Ԋ�7�?�#�ب�
`�4%J:�$Hg����8)jH�wA�䘒Rܝ������I��"�듴�{n98�C�:�s�O���Q�6�� ���tdw����_�4 ?�ą�҇ѝ�8�Y�����i[J���.�t��2�s�-��y��]ͺ�����5lw
�ӧDus2���k�te�e|!`D2Y�db�h�j���8����V��6�1p{�6K�h��2�)5ǩq��� ЙUnx*us�0�8N\;�`d��(�o@�#��B���t�] �����*�����M��!md1q۰�7wYҐ�+�;����G�������pi�y-�$%UY��W���,=Z�U���@q'?�5& ��M�����u�zUhD�A�s7g�j�y~4�1��͒�[���$�3g�(t�v7�Ҥ�IRMT����CT|0��h�c$]��f^��L=!J�1�x{�&P��$�ۈy�'���U�.u�n1lX'��ڒ�j=�g�Y.���sCk'P�����G�qZ<�M0�`X�lBGp�������h�+W���E<�e��J��A�UO�UZ���R��Н=�.��Š̘j����g�lC�,���s>�rGJt��q���lQ������y�臭@e�_�7�k�(u5뇂-�2�?����W��fC���gcD�_.�(%�+��Q�Q�`qz-�	)�c0��;��WʊC��p����{n� ӿϓɑ��h�Wk��}�.?������	��NN\N��9o�Vs+����o
��IV��=����V�G�Sy�+���҃�vC���?S�����	��|L7�gZZ[��u�%�p:���{�IL?el�ܴ�AC\�����\��h��[��v����-_��f�0r�w�N�c�~�!���u�ֵp�]	L�eK2�OK&���.?k��,0��,�c}!�=�8����o�P����M��K���o��M�u � l�S7Ba�.z�֫�{�MpL�j��Ί�@�,6�Ղ
�En���D*O8W�tq&�[J*�w�[��)�!	��+�k� (:篗H��G��a&� �-R�N��z��4��*ĳ���!���pfΧ��{�߼�L�䡅F����+��9�9���T��l׽GzDj���^1X'�O����2��ށ���h﬜g(���k�����6��$^5����W_&5�L�f17����!��Ա��+Q?}���߿�.9V�7+0�}?����zV���3�ă�>T�#�s�D:����Dȡ�~�ͬ�sw�M�&�Qt����bþͻ�Y�
�eߵJ3O1z*?�z�.�o;_��3x�=0,�Ȋ �֛��~����&��>�c�Q�}�
Rk��K~ <��cג+��o���;in,���;�&��SZ���D�(�Q��X��^��M>5�n�PF���yC�`��/⏿e�Ҩ��<x�0��C�(_�o7	�i~�V[���\F��9eR!�����m#�ܔH)�u�&���=Yb�&��7��=�Y,q��n�^+xU����bP�%��"B��.,ܬ��gj��� }�EK`�Ȭez������ѷe�����3���d>���8��'&8�mޏ�L]��`�=��g2P�(m�� �cIRP�.�{��/ю�%sn�,�%C�$�����4=���,6��5/�Zs�?d9���o�Ng�r�-�p�5�"��9��	��]O�E�c�Rg�����K���*3�sRTO9����aΔE��y���y$K��c>��S�[�=V�I$�5Wf݂��V� �Y��I���J�,hp��V�鯭��C������̙{�i�h�t̖�v�W�C%6����_�]��n����0� c�O�L�6��|L���f�P���n�\}���	ʃ[�#�߄ӓGt�D��DS��Gaw�������D��=a@.]����^�z�r/;�ϋ#F&m����-���@�{�E���I��)���CB�ؑ�w�:�U�(yPƏI��G���S���}�F������!O�dtpІR��:�bh#(	���ҽI8X�2ĄM�d���<�յʹk\l4���b���T�<Hm��<� �&K�gf���e�JIe�y��� ������'�N��y���Bd�E��*�S4�/G,vq�e�
��`�`�h�"g�@N��1��-������;���fu��3�Q ݢ�8���LpAa�U�PuQ��x��
�L;i]$�.�s��^O���t=F���y��飵��ײ��=Zh�8���j^%d���t)ȍ`=69��z�m��8,�l�Gp�I��\i�U�o*t��� ;3�QM��z N�A_�V�O�M�/�������:�0��{�E�8<j��Yw��(%��^AWh(�y淮#�S	�Y�k%1�Rlo�ʫ��ؾ�͸�?hB�@�����?��}���C�/
�p���$�栘�{Ó}�f�I��_
 �������\��ЦPsSؼi;�pm��B�{��QH����N��J�y�D_�o!	�0a�8�ɚ�r`-���υ_�x׵v�8W����8���������߻���ṟY�9G�gD��Vn���/�G}C 4�n�9V���wN-~�I��Ǔj~c��nT�:9��MGa�}6��݌�$���S���������k(P�0bR��uq��Q�Z�%Z�������"5$l�2c�GV8]���L�8!� �����l�0���V'I��}�1ͱ�Y������Q[w�r��U7�x���V�5=�����j�<~�DH>WN��"Ғ�א�;����K,O�s{�*y��OJ��@��:���jn(A%�(�] 4���F���
����B� =��{
i#�<P%c��T�&|M-lK�L"X+����t�E[r\%��d6�!Ә*�
MI)���2E.ۉ�'-�~g�K����S�,ߜ�5ęx��O*�\��Q:�td�,#U�z����Dr*�B��%e��(VE����Z�B�}�H#��NH�<�\k�� 0v.�e�'�����񎞕Y���S5x>=7�Hw	)J��q�t��^�ٜf�&QGt\�: ��o�\HipPo��l�H2�x�"�fp�����gǹ���#2�Σ�A�(Y�K~3|�"�{�J�җ�[8趿���b~�w�Y(����'s٥�j���
�!����Ҳ�U����` wgږ�T�	,0N��X�o�I�q�K5���,�#�D�`.�,�m���59�^?������7��@�n5��8T��r*���t �;�8��4��0#;@��;�����yD(�h�����n�8Tʾ��A��lҒ7:	L:��n��4�@I&R��_��@���?N I����p��9�;$����h;��yr`7QD5�,6=����s�G��?BT�=��D�b[��r'$}OEA��� j��\VM�Wa5r]����g��n��g�D֯���Th��ȭ�U���▄�w�c��	Q�?�-݃�G|ÓD_��I���v��,a�W%����dcK��H�KxϵG2��*]_��`6+���ܙʯU�D�l*9i�H�k��ڄ�����E�ۉQ�)U@>��<~�kx��^y�]�]Y�'qX����uk��eb�AFVy�^,!@1���S{���;�9������'�˯����u���	@��	��-��A{�8�a�]�c
 oS�|ص����/p��X' �TT��3�E�����*Ԗ����^Ș�����||V��$ ��]�a����]kWk�ۻ���dPlcwg��V`f�,sqF�p��9�P@�o���K��@�k��Xd�I��]-£�+��Ln\5V"��;�w�}��ꯇM����&��� ����.{�U�0�g���v��.��t�$JH-��*k�c�	<�?p��/�����ڒ���\bSCf0�u}E3k��5���d��aHcKE��i�.x���#��ݥ�M��*4]�F�J�<�*���3�k%S��ϐ��S��{�������%z�<b�H���ǖpc��,>��6�T �(c��> J(�Rk��[�n�;',�e�a5,�v�3{��9��
��P�m}�D[V6Z�� �8�W�d��QZL�������靫p�v��ӝYg�!�2Ǔ�1*<^��c� 	a��9������hi�pQ�	�r����Cf�O�l�Xgz�$;1+㫙�4�����v5�#�wy�jܖ��~(i�����b���b�B8AK�I��9��0��\��I0�������n��C��M��=��G6bM��������/���}.�r�Gď�"&�����K�%�uF�����k��=֢�dL��XNٹ�ي��Ѐm��S����d�Z5z*���L|��N����D�&�ª�M�:]��E���?0|��ʙ
#ۋ��e�M�d����\��'���)�^SK.8��A�*@4`�u7I��ƍ�i�"�k<�*������<���w�ل�CХ�/��F?0��B`��� U����[~����u�:������$�n=�����P��M`�8O)&���]#�W>��Z�ԁ��V��B��3 $>$gF(�V,� ��};P�`l��U'e�����9J?ڃ����ExQ���Zwf��[���Q�(�`qɥ���>DM�lh�j�6�0��Y�w�sbYM��89�R�t�p6W.�UO���-m���n��k�ߖ�^�V(�
�l�>�_�@����?�	��oI�h�z�����0F�� ��Q���Z�jn[6�l]
`wƼ�M`�� �+N��(o��;�_$1s�E����B�W�$*�'��]���\w��y��2wؿ��6M���n`b֫S�Zw�ϋs�8TRϏ6����^�?=�ɦss�$��/j z���ʌ��o�qx&^�\4!�a%����<��nu|�z}J����[F��\�ၱ�D%O������K����b��ߏ<\/O^�(*g����x�/ԫ��'������d����X�@���'�.��PV��+���<,յ��vcf���m�y� V(��Y����x9�;�� ��g���	j�G� V$k&�&Ts?��KE�޴��^��)���M�����-��+�7�|��ݫ2�}��$��ZĲ�\%9Ii��C�e�V�s�h}Ϸ�ff���V����9-)2�0#��4�A�~��蜍��0��
���:�H)ˍ'ҝ�����uN�rE*MY��ñ�ܗ��o���G�m��{��^�ⲑ�v�ڵ,^Ix��g�b9r9,1�Zs����GF�LG~C;���)n"�ϙ��0�(3@q��`�|X�'t�}J����4����2!=�g1/@ȩ��w/�*�>4�r�[yC�`>�W�^:f;G�%�+:n"^2����QXằ�S�mm̨��Hl�*�c�54"��<׸�V	_M!鹻�B��kF��h�	�!h�%7�Nn�r� �&M��"�9 �������s`��4�]H`��c�%N�P�20�.�(Ǥ "3�?Tt@��җ�5�7���~����*�$�A����|s�f%
7�ٙnx�`�������G�n��>�C�v�/�KO>�{"�&�?���K��<�#�%�|t0��ހ�oK�{�`˱��'gQ���%{�j���:H�ՠX��?�����Hn���-�s\�N3��0���.��׮����
�w�����UG��U`���*>
���$�_hP_QTi)����"\w,�j[p�MD�)Qx>U�t����?ai���4:���	�%ȁ��-Hu���P� �U���o��E�NOPuE�⳵���#���O!����q���^.�+�k�a��l�	��W*9Ga���l������k
���~���ʏ�����
 #���#5�ղS�q˟9��x�W���52�X͗�U�늇���5v65�-Zr���"#�`�W�g�rY*~܉m|�-p��<v$vx��u��b'�T���rZ�!��}1�E���{N��4����܇����WɾDݿ)���Ƹ�� �`�r66�-��?ž@�h�Vv��kVt��Z�W�B���b3ĉ�k��2=�VR��+"sVM���ɗ�2r����ߨ6F���	�7�'��P_d��r����l�,$W�j��%}�6� f(��H9��>'�)u)�D�kC#�JP�j��Pݯ�P@��j[DR1���C
�ݧ�p���)�0*�o2ee�֒c��L�!U�P<s����1�nE�}��&Nm_w�'2�WeYb!(ͦ��c+��P-8ĽCװ�'�9l�_64"j��8�C�w� �Ä?ĭ*z��#��;���W���vb2Pr�ܠ��h����BU�Vr_`:�Y����O����bF��']NW�\��K�-E�"5��m��AG�W'�8�ȓ��ߵ��a�N�#%ۧ&Rn��3!m�dJ�*�N���B�LdMm����
�X��l%{QUԃ���$���`��ۀV�Q���F�Ҿ�9Y�@㺐���?�}b�f͊�7j�W٩v'f���$��0cIV���G=R��U�7%����i���ܺg�5P6X�Z�p9�I]/�-2��O�����:�������-��;�{��+�� ߝ2iy�y�g0��,1�nk�%���v{G����*T��[9jO�-�бD��N�p�m5���&˕�� T
P�oǸ�aI(�ӑ�/u��%xr������R]�3f�!��ކQ�|#o	�����>�]�/���L���g�<����`�"��ӆ�	��-��t԰p�o�/�x�Z��u`y�$�c�pg�
3��1�,t�� �V��߇�[<��yE�L�4?U�IR�b&�[e���:�'7�=�ro$T�c�ߤ�.8�BH�����C�`��t}��*���~A�L����Y���wdi��KHw��R�Ӿ1��T�-у�*N�~̋LPu��`X��4�͝����� ��X����"=��8����bI�-Hx����.�Vi���?���vY΃p�If2��[������P��0ב�ɧ0�e��;�h&�2��E�z���t�B�k�ke�NL�n)�[u��M|��ݻ�	�4���9`]��r�/��M~�mk�*�5�WP����}����������Z$<�]���|��^ε)�m���o�<ZO0�a�gi?�&l���-<8(k{?�nu� �c$���H	9���B�[I�~w �R�.� �&T�AF�����`K�M:�� 7WM��O3�n4���a̏�NYL�=)�է�C�]�s�+�M�)�k�鬺�Ԕ�@����*�W�Ug}��e�|OB�>��4ǹ�rB᥌�g��N�n�֛�xF��_�^�4�Ű�W�8xb�y\YY��C�'f�)f";h��b�����Mb�F���z����Q�zA��[xO�ukP� :�L��)�SJ�˗�
���uC��f�.H�
�m��hm4
4��	�at��V:�F����8;@2B��p�9i$�ߪ=� Ó��1R���a�x�[��M�T�ֲڜ
�AƠ�*�܎o�lqмV�g|��sܿm���'��1M��[za���l��x�YӎD]��Q/�\��>4�㾾$�4�J��O����tB���;S}?�.���P���مc�GϞ���fr@���ZZ�9~�%ѩݙDp+�®�aS{e�+M"�+5:!"��� -�v�7��'[`�Ze�,� 'nKc�������}���ӧ�Gk���8��uD>��������i�#Lpz�߱��DO�pZ�+ǻ��f��3�i����1̉QC���<���K���7�h+7q��}��������E�{0�;�,y7���hh�̼h��p�f���{Y�G`�XG@kt)������]
+Yd����<�U�|���eV�ǟ��~Ӭڱ��x�<k�c%���� �u߶
�3��hv��>�b��埛z��]f�e��ӹ�y�&���IT��}��3(���ͻ��G@%q�}��uƽ��O��(�e��Ux{��P�V����z�M�UX�8��ا'1䌚�^�G�ϽOl��jb�t� &�+B�[����������8�Cw-F���ײu����B1{������� �)D
$-1
RL�vȰU9`��<���Ƹ�����d�&��i�o���[rk%2���*��'|�p�d���W�9�E��������(6 ����{�>}0&��:$����`��A��q�R���b�8�0��^"Y�~J����)�9�$�.����o�����妥���2{:��.�T͌(�)�W��O���4����xɵ[��YK~�:͒��e/b��
G*F!�A����.7�N���̅�X�U��,[~E����8X�2�[��H��x���kG�CnTT��8n:L#�Ț�욱��=L�+�-�m�ޙBOS�0I��M��pN9hߠ����ٿB�J�>��*T`�x��R=4|y�Iu��I��?��}����/1�����	������]ҏ��~�hB���l��@�.:�|�:ү��5{�	_�'�0����RN��Q�^���@�>�1��/-M��BrA�%S�/��:nw�K�`��R�U�����Z?��\X���.���D�iٵ�Y_9z������'����DH�{�h�t� ��M\���Ⱥ �}��g����6�>w�;6��oV;���pAV$�Q񖽚p�m>]a��������S}��ڐ�Ƕ���3����]��EE�=�^F-��$lEF5���_�+i�f��M��I�9�e�%-�[��r��
n�)rU�Q��� `M�;J��%^�Z�wW��Z�ʭ<���uR��.�m����p��n��������݊��T�cb��d�gPdU<��8_�n̯.y
�ˏ�2�y+�<͚�1�}֟.�{ꥀX�j_2=l\C"��lh��Gu��@c?�X�/�ɸ���vQ�����O��(�L#6�QǨ�.�t�O�7>��X�ۏK�7�R%1�(I��x�hup�H"��k���O���L=>�L>�t"�p��`�ؕEN5��$ ���y�Y��*�ʮ��֡И�>��^sTX�Y���y�!n�~Tl�j_h��T�y�yRuKe������(�˝}��ԫ���p�Q3#4�nӲT��_��a-�=�I��n�w(s:��h Y���c�A*�M؞Zk��D��ey�HJx�&�Y���C/2i�%���[^G��la@""�C
�s��j �)YQ�wg^<��F�9�;T��u��N��"����m��Z���ε6�_�z#P�P6�'1�8�tK�@�Y�:�c�dn|�^��	�K��5�\KG��W��j�.]����io{���:�A��&d<����#iR�z��A0�e^Q���ٕ�a�K4o��nI�w+�9���6���4�.�"�G�l"�tsy�4=.�V^ MJ1<�~A8fW��f���3D��������	�bXǽ�M�,�h��Foli�-��֐��4�Z��EA._����u%�Z>;���������-�� �D�'3(�-�}�d�#�7���:�0[�t���@#�^�~i��`���ja7��dz%nq#&<�\⒈��lY���RC��� ,e����h|��k��δf��x�K��ٌ�Q��tMf�aJS$?�k�����Nd�7���	#<���1�\I*�1C�W�����E^���|j�:�/��>�"��4�� �Z��(���B��\�h�t\�d�E`�
�yN^�2����*R�6�� baq�9/N�\�jqzn!�1j�b�7:lT�d;�N�S��&�6קÐd �wJu���k�G��(���9,�6��?K�逸�(�3ɢ3t~݄�b �8�,�����M���d-�c����Өqd1�DW(�BPӗ����չ���Z�eJ�l_�%��@���w�� 6��ʞG��2�BB��j�&C2�FUOw�*4<�n����?��@�;Txs�p!r�eT�-5k[��+�S�����=ѹ��8�������J{`	0�ڀ�z�ެ�L3/T�
<,a�pCY�#.�B�����QA	R����"B ���be�* �%���s\~��.&�W.��6��^��� ��P��uD7�n��&��7�m�F+��C����.��cq�څ��hA�����2��:�����#ln�E���M�ˡb��1O	#5oe��>}ٻ0���>��&r��~>t)S��O��2ل�r�b톞d#.���2 q�2�YM�e���K?���,	��C������
�xrwR��Y�����nl�̚~	�4�h�*��k�y�M����X.eP�پ�g�{%���M�:;0�l ����[�o�2�dMqEw�R�/aKx��P�O;@'�#Qf�<9��������h�Ep__�8E�9�)��-9m�����ߝD#�������]��n�ڥ��{���V����x�.z���DI�a�,�s�����bY����́%ZB+��h[�ap���\̚�A�
�T/����Gj���1�_��F�Q�G��-�wm��V��#��[N.��u$Y���R9M��aw@������p߫�$�BD�����0���+L4��Ȝ��a���I,K�wSSi� M��KtK��%5�'���J��Ii��ǥ�<��:N�1Os��hw�!j��Xq�+I����
)���>w�9$�q|{p˫ّ�8s�DKhg,@��a��[���I��������C{'�Y�}$�~y%V���j~�ZU�6�'N@6�����>�ϻ^h0�Ю�ȎK�jG�WLHmi�S~h�~��q��?	C��wC@�3�}l��4�i'�'�q�p���EVYm�`��`	���q����e~�*�YW�m�!(���{Ý����*�e�&[{�	�4l��x=p P�i��s.�����:�U�;?-T	ϤT�u�gf:)�6F`��JG��E�6k1�Z�=�7芼�!�(����Bxg��#���$J��W�˧���R��U�R�P5�r��A��0*��|�Л�>�F���=�N����;����\T����0o�AAVo+�� ʼ\��h?�$|nG>�-2u	�����ʪy���� ���H2�:��w���-�#1������x�|��
�ٗ�\��O��f��o��(�����9��cj�~䶠f�����y�V@�ܧ�u�GcE��Dq+��j��4J�gf݁�l�A-��h�|`�,~���<�L��>�+��O�|,�0�7�z���t�(<ٞ�jp1w}U����,Po;���M�����ԑ��L��#Ni
;��V����| �5��6��^-�|l\8��C=ؽ�Vj5f�ɂ	n5>O�э �1׆ZrX1h���G�
f��W���y�+�\�\����!�4�1ŝm|�:W���-��}�$h�����n�Ҥ�a��o;��4x�_Iө&8�Qv�͹u:!�oSv�t�;V&���}����΁����.��wM(RPm�_S���R�C�:���S�|�=��N2y�:q^��v�'�φӻb���ơ�>7����Y�XO �U��ۄAv
ȐR��~����D�wۖ���d�^����+'D�V��]����!Gٻ'_���;}Iv�!x/ :p�!if������QO�#�����<si+X�1)}pܘ���ǳP���a�	�qV���f�w���2��n�ـ��cNH���-8�	�U�#��J��\t,�O��k�-;���1�s
ٳ�,I�xq�SC�� D}�J�	��L�7<RHc��kXd���FF��������Iv��M�
vT{Y�w�#�:��{���!;�͞o�˝l�r ��g�X-�V!:�S�>=
��k_�jk䞷�2�:œv���rS\4����co�ּ����x3vsZ��<.�L�x���½A�y��dX2������y�g���c����BVOQ	C��Iy�^�2���7!�hPOM�]�0� Bб��e�"R�/@���5$~{Y3�ى�����LŔ�ޣPS�]���`5�ʠ3zQ���F%�^��u�Rw!/S����0��oC@QRHރ���x���f�)��v}� Zҍ�>F�^�j)�� \��`��r^~���	�b�3�$OP�3UP�D��X�f(_���$z�_�!�s��,����t���xSf4Sj�$U~&�n�{���{��#3������ L3�%��V�di?�ټ�ۏ����2���^s@�W1abÍF�z��|@����������W����x[
��M������& �{��Z�$$1��C��a19�;�_��:�D�v�b}�hz(�����G9Y^��y�X_+_:}�k��ݑ��S�܋�O�`���݂1a�!�#`�h��~Q�z����O�la�Qz~��U1�Ӛt��Guߘr���$�%z�1�2�7J��[映0�z"�S�����7y6��o	��� [����3�/m�+R�ce3�c���[:r�/�*�a{�!<�@��7SVa:0�l��u���l>���(��g2
��lt�2$�~���Xf-J���BJ�H�l4�#u��?�Y�P���2�x[�!�M����m�<j�!�O�ݽ� ɼ��+�gO�]n^-��d�9gUjq���Sc}����[{� }.}T�=�S���p��P�^�T����\=�������,[�F{vtЮ��ϊnj|Z��Y����r��U,bJ֔��P��X�.���Y�,�]�*�.0Zb�dXR���f4���ל�9�H��������wa0�(X�4	� �a�ɛ#BF%)�->��!:L
�����^,�#�;(3�n��W�.��1:߅���k���knkB���@q	��U
�ߗX��'CF�"b�v:���t�����n'Y]�[tU�'�b�{;��ZS����ؒ��oca���&�S��;���Zs�00�'����K�D���t��#����C���j�@G���ZP��D���f������*�A��{��0K�>���]�I?1���IOajJ�^�|���c9�w��#¥=�<mD��܄�T����
�=����z}���g�G?I��Z��d�S},�B�G��~�i��;M'\�U�g[!n��5d�_�~ㄤ
�Xs���ͯ����i���o�|�I�<��y�!هB�s��u@�{Q��(X��S0�Y��E���:�PL�Z!�(�f�j��Ƶ�h<<-Zl�A�Δ���3T����?=�&��n5�I2L�=.2ވw�]�=��n�:�V�1	P����W#p[R�
zE4G{h��*yh�n�F����u؀��xy��fw%����cja6�'9��SZ��s1�îA�/ͱ&FC۠��Cta\(��-e4�=����Pd��Ɣ"	��<�qp !W)R�E�G��@��hȗ{�d~0Xq^������"�È��7K� ��ӛٗcذ����cG47А6��G7��C1�ʇޡuFp�7��d[٥���F�2���,�թj�-QNZ��W��^D�D�O�E��� {�H�o��F^��+Q{H����@�"$���_2�i�F	t������z����6�PTr��!k���O'w� ����3 g�y떉�����z$���b-V��0��JC��d��H'4��DK8-��M�1����[H����֤�Z\��*�"��xi�Z���7��}h>޵�9y���h�����ڇن��W�ǀ��u�ɧ�� ��V-�kcH��/(�a9S�K!��D#���W�ӊ����Tg�	��g���7J�I�U12ґ��eN�ʼ�M��g�68�;H6�e�v�Sl��s�,��1o�J5�6d�X��n���f��uċ#�����d{���*�^�Ҫ~o�|ʮ��v���Ĩ�z����	W�ԣ�YN�sW�Y����/@�i@N�.�g2d�<��9m؝(Z4���.ک����Q�m�Y��Lk �N��'�_��{w�
E��:�rA2�����Ѓ/K������F	�oc8VL��Zf�ƃ*�L"�������|��y�O��n���U,�@^h��\e'"(J��y�"B{D�DЮ��qk��� [L-Z6�H�`�Vѹs[�����Xr�[e�W�>�	�wL5��������pi�æ����'~�1Qѱšcv'��`{�[L0��N�i��lz	8r�G�ae�+����QVga9�ݍ`�_NP��D2e�=��i@�&��y��{i�-���u���sj��+��j�5-(�EzB�5I��N"���XK��5��N�e�ñC��"D2.� m�*=�N�X�齰����U1w'�=a/�6Z�Ô��7!h�xi�g�h��Ѧ"�|h���4p���ࠅD|ã;��gb�?n%�$��Ӓ�y��.���ºSЦfOh���uʆ�[���^ztE����\%-��x����Z����ܪZ���;B0	L�*+`��W�ȟ#�ؔ��H��ve�w��gL ��&����ߌf���yъ@�4����]�ZS��Cr�5�G���~�W�1���{<��r��oTB��g����m��e����"��ϙΚ�M��>�'�uv.iME��:ᴨ5 ?�Τַ�,�S�����}�u��B��]�/>;��AMG���V�^y~c}¿�r(0 m�Ǘ��4�w�R&��l�~��a��wv�M��fYĖDxmK	^q$�t�9c��ΣjfB�/X�n�R�F;(��V�s��p�p��'��R/�F���b?
)t/�O�r+���<_�̺s�G��S������j�!��Qy�7�50�.�����ά��F�v۴)�aOW=T����m`GB�;v�XT�Ǵy�ܖa��m��$W�%�Z�Va����S�`�V_#���4���uU�;n�<���3���s�!�7�K�A5X�E�gR�ʢ�Ъn�4��-P�l�zW������̺�0�ٻY� ��_�U���F�??��n��f&�wF�m �T��	j�M�����⋁��:���Թɉ�V��/�P��\���Ai���v��B�F��@}��eg^��J���>mR�]����@3�%P�C��7�FK��A*�D���G���GBW�m��I\!2gV�a=]�Ǡ'�L�t��
R���XDz�`L�3 ,Wӂ(�,\�tw�ھ�)��q��Pts0�>���#�\	��.<�So��4	"A2�J�u�WvV��Ъ*�Y�o��>)<|��'H�5���^��fo�A��K�>�K��j^�7g����`���u�{<\����c��Nd�>I�i�=���G�.�<8K�B���%�5�<�gw�_=Ir���n�s~?����+��>63�q+�@	�z����7����� ����=�Ce$�q�ͼ��+V�^"m���Zr�=�)�p�I�t��`����Z]�������@6��5pҞ���7��H��e�''�:�HD��cR��ɸ�H,+����4�2�d-T�����p���:�z��ʉj�]AO\����v��ۓ��9\)=Y3���Y{�hv,��I��`ο#:�eVQh
�xV�4�֘��y��a�C��X[�
f�H�f�����	�g�!q��_�<�=�ːƇ�h����S�nR~�{#�0Ct���m!L,PNacA��w��t��%��C�]e%l���iD�x��:�W}�M��T
j��y�P��[xU�z���\7t����70H�l�.j�ch�Á:�{�Ŋ�D����m?���/2�}!w��	'�w
��t2�ޤem5�vӥg�
��h��\$���s8ݺ��"Y�;Vľ�/+$ڡ�G��ZNY��ɷ�D��}Z���%�I'����m�{��c4�}+4f�7ʍђm.�C��~dkg�;�K��<诪}Ϊ �-���e���m{_]��8g�tK6���"���0N�=��6Z�_��2M�-�ٰ��?�~H�ey��P1$�.ʟ�!��4��0���x7�Km�!��ݔI��N}o��і�K���{IuW���㌫A�����l��n�-?��љ�~�{]琕�6c�w���&4����T�&�F�h��gM$�o@��اq���%H��/�R���h�=9b.]�3f�o�x0f�1=x��n�����s]UO��	X��K��̎X�̉5�����u��
�v�S�|�������j9�svAe��Aj�c֨)_�)�2�,ṏˁka$t�S�_4��}�k��\1n���g���,
?+t#�ҋ߽%�}H���>󃨎�{Ch�kV'�W���	 @�r�L��C��V�C�~�Mx䶧r-�u���.�=\��a,���A�
��I���y@ �Sx��V�=u�q"^w�V��؟�VZv���[E�r��-�C��]�LdSzx�,������{a;3���:���S>��w|�����vl� ����6wc�_����溫�vj
1%ԭ�#�efV�;��D;��Czeg������1F3�jF���wQ^�Y�y�2��bEe?wb���mכ��Z���-F�o�Ұ��CU� ����xKe�ua��ϕ�����Ϛ6tP�J�9�}�hW�����|�O@��/}��Ȉ}�q&���"ӓY�g�&�"=�b��)��E�wҕ��0�����6�����r ��
��l���8@@��O�c]�x��;T�aJ�}�W�����ռ[����U� ۦfN�3�U�|�J��m�Կ p�*�����[-M�K��[�1�ڽ�.�ly�`�,��n���H���h�L���6,c�c���N�# �R�`�,�8���+�+�2�i��d�����b!M�ܮ��O>���	�� �C6�z���A����P1~p����~7�~��-�R�9L��P���X�=���?��.A�QT=�|s�ϭ�_��y/��4��D|D^;?oV_@kI��mF�oyn��dB;M���0!Lvz�{�#���	�G�[�~�C��#�B��s��6N��Ө�����Z���V}�/���f�TkɅI����uHp���|�J�v�&f��M�L	�d��f|O��e���9.)���P/l��o�F�7��o��0j��T=Px=�:������}�7�c�ꪯcϘ��f��� �M���!�.Ϫ(���.ʾy�������cT(A��E�|p�U# L"�D%y�����8���5����Mni-�m�`��=�%r��f�78����:2���ꔝܴ��%vnk^Ǧ}�=r��"Ɛ��Oh�����}~)�1h����8�/�^qzxЍ-_S{�+mӬ�s�w^^����]�g����������@Q� K�Ć�hy.Pa7���jiʟR~�aznJ[K�F���o����"�(�M&uٞ�����l�o��FΛa�,���n
����fmq��
�58#��t|8�h8�W����H��L��=6H}���u)�� /�]9P�����|��o���aKQ��9�
�0�̃�)�Lѣ�:�ˈOq)F��{j�*��KT����s���eRBo�p�|�5�I��\�b��`���KC�>`i�=U���t�2׾�~�O�i���AU���y~B��1t�@\[�Wr���ƓQ�g�yV���<ΉY ���}������`�b߇�\,�O�[�3�}��F��xԄ7�ys�B5�|�N��Ȗ C<��1�NX����'|�-�@��J�@�Z�1�tF+ܧ���,�U'��py6=�^�S#ޮ>��ڭ����q�7�&"�7�d! �F��z���F@O:W��f���A��"�I���� i�:G��q��o�&��� ����6�1��[�0N:�B��1Ɣd�Lq��;�'x��p���x�}»v�ur�´�Ak�z�#9�M��6>�I�8�V�����]\��˓1B6���GQ�[����{�LOM����)����S�<ҏ��dt���?�s��P�D,���O�ï-z����+�e�$I?�A�Z��b�S�
j�$��\@ߕ�B�"�oF�6YEW�~uaU�=Y�qʩ�Նq��1�^����q���OЪ.%8���V��x�&NUJ�ic,�d�("�	XY�*�B���1�Zz��f�`#��lf!�GJR�5t���Gu��C�q�_���~z��@�ۇu����U���ðX��?��,=��ȋ�O�"�
g����Vi�j�Y52�C��VU�.���'1P��~ЕH>K?8�m��+*2���VE/��~{���Hc�ݑ��2� >nomY�og�O��������лn��u���M��ŋ����w����7p����W7���.-��"qG�ƅ��R8�U��o���G������K��?f)Y�μ����p:c'���{
t�#���8�����DnK=�]��0�P��?�
�$`h����5*{R:��Bu?a;�r-��m��h��W�<fe�����w~R�cj�S/��	bH�7]�����}(��
�w�D�^^b5�q��+�����4v��I��+�eN����bӼnݗ�)����1ߞ�yՁD�dWVD5�~��Г?���&�b7�q���K�ƸBP	3+��Wˠ�1��X�s�m`m���;
B��[��E�4�d��q�����\�oZ�IS�ґ�Z��iצ�n�"��ؗ��Ǎrݎ��`�X�7�T�터H��LX0���Y]��8�o�O���E^�c�T����2rZ& �Ղ�����7Z�Quz�m+t��ό�]Fld��|�Y_7zZ��P��SKc�*��֎5���DWm�w!�A�	h6��CN;�]i�.�/jn�2 iCD���:�l�F������.��y4�oS�"�G�D?l���:Ń���ߝ�����]�g}K]���~���2|��7 'J�e��t{kD�y��Y�)�T�5�P���p�V��n��䶌L������Y�@G���M���H��6�b�q�/�3����e@t�C�|�?���s�Z�i��N�{)A��l!Y-Km�&����~�b�&rMg�.I �K���#�7j`��m59��S	"J������7��!壘ک�S��#-��rF6���}F�מ|��tԾb�3�G���mY�N�_Ƿfks���+�w�m��
~0;�Z�`Q�ְ�������{��}ഴTwbߋ���a��}���A��8�/�ڡ��5���?�Su�%� ����E,�4uS�M�(�dK���� ^ҏ�<��<�z���4�Du���5J������b�w��pC��rq[����?��`��a(�����v��H�#4��5��X�<�N�Y��8aKr**4"di�0�C��lX��r;b�,�M���;��b����}j*�:z[����Ӻ��8,zfj���u�R�����>hFj�x�I���-g��V?{ I+_��1�X����*}��9��c�oY?nD�'�yʢ�vu��l�`|�Ux��%&bm)2H]�l�^����jA�����9}Z�8*��c�=/S�\���?�h@nl�9�8q����g��v�9��TRH�bi]���R5�^�%���a=���ǎ��k`}�@�J�"�#E�4J��:�HT��^ E�=�κC�U�Yx2Pc�ɋ��w��miu.y�`y�/Ϝ��82�V��������n�Մ�:�;�C�����W���B7�V���"$�fT,-% ��[�K�gsU���f��]&��R�8�/7X�z�vӾ���,�L鉅�]�9(��H^�	�����=R`�?���v�V�þ�������p�Q	{�\�`;���yc�L��:9�~٫{8��mKϚ��9H�>
�li<i���i�'��h�y�����o{�Z�3s�v����\5��b�Q�uO�B�#fL�Ctm��>\�4���ً�,.���pFx+2��|��"��5e�X�����A����AK>'y�C��������:x�f/D)��C+=ƻ�nY�&�_
�����M;b@`��>v�C��&
,_H�����f^ ��c��M���v���ٳ}5��63`!7�A���n�8���e�6�id��$����P]<��:���c�n
�ӝ |��R �}Y���R1ޢ!yI���=۠r���k��v��g5����u�!޺;�<L30@�OYT?�H�(�>�u�k�J�SR8�\,K~����=D�J�C�
��7o�&���	L������]{'�3�w��B$�eOC��]d]
���P�LȯB���AGÙ]_f�!cb���Yc���{��r搛0b'Z�jzkMܒ�碸� �K������1�����%|-���ʃSp+ �\E�PWS�j�U��1	<��m�e�_Q|9�������NZ����n�R+����g��1�D6!�G���ج���id� g���^'HX�6J��+a��Iu���&���r΀/j��]C���C�va<=x��]S�`�%���l��PRt�#G�,�闫�I����d����m|<����[,�s�k����{�0g�v;}v�g�Z����t���h���y1(�#����{�l�[���������g������葴h+D�f��:~��d��
K���ad�v}�D��2o��Lmgum���Tr� Gh�-I ge�)�3X���Dc]�]�ħ*�QE�;"�����M��_�BŦ,�rCdVt��d�%sӄk���r���Ed��$-�k�e��fV��3��j�f$&��ܓ�E�W�j��;EUpf�C�,U��F_ b��^�pn�?}B���D<J�C���br��ڲ+C]���}�-	� ��k_�08R��5�OԢ4�x�a;�c��H��3קĢ�%Z 0'��nX��ݦxa���$W�ⵖn(Rp�c�_��$OE�:
A!����V�U�"f�5��Ƴ��㗩���ccf(F?%��Z�N<�����Tl�|��p��5�-cUf��q;��w���xAf�]��k�c�D�ސ�~�1�bX z�d��~G礚9 �o�m@A�� t���n\�l��qM��ƊD�-� fF)V懴Ҝ�2��w���oo��ݣ�O����+�x�l���b}/��R��:&���o�(�o·��h�~5͋�i�`O�N2��_��-�2I��@-������R�|��{K�$�
�/��k�����҆]�1�fHV&o?���k����_.\��W@��	`�R�X@�<z�$���������SR4<��k�� ��T
��]�2����P��k��,:��U����$�-,:��M�=y[���p���y�u�9Nh�˅�����P�	\t�,�|�Յ���)ggYg��/Ix�%6�g��VL>�屑I��H�jY�֬���QH^�[I@��(ȟ�hN6�d{�F!C� b=�CƧr?G�c{XY��#P�� E�ғ��@m��~���jJL��o�rD�~�h{&A�� �%�O��~TCry��l����&:vU�j'��<�,^���AU�_r�����8���/Q1�B��	�QK�<�7�u�y�p-��RVM42¼�,kX�� f����~��-���{�3��2�&g7���4y���X�Ux��c���eDHo�Y"'�ڍ�=y�@�!^	��ڿͤ����V���i��V�f��pp�;)�*^�J�g��\�N�ϫ�����r�H�T��PS)�t��ߙ+�v�����r9 y2Q��u�3���=�L���:��k�c#�{���\/�c�P,2�����a�0��T�F���s!N�tΏ����L��V8.��k��ɇ�$	�2K>Ċb�0��v$S�kd.�o�G���l�t'��tq��3�Y-�5��{CŞ+�ڒak�W�𮛴��Ӄ���匔���Z��]Z#Ը=�?G묘�~6��5�������9e܁"@���dɄ�_�\�ks�� 9I\P��}c2��e�z�=JGlQPO��u��pM`�)NPp/
�*Y�ܥtۈq ~
S �A]A��J=jn��Z�7�IF�4;<^��6u0`����y������#��k�mg�&��O��R��+��"R	��\�c#�������i'u����l�y��C�`U�;=wV1N;�0��tf�"#�N�s�Ƕ�uGR���������Ąz�vM}�*���'�R��N�UrÜ|�����P�҅�jQ�H]�5P�27ꕠLY�z)�zQY�J���`���c�A:�z禪cu�g+���=����%.�#���Q{��W�����^�C��4�W=;��PyШi�QL猸���1�r��i&
�.��N��$Y��(�b��������&t�CCg���[E�0�6Ђ����I�����z����C���)��*�O��G�SǋK��LȄ� �B	�JoC��.0�R����ra�5����B�f�<�&IhF�B��2�y��b�!������ƿ��t8{)�һw!�t�'��$W��4�ou_� {wWs�:S����A��l�}u�W�meQrVd��9^n��Hc0�#V?&.$��<Fqǃ��ԉ��^�Ƶx�:�V��&f!�b����g�9��3Kf=���"���1HlAX�<��i�V2PڏD)���'�i��JTSu��]$��ѫz���L�~�Z׶���1��E'e��>���U�6�h��o=�A�a��L�#
�^:E}�[�Co;��T3���'�h[�CҳD,h1�Ϻ��jܮ�q��m��ئ�:/?�۴v�t&�t{k'�qצt��OE&w��_��$~$k,�$y�Ψ/���b�8����F���z�̥ǘ��h�j"X�(i�Ac��(y�-FMx���?� O�e����64���ڭy��xp�tD�b�&�R�@bb��%&��>m����$p�K���>��3LK�*�{*D�=��v�h�.����Z|{�I��T�&)��ԍ��s�i%�ı��Ǚ���4���Am�[�Y����g0��gj�E�&��i��/�����(��0�.�aS,\�Cs�'�U�n��z�?�"�X��Iŀ��9E�-_b�N&x�o7ر����c{,�զD�O9��l��� 3����|\��d3� ��FA�T�v��E=	#��lz�=�|����H����7z֏9?�l�����Yv�xP3�&Ӑ�3����_�.�|PN˨�7�ϒ���F}�tD|s;rxv�S5T�t������8R����~�x�&�0���ʐ:�� ���e�~TT�s�^1����fP�6��g!r�6����n������֫	�ci��W�������u`��5���.I����O��ؠ���>�g�s�df���%�]N�OƔ�w��/�.�)�Ѐ�y��GAi,Zm�<e<�$�Cg�F7��ܤ��s�������-������|!)4�:	���*}>-M�N�{�{��tpۙ0p�T5m��θ'o���� �7�Ԭ�*TJ���l+�_��CxV���s1���$6(�7EWl�)�de��`�˞J�X鶇���1yf���V���pjKY��:VM�^� r��@��EN#�1�Aa��>~\�M��\���C�>��Lj,؃�ϤS	m� �H�{�"�mFx;��)�p�t�2	����*�X��~���~�1	�N#�U%��)�3�׀�"2<��Cw����L
IX:kV�ʺ�=I��		�"����N�|���՚(V_�g�ږ�T0���G�(�/�� ��zs�3�p�&��J}�������@������� �Z�{�Ia9=���?
ܦ�	K^M%ꗩJ�a��"v~Z�Dp^�g�P�����j�D��/VQ��t�����劍|P���QH�R/ 9�V/zIW��_wz�26B��&���#GU9�M�j���^�nr1�צ�|��n��S})��G] �ՏO�Z`��|�J�í����f�"|�)�HQ\�R����;%���3��b]y'z/&�|ƛ�������+<�������7����w���/�)��y˛����;6�yy7T�Ɋ��G���
%�F��[��x�]T18�4�Wg�׿N���N��\1��֡��i[�������+ԉ�z�Y;O�qn��)OVZs����J��y1��v�֕Le�l�Ӛ@/ڝ�~�>Z�;��1n�����W!�_�9v������D��������i� ��^e�wӔ���D�s�~@��)壹�~B"eã��Y3�a�A����G��7~�C���h�i��g��w�D���<�� o'\������=�)n/�-��A���<i����}�\ﻓ���X�-:g9�!��/�Y-Ԫ������J��L\?"��#�_u�^�����`����!Q�D�x��O���pnu�_���ٹ��f�X��~�աG��d7"�A4d4��*����L$���4#����g �x��(���ٳck�a!� X�N��X�`����ǂ!n�C/R\Y�# �)ѧ�١�#����<asC��N�&js-�r�9	�6uY�%JT��V� VOD���#�(V��p@阁l�4������1l�Ȏ	�����r�����{�@4�iP@�����"ޗwY�O���}��p�E񧐙o�ك��*��g?_�ד��9K��6a^R�x6~��#tF��{Y-��O]�Y����k�Y�:�gk�\X���_��J��Qt���e�
|��BY��.�(�����kn�73�a�C����`���HЯ���tt�s-���\��HrN�u����7[�o�B�L�^\���OXU{U��*1� ŮN��Bh����2䆒.5����&��]ǹ;�!c�γ����@�F�D��Mǖ�AZbf����^ ] ���LRiP��#Z���R!w'>�SN0˘���}0塎n����)�;^��\�&99�6��c��k����P;
��F���`����-[ŝ�]� �׭�=�U�I��ђ?7`�\�,�
S����>n�o�au���6�k0�����x��'��`fzx��.��/�f/�ߑ��k��2al����K-��l4+O�"�x�Y���Sr�����E�TN咑��uǅD����o`'8�}�c6��E��BV ��_}�E$G��`ty)��/`�T�W4�sgX�3T��JOxIA�\�T�-Mi�2�Ba�:͈�-}��Wy����Ă_�U��M�nG�_�R�H�:�2�'�a�X�NG�˞B�G��
��G�[iCvjQ�Wο܇(H��Wi}���f�CdX�5�~�]��EgaQuS+��M�uТ��0�y����w�Z'.����uE�z恎�?ٞ��Eo�ٙ�ZxH��p6`-6��D��٥�s������4.���|z��BC �qJ2+������4[��V�W���/��qvm�P�+lr���9�W�$��1$��)�s��l��ITN�����/ڀm�L�{{w�~���1�]t-S�q��}��P�!��Ħt�����;���zA�N�x���-�Vx�X��.%3� �6���yu'��ڝ*�B��=�p���7߷~�l�)y7[����g�sH�x�1�f]\�" ��;
���5����*��e��O>��o��o�-��J�#�M0�v�%��:�]�7��7�.��`1���L+-]f�i0�:/�Vnh2+L���-I��'h�����z��)��PǼ��y���9H����$j�k�ɜc*C��K�C�ţ�)}1�_��p*�D�0�R�
	�p�W|�$M��� �~e���*�r1P�F$�
��O�)��15G%6���e�Y�M���n��@�#ne���bt�� e0�~�o(8�r�~�f�Pp��BqγY^&]3��;�}��`�¡���װ����?�?�+��%�y �f�?�u}B����F*
�=���2��7����������1,һ��G^�d��B+_��C�ta"ym�u]bb�n�2�C~ǋ�଀�gi�L��o>f� �Kr�n���ia���jg.(��Þ?r ���q	� 4Oy��Z�!�g�$<]�8N��õ��/���V	H�K�U�_K����c�ϙ��5%��c�$4������@�͐ә�O�+FTj�־X�a��E�_�<�	�DW_�4��̈�)�n<8��]�P�J�4��b(F31�	sЕ�<=��+��XU݇0��Q��k����i����T��	h(u7�Ϭ�n����S�Ǌ��������D�$Y��S�@�o��:j�v����#�xu�!kn��I�ԃ �"��h�Q��$O�!�V���K��B�XģY	j*j$�6��>�d�dxS}�D=��J��BhUW�ڮ�(☳�}�뱄�$���n�u�����<����w̇�\r^і�d���f0n�}�f*h6�.����|��K<)�KP:����NG�v�n�*Σ���{��m�ny8�E��/Ya����r��$Q�:���doI����nû��=@��_5yH��Z/���eR���
*;=�gM��� �d*�4Ö�_c$P ��|�5Q]3¡q���ih��ot	��۹'��)��;�[`����c�y�B[4�*��6�\�Pe:���߸����r)8>I3r�h�b�9����@���9;��f����@��R?{��s�k
=��YJ�𾮅a����P���\d�~��{,�����-C%W�-�Mp�z��cK�� g�����UQdl�Z!���^&�Aj�BMs�
+f����#ҧ��FR����W��ĪA\Ղ�,F� 	�^�<�n:2�{Ә4?��,ѩ$��]�$���f�����&�xn
"h���XN!� C��X�2���|�^�Jk/��ӭ�AW�h�oY�j��3�k��m:����3K�)��O=`������"$��!���+��U�D�Hp+4/t�l�nk��5Q�5�G�6tcx������-�x?S��z ���d7s ���)�m(Lcg�Kn3)����4�=�C $&q["�ā�����xd�Q�ڵ���j5��.݇��yU�6ay){��|i��Bk0r{Y5C�PqEJu�p#��C�����(���lQ(j�����C��a��}�d��q4'���Z��7XD�gQ��O�vX��\�E��2�(���ɾ	<f���\^�8#��e����:�`��44���P�!����1�Zۀ����fC������q�_5�&Zs4AKUڿ<S�������6
�;����a�WW�<��5��N�0���i���ڏ�(3�������G�}��c �,~�4�o�����4��>�v]<����s �x�A����݋�H/D����I��}(D��͢
3!*�W���.�!r���\�W�? ��B��p���9�����j�B�
�Pe��|h��T�O~�z�<�!4c�v_Kx�+�i_��\����|�Z�5��0fsۍHNw�u���u�M��_h���lw�
���Bx���M�J�
�PeuS�.2�¦���cX$�؂�F��;��}�����?��'��v����{i���W�5R"�L�9���QѶ��6ΤսW׫I��t�9�ff��~���/?]<Y��2+�,�owYC-#�a�FB�7ۊs���3�?��v�`׃k�
�����&��I�(��#�A�د�_V.o�oLƇ?N6D����Ⱦ�O	5�A�%�r��횎����*�,��{-��uf\V��W<����M�]d�fa�YϰSX
0F
�w����\�w��a��U���ySΗ��_;O�0��hP[��>�Z��gq�U�[S"4.��/ߝS�`և�K�&F�^�c�u��RP�ĤO���Ӎ��!�ɭ�}�ˏ~�V:0�C�C�.�r6����c�><���Cr����?�a ș��t������5����`c����L�{ӈg��<o$��<3p��:��(�`�<T�Wkb�	>mS���;�pdC��j���X�P	���{V���*x��^?�{����>��BB|Zj�XQ�և9��E�4�D���8��Իa�Q�djj���Y�R!��j���j~7��ȗa�!�ѯ% �εW!�ydk��#�9���ϭ¢/��'�5����M���I��e."����Pe�5�6 d�[�Gy�͌�f`��A��?�
ީ�1�l�s���&&����e���j��3Ι?�q1�7,�Qs�_@H����%2�Xo�H��T׵�o��A�4ċ�/�ʬ���m�X-���3���Y`(�U۠p:_���gͤ�b�~�wͽ��I�s�&���7`q���~��z}4����
E:�r���1�i�S��H�O��'�H�2V#p��2Â�0�S`1�J�EM�J��y�b�6�K�i+@p�s��8,f���!�����Vh��a'�;3��]t/�~[�ZW;�gN���f
"�����4��F���B�����M|�Z"�ò����uَ�<�d��tx
����SBNԃ��YEF���՝I��~�%3h�/58���z�|&�2�vF+;����x�Ͽ��?o!48q��E���t�f�V��{ώ,�ç���'~:�t�^��_�͡�j ��i"�i.�Lы$>ԫ��n3 ��2�?rTc���SD�N�(B=�� 5F-�i���+Ӯ	�o���*q�e��|��\ªV����>-}�ކL����@F5N��"'�v����p��'�����Dx��	7�|��}C�� V�Ld��Jj�6��c�)).-R0��etk�P�u�t�R�\_9P?rS��JɅ����i�����ɗ*��i�N:��jx
�ÿ��EFvwpI1�</%!`ω��c$��%��>h��ED�����u���zt����
�i��(�`(�?Z�#�%
������3-	���WxaP|�i��J����Y��+i��^�m�Yo��?��dvT~�p�{;͚�Rթ����PF�)4��:��M��b�^�:�)C���M�T��8����p�:$�o�]�ü>��\��\�sD�� ��pU��D`�`m�� B�XT�R�����׾�'���κ�G�yC?�����4�בs��V�D�p6�늅w^_X�lx�����H�c�pDZ}�y�Gg����� ���R̟��T!kO�\���#���Ȧ<܂��5�l;����ɘ_�փ~���ژw�Qb��%U�c��붬�f ��z�@z��脡]���i�K�iVm�W�k����OU1���E��s㓍����K��yi��e��Ҙ�\�z6�����wlI����ul20`\d�|;{�X��%�X �/�~�L.Ĺ��VZ�y�9��o��#���#�S��R�ָU��� ���L��-��i+��!D%�Xɹ������Oѵc�,
�����RH���B�ࢮ �F��-ܬ�wb� *6����hzi��nn�O�q�h��K�7�{�����U��]U��_cyM&�J�y"�k�n�����+��� ڨҖ��z����/���o5��݈t�Yb���o��6��MwCK�63���`�����$�8�ٔVIѯ��|k/t�,*0iWw	N�[�hPF��N,!W�}̢���YV�sWn���8��Q/�~1��a4�q3*	f����p���}d�w*X �%�5U����_�N�/�~��b&�� �S�`4��pG����9�i�����+�E�3%�m����TUճ�?�]�rC`Qd��*V��3�:���W��	���Ew���g��J�B2l��o6uQ�w�.D��$,1�.�N��I�;��T5�;��7� �H�ۭ�B@_���Rj��sa��;��1{��AZ$�V������F�ף.PH�*�ʄK6gY��$R?�����P�/�"fV��T$�ݖ�F�=O��g2��x�:�D�.��,|(Օ���M���G<��o,�����_{`m����v=� eb^���4�Rs����I�|�\�]�ƈ��em�<�<�C�D*�?���-�c�8�r�^�ZL��õLiȿ!�w*}tݧ0�.�p�e�(g6��08�ɫ�S��)ޞNVnӿ�/h:ϒb�L��&&n�6u��R� ;��S��#���zZ�d���0���oՎ�#��a��n�sfKVQ�{d������S�$N�c�Fwi��x��~o�ҥ��~n���G�#"mL��L�3�K��N��܌��뀺�^0!M��@� 8x��Y�ib���H�I��߄��Y���z�:IWj��	'Y�|���	��z�)s_q)�+����&�H��X�'�i�9��n
˃�6�bz� j�L��ʣ��'�_�R$���~�h'��bC��,���2-0G14��~��\_��XƄ.����v�z���
�L��-u)���e	��}QG�	:F'ӈ�^Y~��y������10l�*j���a��L ���K	S����V��H��/�
8��p��t,*eG�n0�Rn@�EpH�qMē�Y���V��AW�u�۹�h4x8	��u��,�Kq��7�t>�31M�=���֏�Wg��q�ٮQ�;�$�@X�Aj�Nz��ţ�Z�H\����\٣���u�ȋ������.ణ�6SbiD>�]�����ӿ}Б�aH���gfM�kN��+mQB,f��v���5�
��\�Zȫ�VO0���1�|N�W�Ca��� �m$V#�����z��䘳��vk��4O>㧐�O�Kϐ������{C����W <�KN)S���bWfwK��%�&�����q��j����ѿ=]L�F+XNA�1�A�V8���D�px�,�x��(6���]H䳡�Fĕ`����FM�F��[,�:ꫀ�t��ֶ�e��y'���
��p���k�'��oN��z"��" Ͻ�-�I��T'�
˿uM��Mc�ԅ�n��[�[f�q��4q��@���U��?K���y/��A8�g�+ӵ�*%Z�����l#CI��$���U����?�fl$�s��K��S��l��5��s/��/?���l�1np^B�y�����{rw&���~j�z��3�W�Q)@ko�{#�����d�7�?F��_� ����������6io�`|%�W�{9��!{�Ce��0��UG��ԣ�?�7��ߩ�����U���w�e~-�Y��ǯ�&�� ����&�~�&3©	��JklH�k�6�(}H�է�acC+�A3o0Jq�f!�H_����-�v!��\x�CLY�e��V5�L��ό��J*ųf-�^���D�qe������u0i���ץ����4��ò�ʱ���	�m>8�h�M�|�bQ�S��F��|��l���E.$~ l��������s�G�uW(M����)ʡ\v�ʊ,����x�ŋ"*��j���k��+IրpB�=..��um 	�j>�c���e��9�<x�c��/A��/QY�W8-�+T����gxw����F%'"�>��ǡ9Ş��ef��-�p��SJ��%�46`A'�ZZ�?C�-�2n�ũ��X�����S�5�4Rڮ7��d��{2�� �+x�d��L�D42nR �e�%�̡���b
@�S�`�T��ģN��	aj3)�����ƿ�%!��X�h�5_���џ����DjAh��eT j��
�Mz'��CN�~LY��*s�PB�{��$��{�<Y�D�*������qmG�i��l"�\����pO9_�'ݒ��� N}�;��G�&j�7���r�h�v�k7�䉶��2�b���NG x�Ñ%�q�[�|�?o�y&�?���<j�SM#y7𭼰gJz����XSߵ:W�!���`���˝(�V6�^���O��>Z��'�<���P�Vu7ٜʔ��Д\��o���.���R��װ�+������>�1��˒��,u�X,��#��I��`����+�_���&+ߔ�v��y3��$�E�Iig�1���1yd��-v6HU��|�P�Sk`�'�D3���\r��/�*�r���E�cV"a��
ݑ�j�
�?��-2�M�W��`��k�G�����l������7P�����SJ�:_ލ��6�9Q0�b�֦+1=��W��vo�>bV�?.�l�:�i�>������,xwg�A�'������o��#$ϝPgp%��4@f�&F�u����NۭO�i~��5ap4ߟ��\����S[%�|A�����ku���������v���� ڝzP28���R^M�����bĒ�V4�@��~KAرl7&�b\AK1��4�H*~�=�',P3�I`B(��^��O����t�:;�����3U�"[=><#�_�����܄B8At���Aтlxzޕ1�Rz]������t��I1��K֏��4V|O��Ȃ��e�|U~ˈ��rc�[)O�Z1�x�=�S^�
��+n�u~v��]N6����{��{��D��r���r�j�1>-����%��,��ј�0G͞���)�k��7��i��OI',�M޿�:m��)�K	:ke�Zm�ǫ\�&S�8�gNт��9Zc3�n{z�?�6ji<�B�`��!����G���qێ�`V�OW��Lq���J㿪�/�ç?�l��F:ɘ���e(�~kxB7�U=C�ῪZ#KȂ��m$�8����t.�O��0����I2V��޼e+Vͅ��8��\�#\O����WS��D��J��uE���h٥"��Z��N�ѶԬ`ؙ 
~e�Ѩl|d�4����(9���]-W�>� �<��~�N������'-�z[�&��������n������!C-m��c8�^�/�nv�R] NьX9Q�74�]3�pD��D}�39~�
���Xj�V{�ؓ���fX�!*�cƫ�r6Fm;����֬�s5�Y/A�Z)z���{w�Gd}��n*W�R�U�S�p�;ڊ��5@�����U�GP[^o_H������B��\}�Ghf�N^xs�r�Nhf}#I��3��}ab�(�o�?�����.�j�}���"��%7���Iά���Cw���=µh<I�D��D_����Q��i�7�َ�1���h.H`���nT�T)lMYŕ��.��u�D�d�!�s����a-/���}��U�o%�J%2+�G.:�"�=$]��w� ��q�H�6�?H�0�'�������- h���^�I�Lh��%�:��辖 ��#&V2նf]ߔ~��؆�9-����Bؙ#���@��Y޴��O$��z�e������\��;#�	o�ѵ�1p���/
���i�Y���ь��ށQ��ߝ�͠8���`p
6�vZ���Ć�I��A���}�;�E�1�G{��Ve������b\�R��A�����E� ]���Dy���~�
7+��r��~�N������q�fd|S���7�On B���k`�4��J���:!�*��	� ���.��9�W�r�����6K�	1����`t�^���P}��o.E�^Ԟ-�t	�7d��U����W)��f�3�`t�M'Wޱ��G��;�}1*#�]���i�ux?ȐI��T�x<a���8,L�[��_Y����x�������� M��;^V1��z6+܅'��j�%&sU�s��s�Ł��^a�Ȁ������Jǯ"ӄ�f7��l�I,�`��Q�Vô��-� �O�0<}���,�R�������*����=�,�8/�s+�D���="�oO�Ə(��{�M�5B��(j�l�4R-�]��x�T�؊�� &�çA��W~�c�|�[���	)�f�s8u �If�QB�C3�a/�ں.����ju����7����GXA#5�ƿ���g@7M	���J�|wt�oϬʸ�K�J2	�Ɣ4붋Qp4����e=2퟼}�M��#u�]�t!Rn��y�[���E��L; eꕫ�ȵ29�Èhӗ��+���<�+^z�F:��<pG�=��&ȥ�Bؓ��;�D�Ab*_�ч'��μ�����,HDewh���TLi:�34����[�L&O
<p.�0T�e�I'.�t?<EQ���6`7K����ԣ1摜�%���*F�~���U4�F�i7o� k����Fv6[ܪ��N���-�M�%���n�7,���Q�q�Xߺ�@��RV���jwO%�t
����M��#�1P%�����jy���I�]�#Zxd��	 [G5*ԅq'w���MmO�����c�����aH�̛�nS�G�;�#M���?҃��n�,�}�ҫ�6�X.�Ԑ����1(��y,�`�dwĬ#��Spg��0�K�6�4�}B�3�$�,.߱J\1ڡ�&N���V�G�����W9U�RrkxfU᫇+���'3��t`��Ⱦv�]5�;J���LeU���֖^�<��gyՖ���~d�� �)\_�_��
��	�z@Ľ�[#�1��f��j�G�,D���CO��B�jV������>���}� N8��ԧ�a����9u8�y0{�k�x�@�����@0����a,[�P��b*�8��*�"a����Ѵ0D >�\�]�T1�c�U�O��j�޻tV ���LFi�2R�Do]3k�P�˭|�qN�h�=1Ӕ�q�ܥٽ{e= 1��16������OW�[|����A��^������?���C��k�l��Ҳ���%��Y*ȯ�d0����Q�V�]��D� y�<a�W�A�b��O޲J"�U�,�O�\��)�B�$��R��ai>�!������Qp�A�zOY�S���꺊�aM~�A�x���<�'o�� �3�\ԾJ��H1~��X͑�̭��g�u�2�w��hw6n�+}��c�X�1�Wi
�y(/���5K�z��*,�3�Ƌ]	?<�>wa[3=��T��`X-�N-\~�fЕ/>0�u2��Yy��{i��^�0��ܱѠMZ�������[�2q?B��?W�{p4�T; Ԣ�Knc+�+��'F��?������a�ֵ�0���h��F�R���;5��=6H�7y�RIj��2��i�I��i��
&&�N�~���e8A\�I�;�	�${�|�I(��!���K��`Y���󁫅r(�ZHQ7 ��7��?�=QsJ�����4�����t�����ߠ+�v��N�`H����>��:�׆���_8PϤ��	%di�v�ҳ��\�oh˅t&0�[U���#/ZG0��jh�r���_�@�1d���B�����\�t�8j��ɗ�f���~�ێ��j*� 3x��"���Ԍ�-6����.Cx��	L��R��g M����w�t�0&ݶ�Q�z��� �t�|Sú��h���dO�Wy�����G��xe!��z`��]�������2�\g�L�r��JH�ҽ̌��#���"���(>��'"����X����B�� ���@?2׆4ǋ,ЉPk�H}���Q{iN��=~��˷��t�|e���C�� �ި�p}zgIř/J!; !�9D���<�X�ik����>Hm��b����-q&��	=	�S#`a`�%
�[���5�8p��:ϱ��1\�9l�!Tq׏�hC�oMuieN!+3Ux�3!ݟy�b�B�NX祱�!�߰�������y,��9x*,,K�e�d�iuJ�DU3?F��uT���1_�:d	�o��Ӡ�/X�m4�#��ؼ�8�U�דib[[��`i��8YT��W�*�z�A沣XU�DJ��֦�Q�z�?�%<���vjB^ E^ߠܵw��+޴��\���Cѿp�_m�+@�'Dk֊�:&\:��{�$�'�Q��"l�P��aՖ��g�4�H^N��,G<�����|��I�Nӆ(�3�ɶ���)В��5$tBO���x?H�4���&�_�OLH�e�r �v����s��|��]�LW3m<��S���z3b�
��������>�Z����k��b&B,ө���,���쒓9�aJ�'��˭!���uDk�vf�1����gI7�
��W't�1\���7������,Z�%h�.����l�X�&���/��*w�(�z��,Đ�k솾�츼��"�;�س(�B�K��ԡt�y]i�MNqF��>�/�--#(�r���a@��K�/���"�.>��Y��_P��뒞 �1	�ǉ�.]p�>�m���0�s�|��W	:�4�͠]��Z��<J�z��t�Df��h���Uшi�Xd�F�R�a?E\m�o<�W7�d��ԛs���{W� MT�' xJ)#_ E���c��=MA1�~f�X��`�v�}I7�pa�n�hSiA��frZ�t&R�˲��/��E��+q������=���C)��h0L����>���(j/>����.�ir�OKR\��A&������T��O���'e.��4�7��d�a��;