��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t������p$��:i7���)�^_[	�����be���K?R�	��v1���z^5K��)j�7�Q��x��1x����.��
E7����rn7����>��Y�7�%��U-p���Ԓ�D%���=�g�:+~���dV�����NMk9P�~}��p���5�P�(��e�M�G�����?�%a@���\Z�t��Z��r�Kch�_P�.;p���b^��gXw��Sk;U�|�ڨ��G���ܞ4�=����z��HA�ӓ�R'�j-���	թGFDjKr������.c��5c����J��}+���;:Np_�v�Mq\A��Po��D�J ��۵���|�2�Z��7��|ܝn��*U?�����a�q��Nw�к0�����d?�~���@
��N�P=�󵥗Ƨi�P��vv����v��:(���:K�K�^�����b3 �=��5��$���-"��2�w.C��t{a?�J&?�־���7��_��k��{F!�GB`(+$3�;&\E4[o%����[�T�}-�
���UL�!э�q~+��!р(㜈c�]����M��&��w��rT"<2*H����?��w�	7�+��P�y�i�	������t$����i�l���M=�p�j(�N�ً�K9_��W�4���R��ԕ���s&Pɷ�v~�Aˡ�A��X�e�(p�ݍ��rPs e���{�yɕ1G-	a�C�<��b�a'P,���	_����	��"!����GH�;��p�S��Y;X�s#.��Rk���k����嬭�晱���Z�z�;P��kѓ�ۯJL9�+���0��ne)}V=���̡���*mn��T1;�f��	�;�V{1W���,˳5�����O#р�|=w�%�����Ս����I��	>"%�5c�w�m1�^����е�@�{����:���
��9�,�@�|�U3<������'��|7�C��e\(��w7这r[��5N��A��ßpr�}mt�^�������;1�io&�N�<nG�@�[�h"�H �����
�ݎ͏rz~d{
τƂF�eQ����k�v�q�gw+$�)��>��3ƞ
���<��_������� �NW��3�d�:.pv����-$Y��($Z�3������R�d��.md��*�4u�G�kY�}�� H��R'�1i|<4ゴ(��$�����r�]��C��6%�x(��yy-
�y����6p�S��~L���s`~墳V���ί����2�:u|w$��̵ZMtw��L}vy�dIAPJ��6=�V�:�� �$�X���VRpJ�j⣾�i������b��L$؛����Ω�`����~uJ���8l��e������׭^Uɍ��ꐐ[_�a�T���QN��"�u���,^xO�	�JQ����I?���+����_�Pl�]�$�J&O����Y��)�[L��D�+�ž�l����/x�&�fWY���`��ϯL9Yf��qo�bU��^-g���|���AA@���N<s�y�V�/4�x#꬧��ų�Y?����\�K��߮k��JΒ+R'�SA��k���zX��o ��n�t���$�5�	L-:��Ҙ	uS��9H���;M<�����2��V�D|��ԔMp[����W��.���4#?�`��2:�x��QnZ+g�6� p�n���짘wG�?���������$x�'�%:�%�.;g��+ ��	��V��`��r�`�r�f�C�$w�Z
]���:s*�'4�q�s��+J؃ny�1u��=�?G:Eg�@�w���>K{��s �:�l<�D{��Z��J��,�>��mJ�q����X�}׷���=��``�҄�������5�����E���g�������f� �+�b����v�t�*>�(ʔK=�pc�������'T�f������p��\���	�D���i��{��m ���q����}��1�D����sR%U�m�u� r
Zp����/�#4�X_�����������,,7����S~ߌ�;^��N��པ���~�}�L��[�c��Z�zO�(ժ������D�����XL�l���&#�}a�a<V't�Q ɜ�gL{~�Ŭ��I�7[q����X��TQJt�xW�K���"۞u�`'r�� �ö)2��;l��,��ݼ���P���m�q�bW^t2��w�Ә���V�!�����]�t�ʥ1�Mt?ER>�(����flJ�u~�u�W1��
`:ub��r��-��
�~`�{jB �7 ý£7����W[��0�c 0d������n͏�[�#-46�Ѷv�O.x�"��`����i���fa�~��~��tǽ�&!o�b/־�xQM;=���8vֆyyY	P��bk�/D�6��b��n��׼���۠J�D69�t���S'K��"|�T7
璶)C�^-��2�&�ߖ��Ǝ��:�� �������y;�����Q *��碗4JBŁ�\* ��0�R=m�)��
�^�K8�GY9��z�?͒��3��/wWWG=�葤F��kv��"�������ߣ�t{��%�	��nt�����z�����l�X�Mk����0j�K�*E�ћ��/�tk@�x��k" �Ks 
7��3b5�{�?�S`5SHti�\�[U����,N�%U�L��C�(9}c�t�K�HG�| ʄg��ɛ��=�E�)?�E�lt/�7��:潒������Jywe�aJ_u�Aa�Ӄ�=K>���G+�;Aa��?R�������"d��/ s�Z�LH�0�ӄ� �?��g���5&��aR�b<M$���$��G`�.	����$������*�Y�GE�[�0��&%h�.rncz�o�ԝbb���Y���æE�I�!��"�%�.x?>����T���i�Hb��l��ٳI��fX�g�@*�L��o�E+aЭR͡��?�α�|VZ?�A&ȴk�l�4B���g�(��.e�̥Q0G�g<:��^��D{`
��d��H�T_��<�8��u_v�p��1~Nt���)�̬|���*��*�55�"�KW覇,�S]<���yK�U�E�7���fJ�޳��L�9��acͷO�!Jvo��-���L�^lJ���6e�D�.�i5�c"��W:�c"�.s܉ޗ����`\����X��SI^����BI�W�1�O)R�9�������+���j<�x��ẗ���؊�g�Ĳ�V�+�|�8ܨ�
��qA`�J�΅
�� f3�f͉Y	y�ބVna�.��L0�rF��*�o�Z�h^��v��/�\�������d�`�o�"����eR�Sv}��;bg�|�Қ��Y�PB�Y� x�~2l���F\����%��i��q�x�e̙N��#z�M�a��!y;�D��/�U໗aX�����}Ns(i����/T��G�������PV�B:�*��09��������w�u�x\XQ׏�)M���;���Nr�+���f�p�oUO��7MXHv��L����u���	�Ǽ1�D��Yf���>� ��chHU�+؀Vx��&������F�=V�Q�[�&td�t͋�_p^34���7Ź9��0������g7>S�H��R�$,y��u�:��ܴQ�1�H�Q��\�u��gџ���;��#0��Ʉ�������J}��^M�]�G���Y�-�|%(c]�s'���FgP.��2�l�!֘)�fMr&��e%�9� �^�S�a�R��ˎ�c"ˍ�6���%#ԣ߻�%M~���WM�F���L��7����~0��C���pF=d�D�dQ3�]����j�"h���E4�NLD��ò�ev�59�C�(dom��1�(@8p��!�&YW��;j'��V4�����ޫ��TM���q�Gb粃�
�>���n��J��b����C��uu|�#�㍻B
TO���Č���d��M0�/������t���6CV�N+&�C�I������
�)�������+UX�F�J'��ϕ��C��H-��!�W�r*���YL,����wyA!Kz�-/�`��5HHFl:��L�u�}1》�b���$�t
�_٨�����=����dt��+ag�bH]�g�5���eI�#^L#�կ�K4�x>�F�|��.[�us�jy���2[)s�����G��2�����c����Y����ɀ"|�y�\}�'I'��خ�HUqOb�#�r14*�
��������B�7J��d��gzH.ܽ`)���q���������% ��z>���%����C��4���A;�%�/f����/C�@��yo��J��RB3���?���@�wM���{�sO���¬Du�m��6ԩF�uhZy�&E��m��}�C	UF>���[��
�[��Q/l0��k��L�K̨�<t5h��F������xa�����T�9�q����2ζԧeW�vX:y���*�!�Oh�e�֩~n��)~F�0H�Z9���-z�uc*1�)�u"}�eSu~��S�lUU\��L��)dMG��Eg����pD����
����A�m�{�Y�μ�m����+��^��/3���WU�Lј^��s�\���ɩ�����#�F0��O�EV�����"��59�-�, �"�'kc7�G�����"�04@�^F��v����M���tJ�ڻ	��T>D\YF���w�#c�I�d�n������M#>�iLU�l�}4i<�d��tϐB��PK�~�{��á���R���O_��;Y�����<`��qG�|�OT�xU��[�:ʩ�1��*5���u{���-ɅW�]������EF�7��Qiܳ�Q�ǝ�p(Ql`T7kt�SH����!�L�#�&��_���6>=DN�T�w�J-!�M{˨�f6 �/|�Uy�kD�D�\BlE@��w᠎�ӲN�t�a��?=T����9"ď3Ci��WRj?�T]AX��f�Ɉ����J:�WZe��B,^�N���|�8�L��p<�_F8����9p&�s�Dj�\�s����S�&��3�;��'w�_������(޻�j�Z[Q<�ܰ��&YO6���!����a�ף~z�F3��F͓�C�c`IJU�������k>��a�ҮԄ3��8"�;�"j�oY���5���<8�Sb�0� �/&��+��B�/�Fm@[��i@n�m�_�O�o��֯M�2%�3@��=��~�HuiD����T�o�����g�ߓ7^j��,�%[�5ᬯP�)|� w�/�h����P�0ƖO�y؈/� ��&(�ԉR*�?�;w�r"b˱.J�w�f8V����-Vጉ)NЍf��4
��"6�� ��-�nY�x�T��mE���j�i�N���ʗ/0���1j֫H���9�(�Xptl����F�c%=��� 0:�y�<2B�zF �1}ٶo��@ �� ���Yvi�u*_t���z�~}z�{�'��"Fk�9}I�
���{�C��S<Z^g�C����U �p�/���P	��zxy��]6Ƞ�;r�ǉ!ɼ�ǜ�$�`ŕ�>E����
Pt1�~���`PL$�%R��&2�P�F�#�� iqʭg�X&(�T5G'�2u��F�$b�ީ�Ef���m�^B�m��T}@�Mb�	�����.���a��L�W�N1��b�M��҃
���h^�q�*�/l�Z]�L�û�f�j?���Ӆ?��] �P�҉���݈�U��Q�
�]\�� X�$JF@SO�*�W4��~^������\��"e����+1��*E��J&K�h�y��?Z͒v���"r!F�,�A\HQ(��۶��9-����b"GC�nj}}qg��A��c5.��9�z��j��n�l(2�nU���3~�q�v2xʎY��N����<��v���Wz�:Y��!��C*�x%��u��x#�q	K���иUȿ#�o��؝Ȯ%�BF�jN�^��?ƷF�E? ��R+��?22�|�d��ւ6��}J�hIT�jg"e�����k0��O�8X K�ɒ�F���~�A.���GsO��K�(q�F�Ǿ���4y��i��Q�|6�~fH���lؙ��S� ��c�Z��\-���z���Ay�*N p�<`=��SLm��*����6�P�Q�AJ�74��gh��pH�ơ��n��� nR(e%}&C��:���8�1��_�!�ʽ2/X�%���΍H��l��ݙ0@��l:�kC��dh
�e(Q�U�ǑV����\��:*�ݟ�KSG��{� ��u�B���\���U� 7z����Y���9�PN}�a<N�L~���{�?/Y��=�;�O*�WV٠���ѯ!�i<^����U�\���jz����?�S׋�`�CԷ�����s�ؑʗ�笽��Z����vD��Ma��Ԛ�m�������tl���	�l��?���:�Ω4��]�c;��]�K��1)z�����3?t���%�v�����@�:C�C4�f��K	j���--	��#[�>H.�n����6״��ͷ�
�~UZ6��#<J�(Ix�R�b`i|S
�_��ln�H�^\��l��D�!�F�������ЂK�Uݺ\IE1�w
�y���e�{�R~�^
+�o���]�kM�VN��R�,nv�4U��+�OsBq���*6���7�'-H�#$�F���nVx2��˵���#���RM��h!l��@F�;E܋G�#�|^�V'�W_��Q�FM�^��;��6��{
<���ef�K0��"�����`�h/[4�Y	�#/�&�9Z*A�	&t}��4(ߺ`1-]�s��P	t�q���+M�6 q�����B��P���Y[�SV��P�����p����^(�2�i�G�@m���񯴄,$rK�<eꃱ�vf�\��S.Wd�UmiB�dD2�N�:����wژ�E	��� ���>�{.�rmI����Mw`ZS<"�t=��-��"q$'�ZS|ŉ�%B'z���"[	3��׼�F[v��o�C!<L��v�?���K�Zx֔�C&ư= (���V�rj��K���[�,9g�ˠ��V�Z�X�C�iW��]��p�:�>7�hQ)�^I�ˉ���H�W=�U������S��q��9Xy<�����o�eoyӜ �{�'y� �eSq��ƒL��O-a?�iBn����7����ry�k�E�	�dCY$<��##9�O�q尕sK�r������W��qz�w� �����Q	,�K>����Gʋ�s��h�/_Α�m��p�`ϛO����N�ׁӤm�Χ�����Kb��
w�"ɾ,��c2�N�D��7�ֵ�^+��rt:Цdݱ������-�]Ez�cTx�ce���!�V}�7�-C�����034e�E��;��X�zE�qǫ8�S��72.>Q7񹱅��u.�+�
ڿ���6m٘�6��j���!Ht��ڜ� �g�$��y��X�s�E fs78p�u�w%�b)�+IBخC���Q������Ό��wx�݂��S3Փ��+,cH�/�ъ3.�M^��FO��qp���AK�L�E3'�{��e/��>�I ��i{q��BU1�iCY獇�'}�9�Imp6Pv~'��j���H*�(sk�SC��У�c$�Q���p>彘Ѩm�9!�$-N=�������8�>S�v�]��p���7�	֎���r�&�@�$�ؐ�a�^A!v�
��;z#��_��g��kM�T_ 3���y]��ms4m�K�T�r��-F���MG�o�#�2��ԔUB�hz*��A�f��U�*]���ӱ�E��|�(���m��A�>�5Na��t�F�n9�AQ/��\����#�����֍���|��ņ��Y��� {�*�4�i���?�����w�	�0����Ą����������z��.��$>�^�2;O%�r��7\K�NN�O=�n�6lP@o��k��A�9�c�!���0[m�£�mĀIw����G|$�	�">�$;�W�щ�-��U����ϣ��vq,��g�md�8�߆�}I��+�qo�!�
��>Ly�!X�v��v�ۍZl�@���~��I]�7���/�}��!�9����T��sB�Y�|�vذb��)~E��I�Qg�DB��R�(���w~DQ�-*��<ڌ&�0�/�^�('s��ѭ�˷�b��e�pd��E�_��y�Kά!}�,B�Zv���������:B~���M}b�1�⳾iY�;&1�߇14ͣ���=���q�]Y&3Ϊ�[�Yr�f��N��Z�y$��({0FX�6��?WK@�]�7<1G��T��l{�i�3�&�'QUBozr������f�,���Z�\�ƥIr�J{��&0e��밡m~H�`R�im{	��P��Yi����V�j�s���n�5u����,q��1��FPs\�s4���W�n�o��,����n��Z������C\��h���T����2�w�J�b�٫��r,y�Pp|�<|��R�k�.ܐ�W{���^��K�]m�#�#A���;~��E'*$3q���U�8L��%w�l z��DC{$hX�7�t龹i�d�0��l�|<xp2�'q[I��r�W���o<Y����J�?��C����۳Ǖ����P6�H�q�#,�ϐ�l+�
���]��)b\������C��mSy�R���ڵ%�̏�����v��� tn��Lw����m�t�v|%�X�\�� �6���(����tA�I����1q����m���t��ʌ��Oկ�
h�I��s�˩ǿ@�����8�tzD*>�0@`�P�=dᇃ�ѡ��S%�t������I�n��@M��nAe��Ӑ��Ű5�*�揪��x��� ��d���(�تg���O�je�l-���j7!�Z����H�S��Ւ��XD����ʢC�I�������~a#Y%��Dn�}�d6�jx��ua�y�3�p+��I��S���]ޖ���&lQ���M��Ƚ'N���s��gR�E2{ځ:CN�]t��O6��sn�'t����f�1zT2.��I�F����C`��t
�m�Qq��|Q eĆ��Ut�Ց}�~Y��o���uq*f����G�jg8R�8�D"W��iU_|IP�����5��[��x#� �m��	�F�֖F1��<�D��3�>Uq[/�<~i(����kk������)�����s��(k������ H��J%���m��J���b���N���˭�D�&��tbA?>=�Sݙ
��~[R��i�D�r5��ӫR�(�h��:$�	]���sQ>��Y�0�A<B��:d�i��b����6�/i0������?�4��+� �~�.�Me��*X�m��!���,6�@˝��<ñ�^�P�[)?�]5tB�����g �s�$�`�V�[t�k��!M��C�����Ua,m�I�%7 �U�t.��=�2��{(p�N�+kG�  �8���d|Z�p�7� *j�0{����x
nV׳)�͝��5����s�i�7h���j�~��}j��za��&��7m��@𠗾�ۤv	�h��eF_a���s֌(k4{��6�ޡգ}��0�[l��T�K��ߟ(�h�j�-���3��i� ��G9��8M�te���n���8�!v�	�V�K��!�
Ù���;S��Bm�0�Wkר�K��7@?�q[3G|�G��z���Ď:�*)JFB����Je�곍KL��ㄏ�O��VZ�&C�Y
S<�\0�B���v���G�-: k���\q�p����4ҁ#Ak�u���6ӵ�ٲ��Az��>�Ko¨�)��]7�:>6�
y����i�ǱOhDU�9�՝L��鼤ϐ�خ��n�g�A㩗�k�s�'�_�8u��uͅKq\�oz��y�dI�X����NfmO��M�q�y�۟xU�6j�����?��S�צi��&�C�I��ؚ�.5�lDW�e�o1Kʸ��g��A��Z��a�Z�"{p��Օ70����F���U1>����8u���(NU;"�܉������HE"�ӟ����	�CJ��䈠���䒋y�}l�P�rz'��N.Q�~0��{���E�SU�%	,���tk� мڗE�� �ݯ�L�!��2dc"�I;q�L�c٣fj���y��Y�H��U������U_R��9%��4�\�`@2
۴SG�;5ץ/�����rqX����0sy���o�/5��-��Ħ�_a�NH͂R�"h́3gsn��[�z�3|uFP�P��4���N(��b��z��+���]�ޱ�/��N��T�y=���0��d�um��a�zQ�8ȏ��v7E�����t�.��.I7�+��t��s�fo����`��)8����8�$^]z_ǥ�\V�"��cL>��HK|��A�m~�<����4 "���}������)�@��e����ѯ9D*�Y�9d�O-�.�jO� H�n�W��1Hx�/ޯO��c$��_�,	U;.hmURDFj��~m��ٷp�9�nS{2ۣ ͆^�_N���զ��=�n�}��[� ]��v�[!�� !Sc\��פ6�c�<�AMY�<������nC��y�%H���������%��_f�)U�o�m������"�gƚS{4��H:i[@t.n�Te�J(/lܮ�Om������yfn��D�4�Ȧ8�8|,@���2��řc�'��{	�C{�Ȟ�Uz����R�Dd��V+���x�F�6�O��x�:�� ��9Ȫ��<>�	\��ij�fi'�< gɊ�=_+$�~��ǻ>� �������pA�*c����f��f%SRi�1���F��4��e�5LO/*#���PdA:���L	@D�����\�*R�ӕ�,k/����zC%�i�*�n����Q�r�G�TL(�3fޒ��o1;Md
Oր�l1����
}��#��mQ�� ��ݵrx�1 �2�cL�k5�-)�^������s��	�=���,r@'�T]�B�վ�~l�*]K%�ͮV��Y�.�"G=kΫM:y�bxk[�|+�Y-��P�<�N&�ϿǃH��*8�p����y��]U��WgK?�bft�Y�^�}��B����_b�ܫ���^��fS��v�o4`�u��%��5Y�a�����Ć�r_]�����h�v������.�ި_��Uջ��E~E����'l�z�o��;x����\R9q�5�^��1!�s���"��U�2�+��BVN֛ŵ/ f��E�~Ā�t>�����w�W꿥�݃��~N�֧t�d5�"�m��1�ŝS��êjX���b�k5j:YY<�T q�����|�<�WGh"�^�Mu�o�75>�%M��o�lޔ�E��n{Ӯ�Xc��K�h�ݪA$΅��/ӥӔ��o�Z���G&���6�$3!���O�1;�=[$��M2@����t'���Ƨ��f*��(sR��rh5*���^����t�#��ۓv��(�,�ZX��b.۠�hw?�7��7]eZ��b��_�tOTY�C��Gc�Ӽ�eK@���ne�A6�4�5�E=ހ-����Oɻ.����a@�¡ѥ!�kY
��_t*��M2�dA�j�QMs)�̋�G66*F�,焤��qa�m"�N��`����Wˁ��f�GN��%�~5Ǽ�~e-+��:.�A�{o}�6wWv奊Rl�8Đ!��|#���\��A���P�R��R@ŷ�>�1q����Hl���;�E֦��� ��� ��\�yG��R��ѽ:m��d�w�P�4�:*�	��ޯ���8�Qm�?�~�AmJF*b/kVU��/�L�S+&p)�Ǣ<�&�bRd��%n.����?q�nr�%Í?���E��S����c�r�!y�#A�m-ڗ�{V�U��X�":��3RFt�r���Zg&��0j�_7��@�������M(X��n��t��g'Z~������xE<���<�N�cI@��ǝ0�?��+{;Ѻ����N�@t7ZֵryU���kB�$�f��I]3���f��Hm��W�ķ^\)��9�~����p���� ��=�XC�v�?r@ǃ�C&D�?�����{d&
Y���~}�@���֢{DY�4�z5u��<�밨c?�^��+o�Ɓ �x��e��n�xd[㵗�c�<?r�K��D����fI��Vq�C���ɼ�Q;����Zqr�o�t��!_�?��F���'���Y_4Y�f��e�U.���_���!�\O4~V��J�W�%�*j�X�K�S��gO�,w���X��T�u��1�\��9)�>a]�O!e�y�ULt�;/~��ְz�aX{��Hg�{V`m�|��A ��J��I�}c���A�ֆ���8�Fv3�~��LY�S��>����^+��+=���]���+HՓk+�ϱ>��4��?8c����Є���Y�U��$����	D!͒I��j݄,�}yq��j��C�y�R�nZ:�!6�� ��?��t��=v ��͜<��p� ��o��W9c�J�^%�o�Y{@yw��Ӓ��fW�)�3j�`0\%�b�Hͦ�C��:
~\�_���ij"� x��2��+F�	m��.��K%�,�)"�k���F��c<*���\I0��>g5��I5e����QCT��)��>�����{��C�z�kʘv
�ݬO5$�;�\��c0��[������[-s��S��EԨ�&���MY>F){�=��d��L��u��M�h�u	[-�S
Z�5T����H�݋��8&/�2d����F�^>#��TyCE�9I��$��?�Ew 0�-㟡��F�VjD��4MZ��ׄ���jK��(�<5h/�!"J��c<�i�c���������^���3_RT��\͌�D��G��%��;N8g ��y��t$��Z'G�x�����a�r�\C8���\d�y�C��+ͽs:��tڡS�^��aň���͐�zwg����L8a��>rV�:���H�~5�yq�T8PKx� ��E��Z0_*GxP4=�c�
�$�ᇯ+}�<��[@es�p�� �q�:���7c`~{nDQjZy�z	�����7L������>���8�� �&�I��׋n��ʉ�Ĺ��-���|��E����l��0Ё��@����\��� �ҥ��4*8��!��mC���:V��P{�}���Ʒw�U�?�2���O�$�:�Ү�T��&ә�W�r{२�k�|ǿ�[�,��m�9�#�����K�Κ +ȓ��zG���(4��M��:�D��A�"������O�:=r�_�q�竔�1G��K_}��lKg��Tز}�3�R�*!8�D7uٙ�W�0�7	�D/�C�B�X�?َ�a�Af-�X��Kڒ�ϋ�f�So�VD��g�9jeV��)�.��G΃a��@�0���6'�IA�z�XIh��SY�_G[����f�sղVj��9^���q�Ah,M�娈� 	u��sh�s8R ��iZ�� #̤��>kT�M�c�j�Ѓ!�ت0�шM-��t��,�f�Y�b"��c}�W.?���?R[��'�"h��á�����)~g��U�3�A���i������L��@<+(�J������}zWBn�9�j�ة%͟���j\W�,r�Q��1��I�w��Z�����q���#�-5L�.q�L;8D�cu�H9slE�e^��AwW^��5�#�ji������٠�8q}w:�����T]ʛ����A��W��Ԉ��_�J�2*o'}Q@�>�����[F�J	*t�n��:Q���b�d%?����`��*T{�2m�� ��·�ڴ%�I�>��n.���y�
5n�ح{Sa�c�dA��������<g��D��z`QFӨ9�Х�ރ}�u�v���B=U���7�F��n�l��k�iQp�i��� `���ݸ/>K�m[{X��G!���� 7�����5�-4؆Ș��VBf� �l�$�Y@�v
�7�q!�[�`d��3����fut����(%����Ar����0� x�/Z���׵I<X	o��7Gb\?1�\�Ѵ����>��x���wS�|&��Y��q++t㱮�ƁˉWW��8@�_�3�#4,��u(��!DZ#_�r���*���`�W���Ƒߕ��ԩ�}}�*-yC��EC�l�gQZ*��SܛC� O+"��.ڴ�����Y[��(��	����I�O�Q����Nr�����ԧT\�\������ݠWT�kj�OD����Ed'��Qïh}.q���X�b�`�U2�P�#kd�L���Q+!b	�N��������<� ~Ҁ�ހ��p�C�F�nО��CY�Q�:Y�)ȣc\VUc!�;����U��kw,b�P��wr�GwH��ׇS���`��H`�WLVn��I�\<e��&��5?��37<����cXM0�ҪJM2�� �ܾo;��=)�6��w�Doe������v.�K��1�@���6���0��:��+3��B��݈,��+�s�!�&��U^^i:p��|�EH}n+&Cq�G�'�G��^@��	[������$�.���v���K	6VD�\�1�j����X��e��5�Q7ܑ0I�a�>Qށ˲��c)�&Z/�VZ����E?cݪ񠅇w�=�oӪ�0��6;�0�gL�O�荵���]�yc���^��5�F�����H(���+��e
���/����6�0^�U!���!K�^P�����m!�TƆ�
�P<
�G�(��EYn��"�8!_���������z%\@*�	�w����kT_/S;���������qj�/<*�t:ҟ3%%��I�Z���,�<�B�ݦ8�q.�$���C�j��� (T�rNĩj�����H\�kh�.���,�M�� �A76�ݔ���Î�QV�ǧ�G,(p�y��FD��+9e��P������BZ���rZJ���4W��R;:|9_)���0�c�QIk��e��իiE���?b#Z��YL��P��o���G%��9�\�q�f���P�;��Z�D��mjJ�pF&�Ul��*mt�RUԀ��ft���J%��<�����`��,=��ʉ�p]m�_��$|���&�ڡ����g߅���Z�4�S��NB�#W~a�{�p��p �R��6�6�o|�[�K;M�g�8D��b�v3�T���n/�F���A�W�.���W˱7n�P��<|kVm�5L0�d�6.��Y甶�t�g�_x�$��e�g>��æ�T)^&�/=-�!��q����_��G�����BW��jcu#s�g7�n�5Qr� ��2�F�s�ldŴ�B���o��Svl)x՟�d6�G߁��;�r�. 6�ć��b�>�k �ً������|/�G?�1мx�)�$��H��N���P�T8��1Z,־�z�Q�ނ:�y��i�ULN����N�]�{�����G�%��V9"5?-`* �#���#F)�O��c�"O
�gir�s�fj8S�J_��+�Bj!����m`��5��Fʚ"�bP���ؖ�C���4�aXS}�Sc-"FC�􏴼y�	�3*&'��ͦ��_4';�SR�[Ȕ����\��uy`n主Xo�(��|��J�]��x� f�� m	��O��c�&��+s�Of�B��g_׏�6�R�=s����ào3��9�j�v���b�ꉌ$#5U,��� SR��e��]�j%��m��$��=ٻ�8h�/�b��fK0�(<��1�����
2`Z��O�o����Z-�����j%��,g�4�c�IkuV!�7?�������})c
�'q�Tp؊�Z./�$<8[��Ĭ[i�KO�ΖdB�|�
;!?�
�j�K�!FJvo%E�����ּ���Ĳ��nPmy��w��Ѳ ��{}����M��B����h�P�:��Gw��5S4���[��BP7��x�-벋n�S���j�C	� F��M���B��
Jv�YJN6�l� �#��ߑ�%��(��9zi 1+�Sm��1ĥ5`�93��B�mu��dVh+�U}�4���i_!��V\G\�*��\��k��&�Z+������ɒD6���k���,=t�e���+i�8����h��w����|�B#1kO�y�3@�����ߕ}�J��ԝO�}|cc?Zl�`��g"[L�v�A�p=w��#:���7jv�����SM�q+�A�
;貪���2P�c�W�Ew�����v���hl�z����M�q>��G�������c�%��@�jx	B����KX�T��ʳ���]�c���=$7"TE����珿���`�&E�l���D���Mk*��߃��@��ړ�0h�!QuPk�� оS�;}Y�N����u��m�[�,L���|��E�fyADo�5��j�����������?���Z�"Io;]�ekŘ����x�s���}��n�cy���մ�S��O9=.�a�؞$�dH/��y�ʌ��T��υ\D��Ԃ���t�9>M�� ��L2oj[�0?e���0�Ms��=��LѲ�������\J����r��%ut���a���a��2;N�C;���5�.��3�jh7e�0L�q2�K#i9����̲��ū���G��x�k�3�p{)OL~fR�L3��O������H\9��#�(�q��2�k�e� ݳ�����S�m)�C��rʽ?�����@g����VyijJ=�|G2�,�eὰ�/I�}��h���sK�"ȳ�V����)7��Ч`[��_��^a&��� 疏w�N��>�аG����t h�$��ƈ*M�:����G�șbu3�,���ǯL�0��m���F&8��D���q"�9ј�i� �1F�9>�r 7��]����f��s8�G����3�x�+R-��̀�����݌d��_�@����A�M���h�{�%e��_�j�c�����}	�����*�h�av��b��9�c%�vm�V��G�&U�]c��7�3��g:���aa��X�Q�0-��_���V���wy�c�z����vM�;����ۏiP�0�
|_�c��0LH�h�(��F�9��8���^Z�Ҥē8��2�r�|�[tn���밭-�x�,#�g]
Ad����,���ÓD���9�hY�=��i��`э~{�fL�(]�j���'��V�M�[\܏�Xi��±��)����7,h)\�{��b@�'`���`y~S�Z�U;O�F�X�x�_�AY�ZJ蛠���9h�9�`���VڂA#G#�DH0��d����RaX��|g�N��CF��*��s\M����GAcS�8�'Rg^�*�h6U�p���Ĳ72�e����"�J��+���=c���N4�jze� 7q����U�'�͗΅>�@��1��5na�$�֓��H���E��PB�f��F�,n;D���F��ЀyJ�$�5�Y�ͬ�iy�[b�&��yҦ���vm��J�}Bq(o�J\���Zn�Bsn�>�1免f�y
�p�M�k���0�L
�+���TU �&
%����ME:8�Y�h�bw�x8���[6����h:�_�Cw��d����ި��0k��9�:�� ��p�_(��cf�I��=e��yh��Y��m���##1Lh��&�,�h�;��_��&Л��ۈ��0�So��A?d��ON��g{M�w��f��;����z�g��^�٩�j-�Az��`jZM+��$� 
I뱺2D�����c7������M��3F�8*W��Lͧ~Y�����Y�o��$��Цt8��M��}��1�����Ƿ��o�4�xQp��5��� ��f�ؾ\|��������pІ�w۷9�A
t�m%d���N2�l�RCB�a�qD���v�/�1G�Ȍ}��Q�f��e�����K4��A��C�c1+K� ��7م>~�j����p�?���wTB~:����>h�jl=p�͵�TqrE�ɉ������~�T��I̚���	wFM�� ���	k��Z���w|2�z���QQ�/T�`����V���iu�x��->8��h2���k�����E�u�b��EC�� 6�x�RK�{$��%��A���Z�a.�V�[�S��d�`3i��^���	�&dF;���!en�.�������/�)�r#L��mh�`(�<��ŚK�sy䤦7@�ڴϵH������L2�^��n��voF�k��ĜVԒ�pi���B�2,a)	���X,یD��g'hjc�g4����w喭���j���ՖQ;��[r� p3||T_��2��:�y_|s�^`<��&vk���27��\���5�a��?�o�[���J���J�=���2�����C�嗓��#g�p�,���e�ϢN�\�]�������=�U���@!ʹ/��S��%����-�c�����#����v��nR�����w;�	��JNY?ͯ��b;[��0�-��!)��q\\���鿅j�&��h��YEwԌV�"b�b܌$1�^���bz��Y_���O�i4�o9@PT�$�y���8�k<��e"��ƕȦ��4
�`#�B��٠m[�Z�\*�UM�\�|$��I%ޚ�y��ڵ�z�L>\g:�g�0�9�����!\�u��ݛcbV���6�s�mb���|{RH��j��jڶ�ɣDuCd!ѕS?P�7��;4��6�]���ϔ*�}$Jd}�"��M���Xv��܉XR��d� �b�4H�|�c���C�wM�5��&�P9�0�.E��˃5c��X!��M�^O�Ri
�B�ӫ5)žz�*��ҍKk�4�A!�aqG
�_��!��b��r�Q���4IP�AvH�����_���"?�6��%�m,�}�R�x�D����O���%��I��j�!�}��&|��;C��Rr�o�:Q~53M�o� �D2y�8�g/}c_�����ĮmʝzN&����N��t L�<I�@��B��ϣrL{����h�\�J���49,C^����U՞�d�x����8^�љ�Ú���߉}۲�C��e���f���;�@:RhƯ���۵�$�:����=���z�2���]xnI��։�p�潗�������Q�|�9FF��t�m~������LR��p�t��U_nU��L����	S��Z<#W�����X+�/[�e���P�SGUF+P��j>cN�����L8�	�Y��=���n^�A���ì��u�a7��������~ِk�B���	ɁD�{�;_����&�]��|�Ĕ)y�����e�ʫ0��8���0a�dsMr8���iYD"4��F/p������6춢�J��?F,�P_�T�ř"z���.�� 8|�O���^![C���~e4�^�gPd:t��B��d8�(��.뿸1ς'��"xOh�N�_A�J�u	�r��*N:����g�a��S┸����q���R�R��D�@�Wl
^L�X�L�U@����Z��1X d�� ����f��c�ҷIR��Np9�?rEQ&��U�����+���X)��i�VO@a�ȷ���%�{��[�1����ԩQ��i��@�_F΄��7İ�p��'��Q����t��������Z�r�*��`��o[�hHM�+E�\��Nц<�E����Q���'�ҵ�ܻ���C/�MN��B��:C���#�2,?pv{�'Z�?E��s�ֱS��#ХHݒ�a��.o���-�D�Ɇ�(�פO)-{�;E��v��e�a��j��+��9��a)v�?�
Կ�A9Vl���$2�ON�Y��y3����ָ�2� 5��X���7O��j�Ѻ��'1�~Z&k밀�X�<��T������Z�.Ĭ,�0$�?b��?� �4�mH++.5FI@�jm$� ne�������#�ypG�#v��z ����Ř�F;���˓��{zC(csk�$?�I�8:d�JѲ&���\sSJ��ܒg�1i�X�%� ���;-����m���]M!|m@�Úƃ+��o�J-��_�?w{Fd���-#��l��2������O�{e��>�rf�f��]Ew|��:�E��E�R�0a�Oҁڽf�.M�����5J�� [��1Ɠ��r&�֕%��nI"L?�d�u��)��xLDܪ�ٺm*��#$hC6!F�/��r d�yui�XN7�bg���7��꡺M �<��l�uSyv�OW�iˤ�
��)#�j���9���ګ�ן0��Gf���8��ϴu��KwK�8N7HF�`�����U�4d"n%Ss����F��l.��CA6�BT�BJ�t�m���Ʋ�Z��N�S�K�����l@�9�ˁ��_R�����D��?˃��u���P�8w��=5߁�9��cB���}\p�e�)���x�)B6�?=��f�!�i�Z};B8w��J��;��θ�	&D���ڻ)�:��u���~/wrA ����{!�tVh����JwqAծ�|jm�# �����W�@�YW��^���P.�X�=�ue�]�l��{{���Us��9,	��W/�X�2���y h�ٓj-LD��_Q�ߴ��#ԗi���ڼ˝����FL�GD���q[��(����������v�j�o��P{�8��T�9�Т+Lkm�o�+9|������H�N]2{#a
����J6^�h��!���D��
�#<Py��u��o��D�ƞK\�R�dN��������B�8D#���e)U*�����]閧}��]���vU���y� Y�ۭ�6�g��\E�<�+48+k�z;�S��׷��%�
�x�Cw���	��j�eu�vZ�b�;J���'2�G����O��ܖlAZ�F=��+k��5�c���\���ٳ�i�|Z>�ķ�0�@x�ˆd�!,�5�b�
U�?�7��|�� 	�>|��0I2�6��۬c:%7ն������iZ�yz[�X��,2���|��J��g�%��FPm������`��C��p�:��?�c��� ������t��h\�#:}����:[|^�TRi���<�aYΜ08{ۓ��K|K�闅"��s%R�ΰ�$�ϙ�B�Z��?�������B��Vf4��5����j/�����]��e�ty��!ȭwN��л��	��/��B^�SV�~����r��C]������Wi�~4m��T��8�p_b�]�O ��s�-�����I�G��M�Fш�[���5�|ߦliW��*z�,��B��9B��H��:��Ju��	�c�#���3���䬋5�L����?��/��TTҨ�,�Ƶ�G������@���b�ci�N͍��� �ܱj����'���}D��ȋ�s�d���I����^�ԏ��ל�a-�Q��
j��_o~��G������۫�s��ҤP'�Ӂ�&���cH�?��vR���n
���7����S9���^(/���8��ڕ��Xy�~w��0���!~VN��b��2Z:|&M���G~fӱQ���nZN����:�Z|�q�*�������Gq�6uTI�^�Vܟ��Q���\<�3^-Ib'�a/dʫ���J�?pל'��!Pc�X6���يp�V��?��]IԸfd�O�L���&--��U᷎��FCi4wϼi���5m@����2�o}6�T�-'h�Y޼	�Ʒ���5z������%|��ҤLH wm?��L�~��DY �e��[��/�.�ȣ�<�! ����ӱ�HC�wVڇ��#[Jq +}���`��q��" ��s8f�ט�cMWIP�g�jk�f{��,i�P�7k�.,�T�'8�@����(��2�R�A�}����z�Ņʹe6ƒ)�3g���(A5[ޗ�B =5*YMB2�W��َ�Z���Wc3�$@�lG]�	����@Z=kU0�������Jb�\����:��eM��ZM��֛�"}.���.Rsb���0��=
}Ұ�|��.���Y�El��b�]x�~��Fp:P��<h�:cE�F�������	n��D���mhO���Q/���tb("���󥔾���O��;,�����(�<��T� *w>XW�)�"Pm�Oa}}&ǐ�Jʗ9x[?$��\�i�*X�OUA�L�D%�K��D���b�#D��бNUaN����.�
�%^Z����11l�[>�Cm~��߼�2԰���x	��/�=�|TW�|�"��"�9���0}�Q�%�7�����:!F:�]�Z��<�->��8gR��
��pF�䏻,]��-4m�	���e���y�Y��ƕ��Ʉ�"���#w�@ac�&5xiB\��*��X���WK����zz��5$��.�:����"���W��n�<���]]J�T�h֚�`�Q�J�3�7}}Q���(L�`�O$Ib�������`7E��;D��q6XL⚋QjF-�D]h�2BT��V���R�#�)>b��M4�!u)���E'�.4���xK�ӓJS�U��7��*�pK���ph ��L{�<zƭ+�E�=kC�#l'��'icDe�B��o�=3�0ؠ�X����»*�X��M@�{���Srp��[�X�1o�!G�|���(H���'k:W�]�����]�/�2`#+�˭r2�Q��ԑZ<J�,����	�\�,��wq�PDd��9dJݳ��2�N�\�M�����������z��e��dRj{sw�����Z��&�Y��"����@�ܥ"���!�/��M�W������o�{j�����rK� ?t3�Yn������,e/�fp�`o�	��[�@=�w��L.�'NwD��8-ԁ�����(�"n��Ǝ�}��(bh���� �_#�W��]"���b�����>�ט*�3;
e�6�3�����Ґ�c���G�J��́`~KM1��mK�Iya+ÊT��b����gË�ϗl�Л�7�ދ`;���C�xSqBh�������x�a,`�����@�����kcrf��%�H_�[+��Cu���Ϳ��Z������h]�Z�'���]�6�E[��@P���Bt9�hUI? �&dO����Dv����*�a�D�Xb~�b�;]*�qr�f=�M�ԪfI'��} 4���G��r�7H5e&`��qoF�Fp�>e@�Q��.vs��i5W�=�&�eW|k�n�:��מ�/*��mC�bM�T�3���&�1�1�;C[�@,�����+L! �7�S�H�0�4d6?���jR͚y�R�*�Um'zI�x�z�*�j�M"锧��S���H�d-w#�3�$o��o�bPDT'�{�$u�&�7���a��O�;T����U�].��ň!���E]��Ԫ��E��Ō܈1����D34�42.���N
R=���r�D��YO�1C�z�2�W�hs�Z�!��KD�z0�7�2����J]�3�2��0i4�W>Pa�Z�R��Qh�T�dƑ��1���Kz��H�0�A���Q�]y��=e�lb0�!\����ҽ���������M��X�Lcu2�>9W��%m�k�zd����1���Ҍ?G�y9&�!��/^�z;���/�GҴǗz��n�u�^D���yr}�q�� ��%�l��d�$K���p�����Ϊ��c�{.H�-	C��M�I�{Q�` *�8˚�����N�P߅��X��$��]9Z���-�6F͏�������z=*bF�M�3W�p���
S�������/P#�#0�&+� ��2�ɤ,3P�_�.!JY1�)^g��Mkl�C 9����Iq��(Dt��p�'DG�"�}k(�hE�D��")j��~9���-D���t报��%�:�]zՌur����5�C9��ѯ\��U�e�G5�= �}��W��)ÔSkl�-춎���h4*KH���]rI��s8�8]RN`W����A׫S��wT���/��
�����K��jDk�����%�>�)������?�LZ��{H��D�u"zE,��2�I��w���Y��V�j&��!2�C�>Fϖ����LqV9)��!{����`�*�R²��&�{�S�Q~��L���P*4�U�������^Mx��j��r���ɸ��~&�c���A9�f�pB�}]�b�O�g%1݃wzЩPɅV�I��4'�ە��`��Ǭz��X�4��~*�J���Ɔ0�]���c6H�6\UV�������k�l�A��=� ���*�{e9U3Îe2<�����rbj0�X���E(J�a<���ٰ�]�Wܙ��;�W}��|�T���Q��g���� �jpO��5T$�>𤺌v��z*v�!1D��}uS����q�9� y�|�p|14d�"��]3��
>8��b��v@���ꚲ$��}'ȭ~3kÕs�X�Fg�.��9j'�E#��D��x�Uޝ���f�(�}��I�	���8����n�4#�V�SbO�����h
���{-8����T��AV���6�{�t���#O*M�2�,h�����t����q/�n��z}:�kp�g�W�B�m*������s}5�Y-D�A���(-9�\]��+xyx���Lq��f#ޓ̓{�q�XA������+��}���]B@]�W�7B���5�	%풑��@uHӡ��F�L���n�֖�o�2�@?��%��g�<�71Q��"�b�O*���d���Y�qy�(�
|h������P��֚.X턘��ťu�5�$-�m������X�z5���0J>I �|��N��0�����C���Sȳ��ў¼���ې����d�r)�6�M��.h" _32�/�ƶ��3�h	����9�R֡��$�u����Gz�}~K��?��G��x�"��7���i���׃���*�6��ݚ�F�TV����Z�c��O��f$9�2�Dh��氢�w�^P�_P�ҿ�{PE2�����- �a���<�/���{w��G�[P��,'��g��a��h�F.��%P^��d�wb2\��E�O["�^�A}�R=����I��{i�o�T��Y�a��'�p��4�|`�y�@�څ~�l��q�k�2��|g���讕�
��=cX7��*�C8t�9W˲&�p�.*��7�9@�t��������������UV/��W�A9�t;�X�֮�.�i�Y�z�xtW�?��q1�R�U������������J���VԾWK���M���$���{��5�&���	RY��䴯��"_R�`���֔����k�+�\�'~]<�Ҥ��A����{�_1��H���U�'Pe�>e$��|�p����N���W�f�@����b;ߏ��!@�,̨�c���P�ȯ�ofU2�@.fL����m��j{b;��t���/Е����g �Betn�5ߥ��4��I
�ܩ��7�'��� �� Z���SǇ���s'H�׀k�ԡ��^������U8F� V~2�T%�_t��zK����h�j �P_�/�bڽ9�����CHR�3�B�h�ģ5YH�a�g?pP��t���/({�j[�yƢ��8���c�4�~]xczB�;Zޥ :�ŵ��'����0�Z{�����f� Z�$�Ar�ux9�2����;U�-�U�ޕ4W$�6+h�(�"�֮/���?W��%���e{���9������Ç�8�-c�(�-�r�Í�3�����m�s1j��9n��]}�wb!���!~Yx�|�7�h��g����UX��]M%���xYb��a kю�&�n�]��f���W�I^�={�7�I����� m��=����W��y��g�n̉��Z�#��:
}%�i�q��<[
��D���Eד�XO�}DW�ǩ�T=�X=��?��%U�ꈊ�.Nc�w7I1� ީC�X0�ŕ�uEj>�������.mCb��^�x�߫V-8����57�Ƈ%��k^ܚyJU`�>��ڂn��C���`�x�R�����3�A�< >}[�;���E�l�5�F�<P�.�RNq�zB������=	g�K>�?�~�N5ܱ��	�0b��̛�0\VI�=RK���*�z���ۜƛ���3���}]���eM]�sN��ڸ��W�T�`�bn7��L�j�S-�'�t�J�/.��Y�ID�ͤw�T�q�pns����7 �{w�vf��'�MT0:�gSB'������MC���
��{�ߣ��=Ņ���b%�	eŇPҮ�"�DV����L5��Q ���y�I�]#f40�t�7�Ψ�ӅG�骰D�١|Jՙg�gҽ'ۮ�*5S�f��W$k�g��� $+ܘ�:�kQ)�,�K4��!���k�y�W��=�Ţ��:���	^�y�.���~�QQ��	H�f%�x�\h+�Qd÷n6W�2����u2�u��n�t�ʎп���>îG�U!��������yʺ�NŘB��������9���Y�	v���I�����0 �܎z�����n���	nIQ�5/UJ`��AF��(��}��!��T0?��%P���$�IE�$Q�������w�f�*pP�Z����U���S��/��U��5Y�-](�;0#���$yu;C��:Od�m�;۷��T[h1?�`��6�-:�ms3|~Ʃo3��������ǽ�����fk溽� �׬[��.��ϫ�O�Y���](_�E�?�B��3��YVj$�r��^�kY�Y6<���]4�! �-w�i�i�s���)Pf�k1}P�"��U%��N�����ķGw]�o.sh�h/�,���<:r=ʏ�f���m�D���,�ce·���v4"WD��6TU�4�Ml9���N���~���(�My=CM@��Њ�Z�K��+S4�R�EF#/�U\j'�;��4M�"����O.��\����kRc��Ap�u�����E�� 2*�F��.}�J�@���:� -�˭�t�	aD;K���	 ޥᑰrM$�'ӸQ���֞��L~�������D�<���A ��r'���`Ӵ�����%v�G����@%Z�7�F�uU.O]v?X�a�Ob2Y�&(J���	���3��m$y�-]�X2MԆ�'|���X�DqŘ��ԈA��]�(V��^��=�K\R�����ݝb5�򼻃���v'�g+s��������l��Y"߮7����dKVڇW�%t����k�H����Q��f\��V�;�������L���P���k?�J�j��h�,�%<��%�����s^���彗��Y�w���N�}˿��U(�R�pQ�O-�x��񸝰]P�������1�N�ùD��+��!$�5b�K#I�:@Zxb�G�郱u��������nL��sN���������H{\�����)��+\�3��u tPz/���� �xl�H�3a�UQ��5Ɩ��y�ۿ�����"�!���,kb�jX� a:+6�5�;ݭ�)�:C�"��P<�;K1/ᰃ<���zUЫ ]��g��j�ä~�3OP<Mk��J��Pn�*�zh	�m/�X�t-:]Grh�f(�T���K̡Ӫ��k
��s�d��� <P�m�@��e�L�$��y��s����y=�F�#�́�H� D�J��~}p�M ���zXI�ki)�J�|����K��SN'�T�j��}KH�%)knK�J�a�o��%������ٵ �WEl�PUU��
�L[~c����w�,/R�.�Y�������Pl���"���4+�jz�_���3/���B�YٖBc��W��(�(<�A��:�%�bm���L�-�`�*t�;G�[������-�r?%�{Ռ�������n���[ۯ�9Ja\>�[��y��1X0�)iG����q�P�L��N��@�i�QGpN�}���Mi)����uC��v��SD<�le�
�3�諒�Ւȁ��s�+]�>[E�M��*߬�he����JYao��\�@6��C���w�\�Df� �b����z%�Z��&E����Cٌʶ,�f�&����	暲���jvW�Ҩ��4l,L|] �VY�#5�lϐ�3Qnܾڪ�%�tDOd�m�˵̠���)
/ܽ��~�Ϙ����m1B<#�]C��֖�w)a)��!��d`f�Z_I2����/�Ho ��k�|������W������O� ����~�3�	c�p�6��}��A|�'~��$ �g���:X�Q%��fiw�P��L�!�G�b\5�Lr��HcQ�T]�k�6Y:����q�P+���S�%ۨ&Oo��r�)�d�ݨif��M��y��k6���6PO����)`�Q�)*ߐt�>��XR���s��M��q~-���/Pl
�@{fc��./���6�&�p\���P�"�d���:���j�WX$U�!��~�ϪRu���Zѳ��<���dbP�'��7��~&���`�%T#��_��0����M`1�OXIi��Υy��w�܌�w31�ۉvQ��6�.9ߎ��^�͗����3G��/#Ew�3*�>-Y����(���1|;�%; �[p��d�.uN3�/���Ǉ�����N�#��_�x����.*�&q
&�����Qi-	Ӑ��PX@C�!43�qg���_X%��T>ȫ��h�_*z�/fW�pK��6������5�HC�͢�Û�>z���(���_���6:*�X��nj:yu>����<Q%pky�f���O���E{>�������q���aYs����޼�ocr�>��A�Q�Y\�Fk�8I�|�:�x-���g'ߣ���v!(����'���W��+̧R�K{�bE��OsÛFj8�6���6�}%},�%#��-؇�,1�H��^�*#)g�R�M�M`����P-�51n��o=ݧ!%K {��_�Q-�>A�6s�b6L,�^W���K�)}���!�2ab.4yWN��H���ժsZe��q��p#8�|�[Lkoⷓ�e�)�W�����/��mBg�ўd�����۟E'�uc�aX��5��4�g=Z r�y�_m���lv��$�OC�åbS�p`��q��:J�;%;Z�vb$]c��,�_�j��<�kvL�_�E%��� �]~�`D-GEC�����k|��{���x^d�"Ei+�`4��9QDl}�$����0�����'i�}��Tw��[ͫ�[!>{���#R�k�	giR���ǌtS����`ʇ`��* V�aj�v:�6��M��-��i�; IO��gce'n)G��-�>;�	�EP�;��5S��q�tN��Ӗə���W��θ�\WI�}���;�t�̧�r>�X�����4o��8/2�b��H�U��q�)0t=h��� .� |f[3�Z���AMں�����I_��^&ݻס~�F�.E��׮�B�)�JS�ߥ,�-Hݔ������#�p�j��%M���g�\��/�I�q|w�h��ȁ�*�C���2
#�!ķ
�"���d?��Y�W�h:|��
֒�MzIl~�����\�����S�����4f0UY���˾OB(�b��c�2?�#X��"`}-��w-���SX�'�V(ؒX�ind,;?�;7��^K���i���fl ?�	'?�ɲ�X-E�wx�˂����X���
P�\V98��r�>Ч�8�����T=��������8?���&Vk�%�v��'��i���k�Z�4�"��.��O�?��bs�M���Q+��G�3�;rhiy���Ԟ�~����[13R���z=みDl��b�d�C��W�O:�o���Pt�$��kF�p��D���/۳��ƵԽj�lD�	�_z���xi���y��F8��."IfĶJ����?ۗ��N�)�/ˋ�5�U�L#���:1��wu/J/.�z����A/���Eѥ��S�!�l]�aX��d��l5��w��G�\���l!��N���<f��S0w������M���y+�5����A�ߞ����b�����n�s�2%����T���se��7���5¼�SԞ��]�� *A�PF'�N�Q��JG�)���~��Y�b������΀W)r��a
6������9
���D�Ĳߖz���L�Bd�7s�F�4�O��@I�8�����c�D���Ӣ@:t�c�[��p웜�a\�}C	u�����>�'��͍�چ���bt�Y���6����/��0~`K�1ᐙB�9Q��9���e�|��D�ߴ���&z;x�� ⁰r�.g�|�T�k��	˯
�[>�꤅�}�s�e�3w��G�fc�4az��\�/���|�Ɓ���j43�����Ux���#�A�X�� Ϣ��4���
�$�}�ıw�a�0:oP<3��u����x��X����$��q)ʫ����S�wVăs���z����cl "���;܏�V��%f���v�b�Vp����D��K����)n.T���։a���@�z�4�|��3��Lnj����E	��l�C�z�P���1�f�^v.�y4¶�J�Ks��dx5���BH�%f�/���RXru8N2�I�Ƌ�p�|��W�\n�Tb�)�Q���q���k��Z��z~�|�!�Z���*`\���["�N���o��Na7�������	2Q���ެ̘��zŋ��-��G��z����?&�Ԋ���y�M����kdNQ�����F5u���H�Rѹ&5f�1��@bxk��Ȏ��%~)S�%����ac��2��(_�*ŀ2����r�^'����f:s����i��)��yr�����X]�9G˙�!;�Hi�ٝ2�'<mc{6q1p>�����O�\�\f?H�����`��"��׷k�tٚ�KN����wp�����/ �cDh�el�;�ٝj��0�tZ?z�Wr{,�/g�ue?}5��&)ъ�Dm�wV�ڪ��%ӄ�=�W[��Y�UTĞ����u@��z�}:$��������K�)`�������9�c�]�w}"N%�?3�K���|��1�"�S����m.����ui��m5�3/�}lB#h9v��M�0K�ܬr����Z�>����K����tC%3�9F�/��S��
���c-�t���kR?Z�=o�b�R���q*���{�p����+*���x(0�l�G	/�'��Kq�n�隷8;1�-�ܘ�{�]��
�� d��ÊVKL����áy.�8�S�
��"	M�+֥�E�T5��C�Y��ȖA��@G/n�fK�%i]�񇬌�O�7��C����T��zׯ8_�3ր�OtйѶS7�	��,+��h�x�
�|o�gŞ?|�X�.i��2�w�{qK	:�:�v�mV{�v���|�h�Cwya�TGF�%��m�?�E����au�~����o�@/�n��WM�]Ř����q�=����s�Gl\5�M5��*��F��)h~����<k�}�)�\r��2�w��q�X�V�f���t��-�� �;L��y�x녆�A�t-�ß������>9/��K]�	t���E ��w�d���2KK}��&���dv	5%�sA!Cr'dp5�d3� ǽ��dq�T��]Y1��iy����#�pp�|���0a�[>T��O�p�N�;� �2d8~,�f�t����2;6�'1k�50Lr�'E��.l؋�/���et��D
�0d�����o>l_.��&hnw�﨓��1��y�i_���`��n��Ө��Ma�!��pTy�c�82��]@���Q�DW���C&6�];ԑ�[_ǳ.h����W�|�o�vx*}�*N[ /��@y����(@yZiѳ��et�qn�5n��ZV�г�)�N�kO[S�m��}�\r�M��K��o�ߕ�;8Sh�8������hЛ)ޢ)�$f�U�NF���ihV_?ux1���vZ&5���t1:���������86i߶O]���ɠ�����E!@j[[��3����^0�&���
�_ 8l���"
��+�S�~J;��QG�2|�s�0��
O����mo�v���@w`�Q��5���)�!|�)P݌���8զ*�r�=WlxҭT����.�LK!�a�p�������v�s�M�Cy�~�&1A����n��k�4�j�
��)EzDi����D'ę�`�2M"	��o $a�˭"bx�NӲy�9�¿�����\8;���$���:�Q��	�^�|���ya�@%�ʹ'B����_7;�/��_D&i=D�#��˟��8��iUѶq-�e_iB��=@[���g�N�S;�o  �ۼ��H���-�	�>K�7Ƿ�-�v�Nz6^��Ɍ�����{�KÊ�E���i���k�	\�b9��W��,���>f4�ۮ��+�3�m\B�@:]����T��Wkr�T�4�N��A�‾uJ�;�O�;A�@�Z١�T�����+]�u�����������u�|��j��^s\��n{���eS5(�� J&ڌ�"��̥�@��sj�����K��,ߨ��H^� S! �3����97a�֍��W�D?{��se|6��:6QZ�#������Z{�vr���ks��`D��Y;�]�>�+V�� �X���k��T��]W�F�O�^�
y�^��БS]J��x6%m4�iEA��Bb	�U;�a�^cM�#�щz�����{�F@��l����h�]���x�՜���M#�[��0�,�H�jjf3+X��Ϡ�Ht�����V�zь��'���;sNx8>{�G�֐'�ʅG?�2q㥈��<�Ƈ,#b��4���6��	qJ��T�c��Ґ9�P�X�7�9+���a�����#�R���YtZ3&����U8�b7I�1<V��̹�Jy`����PG>��m��c��tuJL�֍�ٯ�%N��Ve��	\bH2����E�_�B7��Ԡ���glt�e.O��(DK�ϒ�G�����AR3-�`*��;����T��m/��/��)%6҂Ȕ���_�Q��3ӐI����r���G��d��Fݙ2E���\�-�_;��<�j�\E߅�>�n.�V���Qgc!?{C���}qy�L�N~o��.
>^���e�ؒW^�C��8��*��͈��b����K�D�����t��C4oCi��׳�-	����z�r���mo�Hb��9�:�����͹J��EFЂ�$}�m�1��N�Swbp�0��2nJUǿEv�
�[^���� V��ӑ��ooS���pL���4&I�z�|t��b$%�^�&���4��֜x���B�]�65��~�N$.��e]��ިv�r����_I#`�ۼ*R��0s�����K�:��*J,����$�G��_���E]�.�+5�`�j����p�+���"C�*���O��n������ Ky��<w�;�ނᒕ���z����kV\�a��Zy��o�	��jf��0ό��v���'��a�:���'�q���*���x7:n N{�l&��s��&~�^bt�L>�ڲ��������ZI��>7o���h��Zio��[��gR:�-��=f5%�����������R?�KvI�B�;�	L�2�<�����ԡ�9�EwP)
�<.�뙹p�]Lq%���|�yU(d���������cR_�ª�d	��"-0��+z	2fN��ᩬ��21�&�ى+@>���yn�Uq!�!�@�~�#m�٭�G�Y�S���?��\�t����Oo�~�@��x�� ���o�{�\�*xg%%�DQI%K)�P�2G�A��Q��xA+Ǵ�(����1�u���U�?�r���Wo�9mѧ�V�z H�߳/&mr/����V"�Kv�0�?��_Θ�>p�-� ����f�?o�%��ۆhM���/ld ��Z�C��6�)v����K2��T��&Ym'i�@�o��&�����|u|8Z\�\c�k�7Uɲ����^�Γ, ����1���/^�PӢi6:�
��$@�$��W\1�
�^f��������f���Pr��h�Ln��W�z҉��qs��իǛ7J�Yϻ�շ"i�m��-b����?�'��TM���S�;O��?̀�ڀ4�Os�6��+d�s�n����Q�D"/p��L�x�x�,�ȱ"����C�|����Nq#Vk��B
����&�g�zPS��F�ӽ�$�|��?��.#t�׻u��Wȷ�Qgo�/۞�U�+�����UA�?Q�(ĴK�/zI7��D��>�F
?���9C�Lpm�[��î��]ec��9�Hr�'�,�l�_A�l��^�x�yp�>9 	K1)���jن_N*���R����Elm3��9��%��\A�瘙�J��`&�ʿ�ȿu
�غ�P�#M��U��_UI%��:��z���O����s57�}�X���=M�|�؝�CI���WE�^F�9B_<�ߣ�R?K7�pyY�?ȠG�@pD���sX��N��]�(]�Q�̎;~^��1�>�m�m�p�dU�>�z<�9���S~g�/?������:
����p�eJ��Y�,1M&�mt���$�M��D�)���F�E.A��n�Dxo��!~�L��9�x��&W�&�[tw&��Ma����;c������	=���/!��z$z'�Z���Ѧ��+%�ϰG&&�7ۑ|0
K�`���L[)IZAg��ټ�
 �r�����?�����f��U�YW�����������vX44�BU9��9�~�n�07 {y(���p,jA�/J��ʋ^mʛ���Jl��ـ�r�u�=�U9��`�@l��Ql)�����U��m��Wt�5��Ꮠ�F)�vLݟd���u"���N��ğ50,I".P�8=�56�YZH�	���ޔ�XZѫ&����d.�t��x�$5�n���H31�ǏZ�e$������G_�"U�<����s&�zb}�c�97�1Nߞ�
X��i  S/^6w�a�"~�5z!����>�W�!���/��}d��M�R��>�����M��X�RAD!�ZO 8#��
]<z�UdOO�/#�&x���N���x3K��&.��9˥��5qH����v8[�+%{���ߔ�A��?�
YS�u�Ȑ�v%Ǉ6�u�EB�_�u��;���g����E�{�}�%ҝmՈ� �71N�n�"�!<�
ȷ�F^�Ҹ�^ï��Dz�:g�K�J�p�ŉ�/ܕ�N��u,"��8= ��}I�[�3��ˊ���f��K1��c?fĖ߈7;`?ə��tp��١i`Ga�|y�H���y��϶ݷ	jP��Jq���Z��������]
P>��:߇�=���}��-������6<��d�j2!�����I�;x���dt�OH�����H��Sů��k�T�g�W���y4ZG[ܺrEQV"]����%�,��{l5I��p�`H��ցF����#;%3�!"�%dn�R�@$�+�Vb 0Z0J�=���4�-M�*���|�URf�%��a�#�ҏ���=A�
���^K^�q�љ� �\ &����7�"5pm�xB��ќ5�����G�'�b���@��\J��H��g����M���X�i��@>Ϊ��C����]E�\��^�IY��)	�z7�8-أ驾C(N^E\�J!���5���b��<��o�dn�T��� ��Ο�j`݀�X���3�؟��i�j<̦��\n�ޒ�@l�5Z��Mp�A
\�fP�)0�}/�(:�E}�˼�f�k�y	�$o��	ê�����H��e	��7y��7�7K!�1*n�|�FuV�3��kR�/l���xU����sϰ4��ʒ�7��	T�5��j���o�LR]B_�q�A֏r�鼻	�P=r뚱�V2A��Ȇ��QA.�z�]�$tJ����gh�d~:b ���4t�I�ݳx��<�U7o>����I��%Pb>�"hH���BD{Sꕕ�D����Y~��̔�:*��8�Q�L�@�G�4�SB�V���wV�ֱ-��l��5U9r�d('�@���8�f'7����MF#t^�UN�uLfĈ#>�쐃�jK2cIS��u�0�z�����L�s�X����{�XSlFrȲ� ���	��rيH��*{y�88�$Q�Y�	�t�T-l,��<0��\	!�o�/�;��Y���IA*cN!U��x�ֆ�vZY�M�Ǒ�-=}@NY����hlV=������,+����fDa������[�݅��`�w���ꟷ�E�� GL��/0��<��#���b9�'�{��D��ᯭ���M;�u��n��Ƞ=��䕌\> ��!��.��x��|0m ��=z�o:�xEE�. GUzf�����0y<0�g�5:	+f���k)JJm�]���~�J�P2ַ�w%��#O
 mFm�'ҠP�2��3�9���֝Hzpm��iJ��~�t�J�h�&�d�+���p��ۇ�0�lc���+��|����U����ϲ��wY�ǎ|}�ljg�~�+�XdZ���C-�n��gĶMc�`�U7��-zO��ڋ���&��mK9�����='q��-��x���i#*5��[����$�J�۴�4F�}��!�gkbVr��o<J��3�65X��z�Vg��bΨ۫_��9W�!o+� UX	��/;���y�w�Ep�%�oVz�1�o�)�=IA��MB	��&�X��4P�SKd�����?(g US1��#��p��wne|P���lx��'�h7u�s'�R�4"�z�OH�u��{�X2���V���UPC0dy����-�.#�ԟ	�6�x��K�����I��9ީd@�5�6?���d�Q��8v.xiuF.��5��tN("�S`�N��/��m0��v��*O��DB@���ޒ6v�N@�m�q��~f���(�����dp����~������0j��X���2�"F���͏�)nD�͂�_���E 7E� ��%\xO��6t��IdS�=/ o�,�$4�Y�E�(�C���#��QB�&��z�#dRb�43��h	ۂ�����\�e��s #x5c��X�&�����\�"-Cn񘉚��s�
/��~e�G5�B���Y3n�2����mMR�T^�U�]�����l�^�툂��oeS�Jg8!���$� Ol�e��Qmge���G"Cp2k�6W�����v��q4�4���������UI���"�F��M5��Q��~�I�Јo>xm��S��gp<���!I��ז#�,�2��S<![��U+%i�fA���;ۺ��&>��c@<G�Bs�D�@U�ɝhk[R�!�.4�!��9����P�1��gH︿���w]�C������;6���8MA:?���;)�Kz}A���Np���E7a��ﾤ����ˍ�+��s��{�5:濒�<�ܨ4,!���B�(��������j-�\�Z2�?�=�F��Kz_� f��� :*1��3�;�W�)`�\_�n�S7�X�5�+r�9�Mц0��z�N��U������ƥ�XM�EbJn�\�'�1�T���ƭ@`�)��!��~h��'S��W0&�tNf
˹�ZV<D��whF;�Gb^;�׍���JyAbO�o�ch
2�:".��.��U�V�6NVj�%�j��!WN�4��UR��g%��ƩA�J��]>a<tY^3���Y���q�'����`_e����VFA+uA��y�h�k��P=R��2��2�KADE�#&�|1p��Z��I�\������$#�W��;�aw*��(R
����p���0y�AG]�Qm�8�.5L�RKw����U��6l��Qv���M��*��Z�m���|n�����L��;s��<̉�@>��T��]��mQ*���8CJm'���?���.ǵ�Ւi�Tp"_��C�Z4�曧��%����n��@*�8�5Ć����9'��eo��\2�O�r��CH�E�6�kF\bMUۡ���sww�����X�7	�{&�_ԯx�O<�/��Ȕ�H��3ǷI�`���(#�[�e��b$�_�Rï����Ow��:��!���~�{��]��=�ƿ1KQ���v(V'C�(�O@իr��={XnR�^T��!�E�:��^��q�"sH�@��)>�h�;�W��}D�a�#*4#?�"zok����ëC�I�GE���F�V�3Jb?&0*�=r�|�>b�I5��v3�V��7��x�i����A���3�y^��k��.�Kr�����l�@�� un�t�"���ȖU
�a\���Z����F'QG}Pb���������It@i�H�<^=�W[]1��#;�&��A����Ps	J#{&`��B8�q��<:j��[�Z��_��1�&\GS�v�V�_bY4� W�K0��N�	�z�{M{�scYn>	_untD]Qږ`����.��%
����{Y�����@�,$>5)�e3�ڲ�%�m�7�d�DPW><���i��f���Ι�oh=%���{��2RO�=ݖ�o��i��6zKg�M�X���� �eω����Ֆ������C�a#
*�q��;/e��jZ�2Y`t6J�-�y`�󶃊~qv+���mH/�!�;ԇ�g�_�����2�S����G�T"G;��G4O�13@1��v��V�2(�x��10�yG�l:0y��,�J�>L��n����WW li"I��L����SȆߤ�=��W�wE�\�����çHg!K�#k虰��^���n�t�;2�p:A6BljM�YZb�|�twr%=8�_���i !�v����0��S��T`���J��ޯ�Cb�����Oĝ�E�0Hz�Miˍw�$�D�C�e?��{]�#Xc�|��%�P&�2�赜G����*�nn5ȇ�"0!�у|$r@EZ��۸@���}���l�Q'�T��Q!�н�P0\�[DXl7�YͿ�ùc�����8�H�/�XRr��V��x*���.1�v�FF&�a���]�cHլ�z�Z�	���A9�X�^@VӴ�90���.0�<-:�1�ˑ���%!�9�vH�~�q��'_#�VEAb����.�i��u����.h��Ę�}�q�b_�(N���6k=��Q��kB�qX�
E�9!����v�Ux\>���YQ��6�R%S]yV�sT�Y� ��S���Ԑ�]������K�*#R�|+b؛*��+Gg?�1��epW���rʹ�M3J�y\�pѠ��!klT6���8����-Gw����o"S�\��:r���}�U�c��p�C��)����Q��d�ƌumw������4o�� �ۻB\/�yL�d�ժ���ֱ���:> ˈ�6{f�X��� `v@f���d�5[��o�<�a��_��"�u,e�i�N47��L�� �/�m��L������ƪ��H��1�Qt���9k���m�����bQV�$y�@DW���٨�+��N����&�i-ۧ��H{���m�ǮyÏp����!��K�~a��^���n��nV^o�M:Z �P<p�p��ÇP̂ކ�[?�n>u��#N������܀�6���b����螺aa;)u�W5���&8�������(L���(S�8�d�7%���d�>ԅ訒B�:{��et�@�����.;�?q�a��<z��#`��W)�N����n���#��>p9=�Uk�- h������2�(���@��/	!��gЈY9�ӻ���!MO���B(�^�2����͙͞7�B�%�}Q.+��y����I�(�C�\Xk ��+*7B%������by�S����x�6l�g�� ��>��]�ӑbj��^@�����"pma�w!u0W�\,C���?�)��?�5l�M����\r �7"8��D�l���롊��6z��!�l9{�"H�QL�\��>�Cxu��yK��+��e��T�#�_�����B+��c;�@/�`r��
��`�g���2k�%\|y���2� ��dœ���F�$$,�^-����6��M9M�e!k#�P�k��O�{��� �I��&4�mQ�f=I o]�1&�l���j������Ą�@��	6�#��gx%s��{^����`�:�r1*F{�Q����M�b��}ؗIM>�]4�>e~�(��g�W���Gkرi���A_:���f�f��@��3��Om�7T��~a�PөZK=>lw4��#0L���܎�%@����6"���bN�py�B�b�'����>�j�P�y�쇟{(Z���ю=�����Ȍ�J�5��1u�c�/��$����➫`�h��p�G����o�9�Z�&H~K�j�[e%�� W�J�CW)��4�MK,�Ԡq�xuA�6)�ބ+��Ϸ�va$S��p�ǤF,B?SY���C��%)2B�%�E�V8��K�ﰗi=��~!L�+I����y���F1;.n�_q`Mmy��(ĕ�o�]��Q}^��L��9��c{��I3�{&4�����aDCR�nUW�:Dt��3��N�Y��jyJ3�.g8�a!��;��f�on�����hJ.�Z32��Gjt:��ݝ�qI�	��46��U���s�g��WfZ����Ҽ���	��I���9<y��>�ܦ�<��&��1�%����8l���d��C�O�ԺD�`�!8s��mB�����y�����7����*?B'��GP;�5�<T��>��8���mV���ȃ���e��W�c�7(�:+��]f�̠��(��L'��P;@
<��|��ϧ9ҳ<`x9���:�tj��&P���_�\L c�dH��N��'�;�p��14�K`'�APg�6�l%oc�g8�(��J���u�������̻���y�V+�+Z���|��H[-�3��m��ݺ�� �A��rxכ�h��Lc�R��n����|�:�Ipm�G�U�K����i,��K�3i�y�=/;��gC,��sC�2j[�� �&/���)�=�(r����\�*V�c[ü���0�$G��}��ɗ�~{�}]�:�-I(^�ک
[�]�ԡ�M�˫a��h�9fW����!�x���Bt��k�è�Ņ�`b(s��rjQ��b��US���BڰUg&{d����;{��88�>���wF��Ƥ���S���b�ussRȌk4�WΕ���ܱ.��N#Gu'��ݣ�Ӫ���F55#Gڧ���QA�U%�A����%�����,P�J
O���0s����Q���~B�D�p��~r]���+���F� RJhU��N�];�h1��u������]�����}.>3���3Syo���4y���7f�	�?}��t�Rlw�g^�$2�-�@��V��������'��J��B<�]`bT���^���
��d�@ӌX�YP&�ZS�y�ܺ�N�8)'vu�...��PsYa��q���+�/��/�R�A_�0#_oI���m=iݳt �
gTX�>+��AvS����K?����U*f.�U��0E�r�<H�wan^�3���Z~������ G0�Y�����F���N_b�����C��c�ϱ�L�Iࣿv�Ϋ$������y���,TD!j+W7mg��v�X�ڏ^�����%�$��"^���P]gɁ>u��=�jt��*��4(:�CL������ _XY7�Xu���]�Pά�x\��g�=���>v��m�/Cx5�G��P8���3���>nƠ{?!׿�k���e�-VfOlzֻ��6HI\�!���N�(H���Wu�����*H<~a?ۘ35Ј�Q�������t�[ú-��]6_3��.�K{z���;����k��Z@�l�1.
~F B���)�fr;`��������2��#*�Mo`�β���u2H^v6�3���?��*|A�F�%ZF���+t30�;�V7mi�;�Nf�����nˋ��ڲ���1i�;�N��ze��.�D/"�9���^[S��'zz��V�<����b']U!А$̎sz�,��7�H)I�������a��WL�-��y���f}(���QP�\�)"�t���!��2��C(9l'��O��+�2"⿹'�^�Ah��A5(��Z��!&����6�L���� I��z����r��}Y�#������į�'������{���' �3����I�Q���e<~[���qD�����roz���=��-Z}��������4߹'��j�.G���x�ƿ�#ܻ��C��po�*���+�oO�Kt�!=�����m��t2w*�=��=��v����п���C= ��+��c�I�U~�ڧD�3DMt��H��~�Cq܃�ڲ�1M�ϐ	r�k6�K���^^I�VMO\Tg�jl�1�S��&w45"QQ�NF�1�3"�VO�,�����S�_6�tq��¨�
f�bI4a���->����[�v\�q�$��ጹ���_�.ŊN6��S3K���%I9nԞ�(ʼ��Z��s���2��wL���ƙ)������А6S���#�`U2p��A�1��c=����}&�<��<��0��1��B��dHA�ߚf�u���'�ﷺ�ݬ�\P1>���P��~!�ʏ2�s�{�p�
�C̕��n��|p�mI��~���C�M�XL�8ף�fA8/y,_D☝͠*��c<6~v���}g �?U����B�~�a0�W���`��(rb<�w�����Zϵ�J͟`�m��F��y˄�pr���es���w��`s����a�r�i�F�^��u��j�X�lV¢�tɺ�ߢ?��rk;2 �^��(�~�t�� `_u��2���&��ူQ��o
�pml���k�-�ªH� |ۿjF\A{���4$(��_�u䳊�O�	4��F�((�T���< ��ͮ�Ŕ��!8�!�Ζu�Pk*��F&�4!�u�.�y�}x{h�Wx��������ǘv�\<i���f��~�n�nM�G��Կ�h��v�z����9��=��O><�o�İ�i�N�����b��f��߱M�������e�eSY�Y��]�Ɓ�-Y�M�O���2M^Q���)!�v�n	�g̑1�춽�^3�u>�,'���"M�����}���п�N5�����Ő��X�(�Lk"��#fO�5�.��T��.�,�c���R�5�u#�(�M��Ѽ����V�:��+�n��\�.l!�����C������6y��b����$\rn&�ᶤ����ʭX�$�e���; ��q���9�zyi���ǉ��͠D���Y[d����XY��QIo�#�>P���=�4��S�<�ZdXk�0��Jgܙ���l���� ��`��l\��ER���y��/	=-�*�PTC"���Z��Bϧ,�Ġ�i/Ӷ>Dm��ING
L����|��<hu�h��}�/��_��k����`�]E޼D|P#U���|�5t�#d�Q�Q���D����_�~I$�*��Г�0�}A x(
� ��m 9��!S�4r�`�U�V	O�a��	��=���q���~��"'��u��v�(�=+Y�?Da����c8u�E]<��j�JL�J���HW���?^�w�8g�*s�&G18�*��ڎ��T�p�������˳����2
�������
SZ�j�� @D�nk�HZ�I� �0o�(�����qI�&b��h4��7�#�_sc5�#�%���Nh���l6Ov�ܠ, �!�,&��C@^���DA=e�;�}��f_��jR�!�v]Ó�&z6t�Y#Tt]kD���1���ΦW���Gj.2����NQz�P�:w�Ԯ���daZ�/-�������jl�]i6:��)L7;Faz�V/Y���X=K��yѳ3D?ۓMԲB�h�އ�ߞ{4��;��~yE/��͋�\ϐ�F�%�ˣе�è�F�c�����}9�J�| '��C��2�} B#�^%{��^��)#U�ߤ��Oo����k;	�W��3�2:(�m��[��dU�.t���	�G����Gy��^��s��ۇ\F�!۳��W�m"�~")Lp�����6������P����W�VD�.�s����Du�w:���.���i��N\\1�j�K�jBh���5j�ߥ�Ǜt+d���֐��x����(n������n���N�e",'��$���6}��?��������"�Z	��L��cBp�1�K�\
�;�)�C�L?Y��_8����8�u�A�^�N��ښ�
��x�BA�{΂�#&�@�(�N�Y�ޭ:Huޓ�A{e�-x���$g���87DOe{|M�ֶ��|/uD�xF�D��(�fA]O��/��xbQ�?�S��˸ނ*�<�[ݜ�T:5�����~�(f0J�����D��Bu�h�Kf�`��o�S�L��F������ʨ5z�8d��;a�l��y-��}l��]��&�툑�����W`�o��!Vb��t���П�Qz<2|�K^�xv1S��N�~8�m�vu{�I��T[������j��43"�T�~��#��v�˯�Ы2a(p��RIo����V!�~�p
^l!<2v�	��\��|=6����;t�IpO
�a��im-V�o�(�&���t�mI�PZ.�f�%~#�HM���C�Z��:шJ�!r��<�<������'`��]�x��+�ɼn^�LҨ��TߜѺ�#�y�=f^�Dq(h�7p	]�w^p��&�{N>���is�lt�}C�X�z�?~�1����c�?�Lk>�h��L��xFZ��d�ΩBVt-u���~<~X���0�N��'�	�~��n1�>>�ߣ	Pk�(4~ъ��B���^8G� �����횲,v]�^9�k�bֱ�9)�WJ���$]�vkH�2{4�
e�x��V������{0��]}�t,���Ȏ	�2��w���x?Ҿ�������L���4�Q��g�頖��۔d��+q��Z�Aݿ�X�%����Mo-rb4�_�݆��YLX~��0sp4S2��e�w_dD���ȓ"�����2�*�X��m?z��
N�,3���W�R�����������_��F�-E�'@�.[]��ُ+���}M2�~��#�Ԩ)��3d�9�B(��?�,S������<�=�e����+Պy�B�6��ξB{Mv:���Ȫ����pd���ղ�ާh�$Qāl�!א �'p�����t&��ּ��ֈ*i$�����$N����j�T�ۀ���!��׈{�P��}���X�|� �^�(�`sK5b�jK��܍y+��I0Ƽ|��mY �Wv�!���ub���_�� ��v�`��=���%�z��j�Ř�SV����E˯lH�sh=EJ���9���!������T���2K>�/�z;C��B�1�/ͨn�'m?����޲i�m�ol��V"�v&
�Rf�q�����ZSxB�] �
5��r�G��@�|\S(J�J���U� p�G�K(��|�Ex�&��3+�le��r.5���)s�''�o��FdV���8�^?���T�AѽڐE�T3Z��fe�
9��cղ{z,���8k���&�p�4����l4U����g��`	�����wH�֨�^�T�
>�V`��R&��B2ݚy��z�
�-gR���`N�+���5R�'��^�vmJM�5���_��Q^(Y�H��#���" D�T[dЦF9PlP�Q�秽S	�U���`��~�p*w.��yn�$B���b;.'��>����wR�%��eD��s�,�_wz0��)\B�D����4��U�8@T�~�춄�Ę�͠ݩ�:Pr3Y�Y��/Ԩ�g�I3QA�5��/$bݕ���K��O��!�,���7��!��:��(!п��e�'G��88��Ĩ��zY��`(�n=)s�H�摔�?FP���p
�r����JGA���ў/�"7��x܈b�P7ݹEh	��<������7��ھ��U����l(���\;�ʚb��������~��*���(cs(��h���&`<�h�1a�s����i+��/�wT�����y����wr<28!>G��܏���Bw�������:Y	�?�rE��&cJ&gfc���2�@�#���MlpT�!Kl��aGXc��u�L��ii����h��8�rqK��f���>�ܩ����(!5����r�vs�͡^h�B�P.��d��CL�T�.Z� ʍ�3y�.���2y"Z��vU�Y	�]ë�]؆ӱ��G�6���LߊI���j�t� d�
;�J�;�z�Pu�����("U�kLqm���7B�\��ijA�1�M�Yc�� �n�"L�`T�L5*x<���"y�|���8 ���,i�9t��$A���A���o��j��%��c�,q ��9��F����sH�@��e�L�F�5�N��vp�U5��af;���%��Z��5��|-�t�R�q�7���Y~*RE�=�p�^R;��Q�*���:��X>�CD#�F�FxV�*I\�i�]��U��<�#�oG�՟a��5�>QŞw���y�z���D-��\��\������r¦V�~��4 �� ����7������|*�2�%��Bi���nbm8�Z�,�	Sq{XJ�P�O{��f#D�8���A���O�&�XJ�����b�B��҅�n�Bc�x����N�����`amKV���(Nqr� �g�3�ŞP�قJ�M�����I���sk}��{�q��J�I�#�z~�D��/���?�����Mo�g_KQ��(�h�qlx�������Tdt�#�����71>F���&�;���߹k�Rۇ���8�ǫUx��M�v�m���O������`���3 �ČJ�SR2DlUSz>���N6�[�"aY�|���Ҡ|Ao����W��\l����)͌�6lw䬒`�W��Ι4C��G/��D};OxȊ���7�?�y�Ɂ�P���E�q�����hG�W��J�����G<��a���xC����2�`_����ɹ��4t�f��Ͷ���:�s�0��%�ߦ1��-}��������*�8!�e^X�6tn j�om�24(�m���G&'��)9r�d�gC��G���T:c��8Ր��)�^�T��=�s�\���Gt�6n���nIDE��3�B�}�,�L�	~���B�>�� T��������X��u2Ɉ.o�]{�����zٻ|��Zo`E�=����	�I��r?�-:�A3y�C8g�@Q��!X-D\J�C�X�чm�z�t�X��
g2wJ��������U]S �gBti�'���Q}���%{Ih������jr��5B�G�7٦�1`�@�a�B@��G5���82���ɼ���c��C9	@A%)pH�z9��߈ϕpRq�����i���`?E4Fd�0!���={0��@��(�>�S�$���VΝ��:�iC�B��������=�	����Q1�0}|��'�aS��\0x��,C��F��4,^~����L�W���<+��Ʌ�%�	�>�E��s��5����y�z�*}�1�*�e��*�B>�0� |}L����XM�0���zo��ӸX�ٝ��3�DяXdᬤ"e�ܞ?I�V�O%�$(��߈����ޓ��/f1/�.���/e�/ϫIb�p	�ťF�}��A>盝� 7<�!�L�?	�����  �9��zX!il�A ����9��B�-)�cBB�2��d����
-˴����m�"�T7�;����)u�b��o>NL,/�h��g�ԴD�b��nv���j�}mrF��їz�LI|�ߥ9T[��K����F

g�>Y!@B��{GW�|* ��'�s8d�y�U���A��}6,��[h�A�(��i�W�M0���F���QM/6L���v��bՌ	�W��)u� ��Uk '�4���C6����,�Z"��\���A�Ʈ��P�L�s��fU�x�L�<[=�ȐX�p ��.I�N��W��1*��?�-B��2u���ӑ�����P��D[p����[��Nk�?����7�@��}cBн�y�C�AB���c<����ߞ��/L��G��%������{7�Og�A� ��R)Q���aqJ�W���ӷF.�F�%w�����q�H���m-�m�/��Z�K��🇎8����@#����C�
�
⛂�V�$>�o\tX�M�$T�ZGs�G-���E:X�l;�x���\gE��
�g�oȹ�j����s��4'SU�$C<��VG�;M�z�jw��
W���4CM[? �ٞ�&JϪ�k�������&L,�0��&�Y�y�X_%�殝�)��8�����>����5#y��aM����|>&�˦U�Њ��KNI:;�k�f�g�φ�:�NJ�]N�NV��-Ľj����ԋ�}Q�=�( o�H�#�eP��A�P�GԦTa�BhC��u�9���r�p�[ͷ�H�c%����b��m�K�)�	�Ș��@C��	RS1+������WG�m4�-Ý)�'�`Unb�w?������yo�Ne�`�UI/k�(��BZ
J�%I��~b=<�k*��Ӑ�q��+Ki<��������+��N"S�-�±4:.��G�Z#�+�`�I���)}h���i�?��L�M&���P��\��<��.�<s���̛��qՈ!|��\M����gӁ�Ӓ�!4��Uy8��J�;F��^&R��O^�'&�q�O�M��}�yj�j�Pf�z]���`�W�k�J�	L�-�]{���xT��Bq�z��Z�32��#=�˚)/��}G�����4N��)�\�\��iDR���@.n^�\d�L% �0��&����Շ{Ұv��1�����#�i���,^�v���s���(���tH�=�l�/���<(JP�m�/�;[�c�BɭM����/ZP�8*�s*�w�߅&�����T�0���}�Z����4s<@�Ϸɠ��)ֱ�
^���(��mX���`woIk����I�4�3Ol��M0j>�!��.�����<"�	wK-�U<$�J���"+TX��qn�isyY��Wj�=4$J���4i��v�p�=:��Au����:����Rf�(b�w�VJ�܌��i�5ȯzDvl2��ZX��ciK��l���V�9��!=@��}{mͅ>���nP�-��l>r�|+kZH_�&��P�OI�tb�IPk���5D����\�Z�P ��-�d���r_A|Lu��.a���и��4p1p�Bɫ�_�svF����|�2�K�m��c$�f�c��w����v���s�-��*;��>��p�h��!���~���qQA��l� ��6!V[�I��1}8�jwL�_�A�C��C��e�L�e�E@����b=M��!^6�[��� �,n���^�Á�.�<2����:
�������c��p8��ZEEs|�U�kmnM���?�~�5��8��H�Ch���~��R~3�9���R�����8�*�t��F����8�7u�dQ�q�O��e
𣳤�R�J(��Hlxa�� ��FaUt�iF��NY 
��*'��E�Z0���m�Y�:)�$��=f��,���� �y6\��s�푝�"1C�!7Xd_՛�Q�@��BVIm�;a�����{���_�t/Eш��n�.hK�4�w&�0=Ww���c{Y����/�����U��]>���ɟD���:��԰�LTK
�T�%N��#V��-�he���!�b�B�
��6����sd�?Qo��Z[��oˌ���W�s�l��V�U�F2e�k�˂� l�r�lr$��s���Ug�6����$��OU��	͙-��)�79ʝ�p��d�P����n�9�A�:e�S<ё��.��{��g֤N�h_���I�G�Q��x��_�]�ޞ���(�G�p���^����_,�A�F��<dƇ.�>V�-bR��b'mXuMs��x�h��!#��UpqRg8��F�T[Y��.�ee��L�|?Л+��6��`u{^�j/>��}�̈́ǃq�	���\����1XS��0����ЯL9X�i���.�,m�r�}�#�?��ǣ?��A�w�Սk�d2N<±�t�2 �*��擋w�'�<x��.UO����:��=�4�+���K�#�|�0-���h���Q��i���ͯ�Nؤ�?�
�C��XqωR�<�@owJ��Р�iJ�`�@�5҃	M����QGW��P��B��^%��~�QH)=���,��F����8>��i��٭�v+���a����@Pg�.��x�F�b%�i��� ���=�C���/z#\S��1�����������`��������_��q�	 ��
��NkmG�=~P\��=��L�-�\�i=�cGt ����t^C�C������<�ֆ�,x�|Q{�To��!��)Ζh5a[=T�t$l�&��>���½��g���P�n}��~u���0���# �
��Z\���O�'��G��_ I�y	���՘7��f����1�D ��.�kܻ��\��R�x.�dK��i�6�no�{1"�7)��q����	;�4�!�8*J���L�滮��8B�Ӂ1��o������L]]�����2)c;Vo�r)���q!��o����#�\}�R瀁��/#m�VF�w���}k���j�����906���?����b2�M�ا�Cb������"�h����qICc��h��xWu�h�Gɵ��]yvtX�	�}ɐ� ��	'>�ꧾ���z_W��w2����Ⱦc�JDl���Έ�M�#��ur��*��R+?^�Ɵt0�<��{��̣�{�}��
���R�KT�c�5��qHA��뛆��Ǭ�5@��C�����z
F�R;�98�'3}��jg��|Z%{> q�ig��q�Q�&�#_��KvR(�D�q������9кם���@E�5���,X ���&7������8|�BA6]BZE᷻�|���ϣf�d����l*�8�:P��+�aX����ha��!�.t�̞l��'���~���D:�˷�RZJ�,*TVfV�!��s�:�sb���&}����L��Ƅn�G?F}r;z3bۢkV�B��8}@p����([��J�N�Z���q�d����D�x���-�+����z����%�+�S���O�����;CpyZ�ftѾ�= �:ÎO�<YHhG`�&��H[��'��s�'�6����?� <$���T�K�|	��H�1�ǩp?��]U��ڭ�3T���]�D��D,���K�获�дjܚc�2��)7P*��nc7MM&a@���v�=�?fg7���3T��"�R?Q�8�I�+���8���8�&�&������	`2!=	l�)�O����t��i��E����9$��� �S ���8`h���1����$jY�k$�օ �����]Ǒ�6��u��tZ[н�#Q�:V��8���������fV�){|=5�,���M�919��+fds�8���4��n�H,�/J��?��@%e�����=�T�evs6'q]4>��ҚZ�§B�`�_��Kr�+7��hM��~~���n1�#k��(�ʑ�!��n-�^��Zʍ��S�R��?���E��ߤ�o� \1�8��t�/B��fB��nĦ�¶�b]�kza8�x��?Y?|��N՜.)�O� C�H�`) �Zt����F/x<�z�@�g0�4�F�08���E���B0��ʟ�&����7�mJ��"�)��m�G���˼�f�X��n�C����?�ͅP����-m���,�}߫K��%3#�09�����x�@�?�y��Q�8�eE���
/��+��MF�w7\�k5 �ܓ�6�)�un�65nBiMc��QI��s_�"	W���{K��=�o%֢�쌵 �][��KȖ6�U����yh�)�s���# w� 9_�F�L-�K���arv�c�g�pL�:�aU�����ퟫ���-:�e/:�M�c�L�q�*�xgs8�a���k�
�S�j`8n�����N?L��A��ԛcmH�<%ݟK� �i�wE�����-����
������:;}0yBv����Ai�_�N��G�4�vJ��T�վ�7\Dyx����ݡ��t�>	/##� ����������s	ߴ���z�<=�z�ɻ�g@I�8P_�`�� �:�����A�]R��'�3�N�d*�����Pf�����pd3��8*r�喯t�T?&�6�;�jx���7�U V+�^�]���LA'Z��|�3�V��Ꝇ?p��4pC/K ���CW�d����!�s����WR4�T����U|�}gZ<��D_�������V@3�����i�GH� &��_�?�p��^����aoW�C�ݪ�yop�+)s�.�h!g����A~��{��:uF�a�B��]�Q�pQ��D�&����eIi��WYO�����/�6�6�`5��Dh9��Ό�����e�����X��
�g��Dc�D�߼5�^�@c ������#�������2	�����n���Uy�$Hv0H)}́(��BvD��$L1�5tt3�a��zG�<��2�U��9�n�9���r�˩R��Y僁��/ɀd�; 5a�����s������������?���wl����Q�*���ݲ���REh:=��"?i?,Jϒ,��)���
[�$�@b̢�BjM'�J�Ǆ����뼌a���^�F?�^k�ȅ+;�v:�=�$��yʿo�_	+�s�����P���q���'9\L���M@�ι������z;��P��]n�1�N)kT*�I[���	ҧ7����w�엌�2��]��'��?����U<)P�>�f����'k ���^�%�����O���؟S��a����0
�I;�MD�Ĩ��� +�S
���20�����%�?�\��>XV�e�j��CNv�J&t�o��� S=��k;ȅ�}�3d�rgwrv�Ru��tUd�	4H�? F��iT�3�U�G�1��[��Թ�	i�D��#�B�3(������=N��'��c�7��iɁ��F���ґ���dlW+�`���]Ӕ9�0;"���������_f���*�DQ}$�Z
���8�1b�ѫ�3g٤�/x���&m�������0�W�f�p��I���(h�2�&�A�h`��R����ײ6X��;�_�R�ǚ����oR���L�=��Eo��툡�]^�WAG�"o 	바��*:9�������Z$ֿ󮙛����J�g��:�XH�Ʀͱݱ���ܽFE9��6���y#������?��t��-3�ȳ7�Ļ"P�t�P�T��3}����dȆ~��ʾvIV��"��N��O}1)�9F|%���^.����z*�Lܵ��ε^�F<�w�����}���_,���͉u�KEJ�$ٳBh�.�b�K� /櫠��ܨ�:O�4v��c�a�fca+W�ՆD��wh}i�Z���9��U�'R�L���I�5�"�Wޛ>��r�$��r�v�?����nh"��n#�	��K�<���#���z��<����eA�� �]`�o%�!nȚln�k��%�9d¥O�\��ju@
��u�=bķ�RE2<��'hEZ�e�N��BUD˽T!#ժ(l�h���l+�az���1+�ŷs6A@���'�owA�������WH���/)����!� .�y٨���F!��l��H4h���{ ��v���[f��K�5!��/+ΐ�T��{�}���u�2$���g��"����4�;}#���"�U��}x���?TmZ���<�<n�;���.guB j�д�t'X�����{m������Z��<�Ta�����J5ʪ�2�� x�;fR��j�7�����g�R�6���u;�N9)���a���K'B�lQ�'�
�1LBhܙȜD�bN��%�B�wLqR�V�|��}/U�n\Y���J�����Aa��_���tr:~H���+$Msv�������]~����*mJ�!����;913Q�I����$酅XR�������� AѸǀ�4$^���+x�	��<&Ϸ�mNX>	���d�	eE"�")e+����󚞗�� ��J�
��j���Le~���qغbЂsG�T<��6��d5���d表��i�	 �H�Ltf ����SG��?%��-�UO��F��#�阺-9���V���A�ly�o����ل�$w�,2+�b�#r�!Or�Q8Ɯ�X��[���:���dA52��/Q��hX�D�t��FG����$�L���j.�:���6�����4\�IJ��F9C�]����/��"�o�;#l�CЃ�q@nϾF�����*Ý�ҁ��\�k1-]�T�/����O�o�O�`�M>,�/�4k�ꡗ�i,��F6B�:�Q�L�GIpO��Oj���+I��!�.�0uScFC��Y�G褈��X�p�/eW�u�q��ڽ������uI��*TC$�S�{�E�b�`	�UK�l$'<�N�%���qWO]����E-u��"aø�:��G���i)+U!����W(�B$��#.�ׄ�d'����;��(	����ǌ_�c�}s��J� ��/.�zv��`nL�|s��{
�����X[Y�{wX洀�30/B鴿�k6���V�#5a�=�Lz��  }�J㨉s[��uoA�!����l�
�y�H���핀���!+�HѨ�U��I3Ĳ�k��;�g^N��۸ॾ�F��מ+nq���z���V�~ѴF����]Ǐ�~��.&2f���LLY�mx�TM�U���<`l0������ˊX��6���c}��]U��M��է�Y�`������( ��=Yó7t�.�"Lh�f���Y�鬒F��R<4����VT��e)�:������ߘi}QX|�ע��7�֟{���^ޚ�׵K-��,-������f�O�4�e:8����A��){?��t|zLL��giwR��0 6"�U�%!��ٸX�A����*����ƥ����
=�;~)|`O�*��͹��59�۽F�\��V�ht�A!Y���'_
]�����:$�ߌ���0��v����r<(���)%��������&��<L�;���K�$Z�&:��=[�S@���~�O�f�����q���.^CW=
�j��s���*��j���O�,ui���Q��"f9����P��Ά5�����=A洉��jd��"�?S���E�/e�IlCGc�C��>��-��fJ��h<�
�o�	�{M�TA���/n�3Gb^��R��E֧��ʳ>�aB�e.����k�ox��j{����"{H�����S�o���,���4��-{M�O�Ȕs���v����gX����V>O#�K��crE�˧��߂��hA��w
۶��5���Pa�C�(�[l�����װ��G��f܎\��Ҍ��N5P����N�7�@�7���I;��`L�g�s�|�,g�s�љ��%}I�*4��x*H�.n�C��d]�1��X�n��zF9�
�����`;�[S�2o炶�����U����Q3:׸�1bϼ�z\xҽ�����Z%��^��/)A���ej����O�t��.��ic|R�ȅwVIձ=Y�����w*������'^5�����N^�k��"L?v���sF�̖N� �b�>�����P10u����.J8���I��[����io*|��KO�}��:B���	 QCZ��b�~jӨ�8h����a԰:�_�++�����R��F��f��"��gl�ڊ�%rjk�!���>OE��鬿HƔ��Ȑ�v kx�w��&s��bL�	<y�(���;^���Y��jmi��4r��S�CfV�э�������BU�Gs�'\�`Y�w�G�X��ݣ��78��0���
�u���~Q@M������R�~"B�	ܙR��m��P�nQg�Ef�*��&��Fa���0���Hj�\�+<�B��U���US���o�%G�]MZ�A��������0HR����X�<��r�y�{��#橇��:NLQԀ��m���=mH��)��7�R��Ԁ�I������ ��Ѹ��!j���
��~������H��ӱ�����fY�0.%ٌy
��؃�")�Y���J���6�6䑺ս7.1W��;���(|A���^���6�-Y*�ª7R�n�~���y�0�[<|O,�>��j8���/2H��Q#j�^��|�z���N���D{uvt#�I�+�
^���oTs���*'��47�=���7��ݳm��xS��}Bz!�k�2y����DL��b�c�eU9�پ�`��<�X�P��^q2d�!�br/�~4:F~�K��H.K6�K �t�n�D�x��'�`��&�}�?U��<*�,^�dm�;�ۗ:�|U�����U8�\�o�q����kN��<�k./����
��L�Xg<�%N|�� w�w�c<�W�p�T3'���菷�_��Q,˴&Ƅgsʈ�o�:p{�HO���L�G=��H��m�GVue�N$�79�����i]�4�a��9�=C�)��h3��7�S2��k�*����Ĥ�?�x�7����޼�M�٥?euK�o��[�sUX�h�@M���uQ��O��6���}�I��.�{8���]�=�����ܗj�VU�G��
>Ijŵ%�g�����`�"A:������oOs:�uO��'���e\ƃ��wr��W���*r9r�N=�+.��D�f�@�m'(���z�+��1�rB¥���T�cGO�h��r%�V#�1��[��rHZݳ���0�{c2~�;z��w%����,��ԸQ//۠�:�\E�������i�S�jL5w@�k��tu ������R'���,�?I�S�Y�N��gz���6������S6�
����X�p��9Ӎ�+@Yc��i$_d@����/9ք��1����W�3[9�uM&���$�^X50���Пfr���DTP�c���O�$��_�e$>I��8Dץ�G��r��y�� ��}e{� �E'lr�<�J?���"��m'Dt1�*�3��S���ᠠʱ���3=&{�#����<zz(�v��8���66&�6�SX:&�Z�;TZ�3��ES�D���t~��(�0��?9���N*�{���A���~�$_:�in�XxKA��#��XK�O��&��'��`30��h����Īsy\3"�ݏ:�`7�T�/����n�T�O��>%I8 E�E��8I�	�ꂆ�]��CcRE4��#���D�)�p��f}k0�D�5����ؕfX:�XpZ�F�t�Wܗs����K����,t�j6�:T���8���d(��G�F�el��IC L�����[R�u�Ǵݙ^�[����U�_{��0��8i���S�f�%��~�L_*�K��WH�"nww��:�EA0�J�
U.��>�{ e�CH���~|�O_�+r�#�ιF1�ěWF:��(�/d�����ݰn+��
��I�eBl5<R޶"1�G��`�DP,^3�Ԙ�:�rl�pco�����	�����i����]p�z��-D|Y�@:C"�@��@(��\mT)�1s`Gւ­@=v6�៍P�kL`�_�
Jj����������}ʳ��^� V�a��DXOZ%�ɀy�:{��.��$�G}�z�u��.�D=�$oMa^�ؐ�v���s���ƩŶ���@�G����s��U�ň�w�G:��R"�I5��.�� ���j}\xF��$���6?�R��1=�<`���p��������m]*�I�D�ܲ��ǫ٘vr����Sˍ�_x��Y����{2��*��4�\��W>^�����`��5-��]K�����N2xo�`O=�	=�1���ܶ�-|��@�[�!ι�G�{�'�Y�J�m�Y��xO��Ew�z���'y�4�l�1��c�H�V6��A��.%��a=/H���#o�� ��kZ ��f�E���7X;�5/t%l�Tf!��fp��͎j3<���?+�'ݻh�S{j�8��P��=;�C������u��_� ���@�k�_�,���̍ﭕu�8��^K�@��r���%��������s��'71����OS:<�o3�]�=E��D-�E�v)2��^VYUB���6F;8���Q�v�L�33Ҧ��[;�������R�c�Jđ5F��n1�MM��Wl*�*:���=*�6F7��ăΝ�ed0LM�B�\H�?e2�Q{� �ށ��c$("�a��:|x��bO"�X��M�п���/��,�%�Vܢ�L�<�(��E���!���1�{�����h�燓��DE9���gȓ��Ѐs0��z1e���Ն�|=/I���i׌��*�S�6~yk~�d�U<�]�Vr��<�_��E���$��<o�	aBG�� ��
=�(�݌�b<�R��빖��n�pKb��m�������9c�f&���&�Z"c](
�� ����p4�KVֵZ��N�5�X&S��k��
2�(�����<�#nr7����G켡�m��2�"�ײ*�w�⼁��K{�ñ���1�h7_o�@�G	�j�E�|6;u�+�%����+�q~�~z@^�$�rUy�t�T$8�����Y����o������g��fØ��q5,�����Qn���i`�
N�ׅ젿��t��!�tQxIL���4�xL�`����SL�� c@��ir-��+C�p[M�,�o!�NV���K6/���22�H�D�Eamƙ�%"k&j9YЖ��Z��Ե���v'�� �"���F��U
h�z��:Bj�*UO�=�k*c;��B_b'����&�r��Y���S�⮋���]�\���:��� �|G�>{���@S��a�p��m�:�Q}�I
��ͤl��ܢ�� �kޥA��涕�.�� �q�T%�S���p5W@��E7v�!b���+���=�*Y�b-F���HBf��u�)�f�g�t�a= 
 ��pg��9]���'��W��J�}�[��\�`@���&b�n���u�二䧲
�t$�����K��4@;pS͵_�¨<�ԗh��j��i'�iM�X|8�:s(�ƽ/��%j�Jzd_��l�={n��wŀ�'�(�����~{<D\�����K!���n�,-�J*��P>~]�տ�odh��'8���b�]��D��l����+�"/�;5�f��`4��8��
NH���0O�w��φ0h��Ԏ1��E5ށ�����_������x�t�τ�D��- .����9�3:\'�����.'�k(�ԃ�秌��W$qtY��B�؜6�O/�΢:|�3g���q �GiHR+`rk}��-a� _��n����9�����ΎtJ��[g���n'IFSQ�G�������.)x�104
���a�ԗ��m>j�����/�^�]99l4�mlO�$�5'��#��ih�<=��tr�b:	���ۢ��F�q�։1��I-��i�'ι�����K�p�YhT�9:��N^ݕ;�WT�A�r�,��� 0�D�
�ݓ"�P�����\��;R���%[��48ĵA�1�Z䭪q-����!��D�/�ްl[��������񧃹�����X�����"1Y�.AX�}����ϟz0�|о�x`T��颶�YD��b��
}�;���%�"Au���P�2ޗ�ƺj@)0H3��;��16f:���Nd:t��zoX��|緒�xm`x*���r8J��7k�3���K���m
q�Χ����`�W�,�����0�ٮL��j��v�5��9f1�Us��4��~��n�A)���gT��c�ǹa�v�+�����{����V����}�������Qǃr�ཞ����4�+K��0a$
��rNSm�4�씒N�qP�~�wW��S�2��P
�k!;���o���yTtB'��.���ٱy��1���2��Az;s�3�J�`�
�F������ܪ|%C�H�W%�B�"��O��ù��,����;�d�������~]I�E�&;�t�Ԝ���9_���:��l�NV�p-�B�"!I� �?R���I#��io�^C�w"P碶�F��se����t�ϟ�(%M������N9�`(+�7�c��o�Tꁤ�.q����)�3��>�ї�6�XnI�&�ɏ�Ge^��F��ſ�C\⊾(n����꘼���.�# ��.y�^*sO=<�nv��
�GZ�`Q$s��ٌ��,$'�4?}���H�㽇�L�O�{r��J�m����ޡ�sKAK����zw�0�l4"�����ᐎ�����j���1g�=�5��~���7Ct0ɣ�Q�`�l|�Α��du�2&1�1�������d��iqB�Y��<S��JfJ�+��ä��Y��)W��\��'���qt�
����0\�^��(��B<�l9�rp��u����(kº^'n�j�#/�M�嶈��6w�X���m��&�(w����>�3�8�O�q=lJ]ļ/=?&��!$��V�\�-O���D��Eu�f)n� �r|E[�����cV�������NF��3'���ص�)�I`��K�����&e�/Y��l���O�g^�]�r�`˫��Zr"�?ڄ����苼l[��Z�Z}�8�b�c3/�qZ�}����R��K̫�8�"���|�E�_��2��p� �e����^7��_��q��Կ#G�Q�/3ݫT6� ��J`�)Po݆9* �㋁"��I;��V��8|��u#$����1A'��)�Y��4<�P�X��1) b'���w_8�lHXL��g]�f����"Tk+Yc���p�"g��s�c�5tͺG����W�mOȦl4�\F&g��������V��
|�|�R��+�]�u�4� 
��I���V���>�_�d&i�3��\�i���n�͎�mS ;
ꖬ�'5��p�&"�a,]o�&/�_Em���,����t^T�.�@����B�=b4��M��	f��r��G����]q�5��6�I7:�_�( Q�:M W�sz�4X���$X�,pcK	-c�غ�k��x�D]�uk<�k^�Ң�x����aM�������	 ��,�����ƻ1/�I��إ�{����q]�-����gX}PJũ��? 5d�|#A�h�з�e1E�\�ߑQg՗�Д�D��>=����/��p�r���Գ4�y@dx�������۝���6J��6��څu]z���c߈��eM�	�
:1�C����;TrA f�/�ZW= ���В.]��{}&�-��"���dܥy�_��/ر�d�7;sf�e��Q��TW1�ɫf4�3I޶8A�:w9 e��(���
S��*̒�:�+r�Q��2��i/*1���w�SP���Ro�b�Ή�~S�aQ,�J����ż�����2�uQ-�
����C��Z�7��V9n���U�37	\㳹�mVbB��yuJj�)W�r�<M�G�^������Cc�y�g w���'7�q{���:z��/�
-��M{�����c�,��j#)�y���Fy�����s���8R�η�B��Y��H�TS��jR��^{��c������:5�M�b
�~�����Z��63�V�B[@8k�� F{œ�ɿ$Dr&������7�
��kfއI�3fN������U�@u���Q��*�=��E"��;��E%oJWZ5��`Y��:��z�¬�'������G)Vd��+a9:P�Al���TGd��&�몉�n���n����E�{��4ǆx�~-���e�!�㞣���I)�Y���x�K!���F�Pb�Ug���ܥqA��XYÖ��?���i���Vߣ�#pri筡$)Y]�[�J��D:�S\���/���OBĒ�� ��")[,��A��*�xT�����G�Ff�y<�\=/��uƬUD47�9�x�R�^�&Ҡ�}��V�e6���5��
�F�@3AFl{?Tշn�Đ�]E���u6��sHc?�����	�X��G~����t%G�,�UlI"�1��\N�e�f������J|_�a��k�����1���&�;�w����5�%JGI�>���b*>*�|��9��6E'�P�D�qG��af�c1i�؉������9 �����iE���l�޼�g$�Sa0r�ց`����IcM��d@�S��2v��D�ji|҃�٭�����Jq��#��}*-�H�f��K�������̭?��)%�)KR�[��8��<p;��-�L���6�h�%$,R��,5�i�ND��|$PJ� ���x�59)��j=n,����y�?laևa�(��އ��l�r��(�.�U^ѭF�nf���w�S��OnZOo�*~Q��N��_�*�>�D��eH�Wy2dH~;�����&rr[Nc�M��'��o����X�3ְHF*�a_z�y��&2�9x�pA��ȩN�9;�o)���n��:����!l�E�.�[�Φ���6�~��be�Nn Ӟw[�#����<�[��	 7�#�hUJ����N嘔��V�Ѷ�)�`
L%�=U%�(���n�[�S�����A�S�~���^ݎ6 jyM�:|��\f�����QP*oK"y�J� \���'D���	��c���E#�|A)r�
�}����(�h���ʨ'̀f��r'܌��;��BZ[�?�*������A�A0�?�ݦ��۪��i��h�lJ1�����G�W�����`b�������R�A�m��L8�:�۰#W^<�5d���U�pb���TW�b��\�6H�X)��^<���v�(R�2E�C{?f�����}ʫo;��Ÿ�hHnљ�p�[������^HF��E_�~�M�!!qP�5�R����ZFa=.愮�ӑ
w�\Ha��df�8M�Y�ĩ��[J���ܞ�-����d�ؒ?�����#��N�vJW��`�~�?O-�����@�j�V��miK� �^���3�Q8��89���|ӑ���6���v"�	�3%H*?K�^����I�̉��;AoW-7�T�2$J��A�C�@-�*����gʙ�#�V"=&R%��Ń�����#N@m�s����/e��v.p^�k�-���P��gՕ�c�u>�]���EƩd�7�&�l����| ��o/K�p2�U�*�q�.���L���H6_��7o=�߯F��P�jф�w�Q��y��y!S_m+i�ٹ�����Pw/�4oTL:����9S�݇�)}ΟY>����yWZ$�Q3\��j��M�m�� �OG�H����Qo� 	�t&��1��x���T��,��gy־�5s監�1�A���*k!6;�m�6Ƶ�-�� ]�X�N��8R�3/c	�yXN�携����	2���QD*�M�Q��2����<��
"@'$u�2�z�1	�K?}2p������U\[o\��q����[iE:�wx9p}y>)�c���G�fm>�"��0�jt��57���x:��#N��T'+sV�~��Ԩ-a�0��4�T���8��ы�����'B>�ZԹ^�^�5��--%�1f��#������nQ7Ġ�Ys����'` 	N%�s���ׯ���>٦5�y)�>��
K�)���m#	�ׄj����h0I�z���8�t�ۡ>�\hk�o����1���!�;�3���J\`��E�=�'��$_�T�U��=0.��[���w9�����Jy�h�����仹�;�`oz����̬�8ā�	肂�@�k�g3��Az�߁�6I(߶��"��g�ߑ�_���a-�->:��XF�t)$���r�0B�����E���1���J�-�b�o]�n�׃�+��^�xieI�K�\^D亪�F6�~�Vv��"i�����1�!�)[?��
L�Bh�����g���}��$�&�~�,���s@N��\>���_<�X��)wov�>�*�O��S�E-��vşb ں2B�P�ڢ�V������9���䓱�8�s�sF5Z"�]�۷�C#��{
���$�&YG�x��3d��O��`�㺨%�
%�3�=��h*� ٹ����@w��6	���B�/�&�eN]��4���|��|`1���-~Rul��Qc?|F���Sy��M!(��Y[��1vȁ�e���(I�8y�V9_��	. �;ރf=��Yu҆N�YSY�"d��fJS�v����bR��b
~c�H��Nv;��+倀�.(�ߋ{��&����.	[JO�5��H���Y�QeJ�������-jM����=r��2c����䗏�sct�������m`h�+"as��]�fy�l�s���-�D�T^7�P�=G?-_�6j�ýؖ[T]0O�J���h��G�t�pI$���x�?�oQ�)U��)�	���I]���K��o���Q��nxp@�~3�rH�^�g���ö��EH1A=Ď��v6�1�b�����g�6��n�G'_�"J�t��-�({��l��gUc&%��(
����m�}�dbw|W^0��?y�I�0��G��Ȑ�`�EI���G��Ԇ�1K��P ��
3�r�������{rC���������Lex���-j}���^C�J2\:TѬޏ$�t6�q�`��RI��z��{Rb��m��s��6�ݤ3��]�C��M����	�\��ZT�-H�Z�{b\ï)����|�',�Nc5��V�:���5�/z��	��@�T�ݹ���UYݕ�+N2y�A�@-�y���B{(rzv��隥,*P�[�b�F�ZG��>��.�L�ߔ���W��f���(�VsZߩ�f�@>�V���w��,�9��Q�L�@���Ìa���n��I1��cj���0h
��<&�4x����r����x?w�M��h���s`�RCM����ퟳ�]��u�p���y���lGs]F�47ȫ�z �1k�^l#�W���O0�o��;�׾�q��n˔b;�|��Ҋ��l�z��_�q �Q\V����8o�"��}�������1�=Ż��Lʣl�D�o��m�<fZ�p}����w��_��+�퀭��䢨P�íGbE���0�|��ر����
�MrV䣛2��_�r����a�8jXa[, <�Xu��
@�Q��������Pr�ZgN��͢��,ݏc�c�>X'�;Ś`F,�f=ғ��]*n)��+�� *�t���W��OA�FY#����5��h�H�o�n��O�TG�c���U�e�*�ҰUW6��/�MZ�fͰr<�d��a?$m�G�I�N��ɀ��dB�7�� 6�wr1�e>�Vtn�/��zy���e�q�&��`���+� @��Ѝ��TY��z�X���2�Gߎ�.������M�Ȭ��hS����i�k�Ͷ�5|s5T4�o�݁r'x�ϗ�W��%d_�fs��ʡ;�0�t��Д�PZ`�J9\�g��}Щt�FW�_��C};4n�r��]j�0m��qR�-�T��`�B@��>t�i�jޣ�e�doc�:��Wh.�������=��X8��>9ږ-�XE�P���nP����|{[��n�?m�mg%��E������g'����6�6����j&>5���foL�����j60��()ɑ�4�_W��I�Gs��5Z�����$J��J��P:�zGG�@F�̵%u���z
\�R���G�l�E������^'���./3GF&Æh���������.�����t�p^�9[.2>ϫ��1m+.o2�6�ܚQV��I:�j �z��ޠ8��hr�WHL�Zx�胙���/�¿�!p�q�?�0�K4t��v�a�'�������s�d-�F\$����;byW8�"����y���u�w��j�'���gcH��M�]��?+�OJ�T��f�#��y����.�R�IF�܃̆3y0R�W����{1��ɣ
��|�@q'���R�kZC�g���:�0�4'��(�q�*IYS����SY��'V�����:�0X��m�?Rg��56()p�V��%W��dXVd���;t{�\�[I����{.ٛPy��#�!^�8}��B�C]'t)"���MU�6�
gFe���b:�W�i�J��H%����5B�v]|Q��1QlJx�_��>5V [�������'���n�-#j���&UP�5�d���#�*RS��2]��D�Yl�>�-q ��J���QU��}�����UM�,��*<Lq�@E���5 W�@���t�����t�#,��mk��w|a[�*Š
���� A���
�?���>�L�]�Im�>T�;����o�a�+ ~8z��͌<e�x�K2���J�:�ږݶ�]���1fq��59F�a9�K[=*c����9�:�ՙ�_Ѱ��*ڋ���t��R�gI"�׽��xӑ�[ޫ��
�pC�b�Q2��8S�ZrsZ[�k�X�?��	*�'l�"�";��*	b|��6�9D�U>�)m�3��cٜB���J��a|S搾�r)�x��f
~���g0�"Dvj\����$z:�ՙ�]b�lET���P��{KІ��f��̯2������8�!��kĪl��9dOd��Y�\�����bx����NJuQ�2&.W�G],�ha���KN�w@�WYp/D�c��Q����g �$�D�D}+� ��(O��ͮ4Ĉ��B�f������qԋG��?�N_�Q��^0��J�?����pt����m�w�D�[E��cf�*�=���܈���uր�����.T���}I:w��?B�b��۴����p����<g��^�<O��؛�6M�u�W��S s}�-�T���=�w��*�W��W/����2�ՃJ��^����o�+o�y�3��4���+dy`�v�{Ĵ$�-[�����n�����!s><*m_�+*���D���P�I��j8�GmֆT�M��v�'�Yl�Km�ݨ���n��n�r9_���6��E�L�I*����&
�ͦA2�E	�9TT�^�en���:�F�'��T^{�zPdb)�R��\0���.fS�l����{|�یPN7-�P��L���hf��(��y�gg|~	���D&�0Ѧ��EXX�(M��ڳ�����G����بY3i��Cܧ��)���޴��՜�}�:��ϴ7�1nQ�H���s䡒�����F�O��RA\G��Qu��p6O�����|����S��Ϻ�tȭFI��@����4l�I�����.���f$��p�p�Z�[��㚊�;H�v).�����!�o/����k��M@#o�7��c�;N���`�o���(��:m��o�(��H���D�J���11!��5��.�;-��x�b�z��P��:��I�o]r]`1�e}��r񟵾st�*�����Ahz<�,y�Ł.���HQ&Ev�G
z��;�82PG��U�L��ZA����1�i-����/X�v�2D�I^�>�:���Yˡ��t� ԣ��:]��{{-l31�÷�F}����x��/��x���q>�u��|���o�kg�{�CS�O�pJ�W��NZ��nLqO!r�r�բ(9��%����+|������z�;� ���bȾ]t7�Z��N��>�¾Q���/��57��k�t�(_*d�l;�׀�4Ơ��9��X�n�-��@�̪�sY�^���8/����3p��r)t��!"�W���܍S)��d��4�&�K�g���I�UFn����tøX�<C����}��e)Srrd-�uL�$��w{j�Nj�l���˧�8�AE����#{�t���vs�EUH���2�*9[����_vU�"��6P!��o�g!�ڻ��b�k�l&%��B
��O�K��Q����r�7�&�\{[?`���LM�<U!��J()�mL`�I��𰮘0鷧T�T%�7��kn�k��Q�B+U�Z$rQC899t[���+�͜�FP����ߏ���_��.�t�{7���I}�弁�;zR�Rl\މw=�~r��(��IJ9�U�:~�b7�_������E��zt��׽�h9fFb�Έ�Rx�*���1�b��c�c�r��%��Gp��s��>�m�+`�QK���χ��t��5�1�!Q�<*������~��.g'�OLb�缾�M{�l�bdҬ���3�YC�� ����!��_Ш�����JeBw ��eJ�q��E��­��ae4�[��G���Dm���Z�S��ї^���I�#`�;�7y[�8/#9yN}|Jl�%=a��쀑���a���p�0�
S�|� ���,�'��+Þ���y��{{�CZ�iJ�sɻȊ|�+_%�b��e&jeX��ϠT���Q
]Ah���,�a6�@SԖ0�n�l�k�%�V� W��=��= ����Q��W�P��N�G��/c*����<//Gv�} �8�eYr�LL-������Zw����$���̆�&ې�"�٢lkf���!���,L*�[N2��� �T�]����$DyT��ׅ� |�
^���R��C�B6:s֐���	 
Һ�f�2�7����?LW8/[�i���g�
H��i�?������ @��~��6���ڈ��ng獂g:�$ �BQ�wg,�Rtb�"��ey\��gy���l2:�)_E4.���U���3t!�M�W�p��0��k�t>�o��C��
�ߗ0`��^E^�����*'�^��>9Am���Q������c��<�,o��~<��ݚ�K5���l}v�1ʜQa4w��O}y/�7<rQ}e���	(�`/�V��H���o�}�9X����|�Xr�P&��9pM����.�'p:_i\ߕ*�ax��rZ���C/������śi���Hu��O O����Ă��]_��Oc���?3�d���@�ةh��o�a�f�T��^mfw�Y��x�&�?��՛��)܅[v��J�o�yL�~���c���6��F�j�?L�f�ݴt��wL�̱&��.��_�d��� �f��e���~Y2;�J��#�F���A[Z���s�DN�Q�#!�W0���|�3u;�v7������M�x��9�ƞI�g)tsVߌk+8��a?�m�=� �}�3�g�t	�g��}A��evh���u:�e"z�G�M�E�*�~�8��b�����j�;�y���:�=T�<ڷ���;|K�5elfn���)QV�~�/U _��t6"��p����F0�@d/(�����:o�/�W4���L�R��(�4X������e	r��֘&N��[�͜�&���|�孻�
k�!���þ
�Ά��B��W�m������Q�C��}�%7lv��K"��j�xMB'�����Z��'��0���7)r�R��Ʌ��4�I�`@�R؍R?!_��?qvqᕍD6u������4�3Ѩŷ/��>cN?���)d�)��(�D+Σen�}���Bƥ0��a�#�6��)�^�IO
�'9ekR��x,B����A�`�5�!ߦ��VZrM�I<��<��e�K 9���L�Z�$���
p݁�	�dd��нNZ܇�;�O�y����]�{|�l��ա[�,>Hj�n.)8"�\#y�����*9:��ZU���NVKe�??���aFyڭ�g�����}��U�XԺ/�s.�	d����$�l��E�-���4 ��Sk�lES(G���j�}��p�"��s��V7�R�<y����l�$QjA�#�]�cc2ף�	���1;R��p{)牢��w��@����p�eN�ش�
�7"j�8�^l��x�6Q�A��M+����!p�VF@�\��,]O��N9��yL�������7�#(���:���5bY�T3aCb[O�Μv&Vr8��m�S#gb� �a=X�kz
�;��T��5�9h�i��ܿ�1�񷶔�����!<f�y<�����V׊)�š�*�c<0|�����2��kB�7l�1��>Ǌ�x���1�&��4
�./ j�G��m-]� �ZV�n:ږ�/� �N��8�#���C	���_Qa/���l�z��v�5S^�u��b��Wc#ӹ��)���zd�h���ԕ�Õ��	P�*M� ��-fV�zIM��,�㰺�R-��Ͳ��8�/v ��Y8,s�e����H~j=Td�́��`6�W6����W�6n�gp"��X ]l���wx��@�B̤�?�T��o<&|:Н��Xz�5T��3�jU,l��D��I�G��>br�er6H�`�/���+���*9ۅL�����!��{� 0}q��s�|]Y�v����zV���E{
ht���t
��Rr�6�XƢ��)"
a>��3�l"�l}�	X������T/�mK�){��.6���Nvp?'<Sk	bn��`�HAH��/]'YJ�ڠ6B������Lm��by�>�t�%T}���^�/Mϗ��J�w����ua��:��^}��+��q�;hP�ږ0""l���,я���W��XC��D��n_�G�41�@�N:����xQ�G���H��[����4�R��Eg�P�9�u���a0�"�dԀ��)�!|d&�q��}�N5�(�.`?6�.����)���M��&���s���]�C���N�	��eG��+U>f1����Y�x��#}5��	����ܗ�rjf����B�<9:%ĔI�N�p�O��]󠈏�G���Fy���>�ɐ��~�c�a�����=@�o+�M^:��"����oa��%Qo���^)$�H)�^MA��3sP�4M�LPe�i�K�+(�C;������_�����5��)�tf�Y>��D(ispDK���d�SH=��^f�R���E�B8�4o�G��z�R�'�X��&#��.�O<�S6+�y����Ks�3���H>�YA�!J�-�  am��*�k�e��8�i)�> }U�P,4&���xZ�m��u�)U�+)��D�e�һ�Z�Y�A���L��<wX{��]⩴�I�=L�
j�΅B�i� ����j̺�V�3��5�:��\��q���{��sB�y�5�+��&����=ug�ݷ�V�o>`���wיN�&�Ѩ�"����sB����i)��/����9�I�ewO;=��>@��,��[j�!7��	�,4iѰu�WpP��>�>ĝ9�C~���a��'T� k�l�L�J�t�0�`�$.4w�@R S� 2h�-������1	����J
���4!�M�ш=f��0��{�d.�S����n#�)w!n�vNp�u��TEn�C?�q�� [��Nbb���B_o�����Y���%�sru;�.~Q��"�}�4<)o�=�f.�>�J�*�p�4y�V�1���"X��O�)�����՟���&�Y�q�?�`��F��lڑ����@��PN�3��i�3�E^A�i��[ �S�e����T���*!���1���)|G�ĂFt�����Ƞ��p5<�\�1d��#Flo�d�����,3I�����yx�SF�����2S%�H*��j�e��Y�������ӏ�y�K��8u�u������2θ�+d���F.��[��a/b2"�݅FG�C�%�kNrHY��P�nG?KII {��F�eb���>�����PװF1���%�V�q�E��N�R� %�"2��~�t���;�%e\3�>�Ζ���t��%+@�P�b��ں��ٚ�k�M�^��0�5�z ���s�~X��%Y~�c��w��j/�%��\�������'�|���6Ni���e]��t3\u?��AY��w��/+�A�m�ؤ>�:�P�WP@���h�/��,��q�|��)7����B�!��ǈ��~���߮�=�30�d{�}�B�b�8T<%lفDU^``��Q_���T��@�c�>A�~a�9=��h,4Pf�H
�W�
 ����0w�� 	����$a�%�4��%JT�(@���?1Y��p̍�yz
O�T���r�b� ZwPQ�婻�Z�B�9kN���G����!_��V�^���~����,s]�:s=�A���n�6^X3�1k�.��n�.]��w_����yT�d)�$�z���\�$ɧ�=��|���NN�9�a��@�sZ�p�fEK~�lM�b�1�KmvO�fJ�H�j��q�v��Dy���L�ɦ���
��'�lD�9�\��ӨU����!�@�a<}��N�|rI0�H�۠ f�xVfr� �>���-I�_􇯴�V�d�e�v���#�#�t��}�dd"^Ŧ�y�^ɶ��(�c���0!?kx�4�J�Dn�ށl��n�E��(x&]�:E}�E�οb.F��?���̽!dr�ƺ���|S�q%)�X;
�����ya��b}*{W�愢ݯX#�z %��U�t�$J@�9@�ݟ�Ra��Z�����>��أ��FM���+~7��\�>���|0���-��J�B��t�8*�cR�4�άQǈwH&�\��(C@�]�k��j��
�̻��LiQ�{��
%��nlxL#�DU�7r��z�r>���oCةR�j��`x��-�\16�~����2gǠ��!���wW-Eys�wX�[�\���ޫm�UG5p������攉V��D�m��6
1��O���������pV`�����S���=����ė\���d���~�A���S��l�/Č�)����Q�Y������c����ǥ�Z�˴�"ޛw9�������	��h�"	��SU]��YK�|؋�L����|�U������>��W!�	��p�̿A�����GH�_8R^,������-�V�I�0X�἟_4�+]�eۃ��43k���B��`�g�[�4��4`�z�op��'��&*y�T��IF�H��0��>���9q|�}d��J�ޭ�֫���$�0����T�2�Ї̈���sn�+���]�@K�\N�WA��	��ʅ`���~�K|�����Z]C�Wf�oR���klY�D�H���^ʯ��?���!��Z���*"HP��z�K����r��)�ȫ���c�����j�������t��dϠٸ����x��j~�R��97wJ�E�6�V/��.��Z�t��U=r�J.�.*9E�4��'q͒7�����P�a��՛&z�A�C��k�m�y�2��G�ľh>GɈ��퉲/�g����0�+w$O(2���1�p�{�7�F���G,M]��pNbFM�Bw�O/��H?3aAi�8�=��&��K��~FX� .��Mr!N�%��{Th�/`���%��}�y��k8m����"{���Q���PۇYP&�-n �p�R�8_� �l���hqY�|�1�y�%�R
%�ʟ4�1+N��Q&���^�������l��^��p�_{�B�������Kh#S��l��"�,��u`sc��<�v��L*��^����h� [�~���P8�{Z��� @^*�a���Ώ�F��w�C3Gz�w�+)�����[Bh]vRt���L����г�QL�Z��P��a�f�����^��ĸ�I�i�jx�-�GS:shB�s^����jYb9��Tfp�F����es0W�l�"FDG�F�QnD0�n��M�j�*��.A	(qj��y��O��z�e��U��kp�dE$�$�q��J����@��=B�4i��T��Y�TnBHcO�ϠM��Vd�
�O����u+	�U(�/���u���L������%f1$�92��JMG#�^�g	����뱛��3K��� �\5=?!���ޞ�r9tO�]�9����*���N�I�(��N@���eϸ���k�*m_Q�ni��s�)�nj/W�ة��}o�/�����G,�!=�K}�x�7,f-�
'�$m���q�Y��e۩����}0�u�E@7��L�f{�1�mIr�1����E���4GT�$X���ڰ	��J%,�pz��XM�qRJZc������b��/V��r����GC���6�ka�H8ݗ��a�#��\6r߯�6�B�J�#�]7�%YBW��eSykoTb�E��K�>oa��[�����r���(�9�O�>��/�������ڄ-~���	ĭ�cɆ�0?%��ʪ����3�t蹗�`;�����.�{1L8]wM/Y�-(XA��7��mo2��"O�e
�a#1��g��vy�R�'�w��sы�&,ն��xٴʻX�t��G	]�v@U���5`�����k=�/n��~�J
_��ņ�](Y��q�K}l�O2���߂dûDy5�N�:k��<Y?>�B��N�,8��]��.bT�����	�k}Q�gPf����#D��A!�}[;�ŵ���H�Z9)e<�!�ҏ�5UA����"���@>f$�2�����r�s���,Y���ܟX��:$������؞�|��g*�[��lC)�!d����ܮ,w{� �3�-��t�
D�?�
��l�SJ�\ި��[��5��.�F�w�륒e�����+��K�B/�����1%Ŏ}�N3�΀D��4��Ņ{Ж��̌�SF�� �q>�%�(B�/���B^Kȷ���P*�NB8���"����k|����x;dTd9k��[��H�]Ò��,:���!�|��F���TwT��,���g�����c��q�5���ٙGuY���������.ф��q����c�/2���}���vAxJ�8� f�^|������Q�e�!��h�v�a���l*�j���^4dW��X���9_�IW�����)�Mk�}�ɽ0\��X��FJ��`�i.���s�g7pk�z������4qSHV���ɮؐ�m��7���sZ,�C>�e3ʇY^+�Q�I<z�1�f,��i��qL �X���Ǐ����f��r�&�T���:c�kӋ;���r�/4�]\>���Vt�)qCu��4�P&�Ͼ�f�;�`t�H�K-M�Ϙ|5Nz"}&��Lf����S)����p���Ց�k6��E�ltOk
;��Ӎ�M�4E�/	������fp���#�'-�'+�i%���@Y;������tL��2� |� 'E�]p&�ˋd!H��4ɑ���"�5�%i�e(�'�_!����^:@���c}�A���׺�X���8�r�Z�!���8"�&���"��y������
NS6�i���^�Io�$�M-���2J�u'�ݯH|��[P+X��]�yLץR�c^���7�LC��*WB.0��Zg� '#�OV�z;'�-+�9G�B_�|��M&�N���Ȯ��h�ʎ���;��i��6�c��^"W��`�JL_I��S�O�OFw č�ܝx�+�2�"�S����:jB�,�rjB����:_'�n�@���[�6W��|�.��l��?xi���=�Rږ�!�����2U�p���]tE��>X����@G��í�b��m���۔�Y�)� .�a(�@9�M�"�r ���b*c*}/����~X�&s6�jIU�z�8��ki ��b^ �/�wr:���t�c�(bG,E�i@l��?����	*��oњ�w`	�� Y�̰�[H]�v�L�wPD�����neq�l�~�` �`�Zt)�^4M����R^���]�_�mC��)��4��lqg�"Q~����b/�e�r���)�":bJ�~�9���8�"ќY�Z�R�f-z�*���+��X~8QW�1R�ä�C�������ԕ�ܞ�	�0����7RK$����_~	z�a�:2�#a�r�jA7ج5E|V�}j�ѕ�#�A�����j�$��m�$h_=��ϮM@^��F�;�¹���g�z�nϊ�f�l��~>��}3&�妢��~jz�6���ӫ.����mr��5?%�ȓt7����".�������e"9��eՌiK�.�M'.	nSa9�5��h��gf�����	g�$F[��(��B/I��QA�'o:���:�|q�(i�<��J.��=���~=���`���G��
�ɒ�z��'��C��3���rG�&]��uO�}���cW _f1�B�I���W/�X �(��B�dRk�AH@�&2�5J�j/���O؏�}���i��)��|H�t�k8�����?]1�[���AZM$s$\m�J���CsG;�q����ĶdW~�%������
O&E�Z��/���M�����r��Ju��svzi��GiJ��dc�}�z��wYi�XHB����z�� rږ�\A��֠�Z\�W�nocy�=��&v�vS���|�Li���:x~){L\��02B�,42����o����`�M����Ha���'-`_?�Aib<�jh����j6\g[R��N,��jq�UH�ق)��_�㬵�q�l՛'���V9+_1�,�RN�l��ӑ7�i������<$�	d4������[,�a�����(O���0.�}�|S�4ش��h�R%�\�|�����P�P���9�]]!H��i9�fᒇ��Z��u׶�18����ϥ}aE�8�?/�]�,(����O򬴷D]��ċg�M˂�VP���:ߡhdv�=5`�g�p���K;�̃���{�u��zx�.��G� W��a��
��
x_��v��ؒpo�mn$��B�?�LR�u��$�ԗta'��ٶ�}N�F��p��.kw���y����4/3$@��ލ7�Fp0ȼ���c8���1Ȼop�=�e��su(Do�I�w�JW��y��I]W��<���� ���Ր	#�,�"����	��Y����w�Tx�ǂ�Ժ����֞�hlw�ö� d�� s찘������Ӫ�`�K�>9��W�t���6a�0Ko;1X���P�Q|�A�4��_f���y���6=d� ��R0����N�1R�f��Jdg\�r99E��	�b��ͥv�h�/�2͐˟��ߢ�S�t����Mm��#yK�wj��\��:�rO>@��@�k�.�(KF�3�f�=�v�j�N�}7��	�Ž]��XT�����y��,�]�5�j�| ˎ���>���ѹ�L|fS�9�CAe\
_����jRMl�V��r�D����u-�J�@P4 #G7Q�XTX���"]�j�6�C�_���8E���
]�Xf�r�HV��ˑ �r�JRH�,L ѽ?�'�$�_���7)�ʭ�|�6�gN�؂Ǡ�u�
�Yk�Z��菽XGd+_<�|.$�����P���i�x,��At�l����&���)HE��b�@
f���4���c0m4�1��5�q
{��L������/n)�r�gq9��ܢ�5�beKS���޳y0��}Nnq���d�۫��O����
����*�Ԙ����M�\j�hvB.��
@���p�4����S�Y�R��0�t�r��2���j!ҋpgz� �X���I
`��_�Ä6
'�O�L������R��P��zV�xIz�Ƣ����]m�����!�N����Xv]�c�(��%&�-2S���W����u�F�-N�[6,.*ר���,K�.K�!$p3���I��I*�Q��_��7H�#��\��~�� I���w��YQ`d�ZXGu�v:Wn��|���ӱ|k+:Y7�0�'iL뼰�5]�{�:I>{��m<PL��Eǻ�ͣ 44`.�ҕ[X�g���j��׼x8�h�n�?(�'c$hlc�srmn	�u����=��X@|��H�'|�a�~��,�f�} ��n���,�(�-I�Z��^����
,u�l�����6t�#Vo8�p�4|������_�&	���F9&�M�Jih�,<}8@�s>�~}�4 Xې��a	�Γ�Td����:����*p�̋_b�B{H���;wT����k^����!���b�����֓fz`�wv릯���EQ��R|D���88N򀐋:K��;q�!�i����
�uE��6��/��2G�{VZs��LL}��*�)��L\"���#P����6E�2��S�#C��BSW�l�|'� �tmx~�}��&)D LƮ�[�H�V���)��o�1�{"4(���w=��ey	>g��N.�#��7%��n��pU}0s]�e�D���[s*>n�U<L�T�zzs��}�o��%������]X�8�A�T�J�/���X�e2 e��w!��<м�!��{s�>�.m�_5�\���6�Yw�A�{���XR��f"�;�0u��<�L}����E2FUC�����e/~��/��Wog@>������qp#�:��!���P�]��� ��;6�{g�;K�K0Q!�gD�J�IU�6� )�ay=bݯ��(>���f@�����2��?�r���!zeW��_k �Ѻ��G`�Qԧ��!w���f]��˾��)�j�����锂V6K ����p�:tm� ��	90���VS9[�f
[ax[�L�멂�R�Y���PD��T��]��PBxT&��q"�$�1u����s��D%r:����5�<��Q#��千�AFS\$|�Z�(�})A>6����,(v��#k����zP��-:"�������z���%zj�r(+�P�b��������#��P���O�����Zc��[yM)b��-}��7M.�5�|��í�Wa4!���e�C �_%�;>_p;��y�������(f�QHh�.���s6A޴DD��K��[�L4��P@��*���.�=gk�yb�Wk[�a�y�X����g~���~���S����O�֧	��Ō
G���R��d_t�dP�f�pG�n�g1��_�����z��VU�t"b�:�\��8	������<'�1̃������.��&I�����B��*{����akFi���"�t� ̜��-�����Y�֦�l(;d����;��|�}Rc�79��JW�J��S�9Ќy[���l 庖�K"��?|V>��?ř|1�3-������j�N�\ֿu,D�E�8�kN�s��i#ג��ϔc��um���Yyrc��g�g�!M5�kX���w�����d���_%��,��Z��G���$@К�6>u�N{]�dnCn�52]z8�-��Ԫ�(�
���~��N�KO�����F߃��*3���=��t"	��et6��%J��Ľ�R�\5c%��B��9!���VL����<�Уu��<�n�W������"�+���z֌v2~�	�*�w)*h�X���>c:e�Ro'���$��J�u���0�l�u1�¹�^�E���Z>V��Y/��&Њ���'��q^6��i���6��������񥸄V�aF�W8>� �QE-�f���@$�.Z���\G�
�{����t�����X��⟷Q�f�&%��i�aI��n)p�k��}�c�3��/�+mږ�.xƠ����a��dK�t�@��_H���Tq�v�������Z�6.�N�#(�����m#-��(��&�
'�lr2g��ު��g�d��8Kue�\�N�i%n<Ѕ��#LW��B�������X
c�&��� ��h離�ݰ�!m/W��ᦶ*t�|(
:UA�kC�x~�1�UЅ4�O��.R��U��u�g�\YC�|��nԋ	i�<�j�l�ۆ�d+u�~��	,W�Q\bF+��,�R�8�t:!,��݆�X�m�ߵˉ��{$�aԮhV��[���TO	D��&ʓF�R"���lKBo�B�l�c72{�S��a��?�f���P��R�D�T��M?�9U�v�0P�X5����t�;�P���MTe:�_��H~�w>S��3�d,�% M�T��ż�l͕-�$�4�7�o����Ny1#���]�w�ό��X>�4��!-�� ���ԓ�^Te?q�y���.�u��R����(��ؒh0�y��nl��	(F�mv�-
�d�n�}�LL��L�:�P!�}�����wI��m�M��Ε�2�l������m�V� b��(�2
!�Y�̶���6v|}�:��-��GM���5�@H���ͷt:�_�2��E5��6X�ދ:q��G'j�)�5�>E/w<��Sz秊V_����� L	0��E!�� zj�VL���(ee��	D�y�Sy�*՚�:f�
c���b�\z�t'��p�~�H_֛��z���K�[����Rʇ���
����$�s��ySa�͕��Pum�M��vji���K�|�)V�D���[[/�5�G����@�h(��')}��d �N��hH�;����{v�r�)�$
^z�m���>�X��@��~\�Ժ��j�}{!�>�-M5��X#��R��I�ɕ9����+L��}�4��8�+�6�܇�Hp>����}b�U�!�0QA��1qu��Y�������M!d��/����g3�K���F*t�у^�y��7����;a�|���B'N	;���#h��cr���)�&�T���[�N[�c���#��[�A�����1Q�C��[6��)�|�e�6�x� &���N�M�D}{%��Vȏm{+����S�<��Y�N�6�{��X�z|�o��X~�ffm�xN)l}�>e������pi~�������Ou��q�L��M�J�H��6���k˸�[�|0\�����%ZTm��-�0�9��2m)�@��\��q��(w�~
�j|�V�XV�@�W��#�nĊ��<�|jm<%�zᐋ�Z�� ���-��U��N�|�{����H$�sC��đ孌������4���䍶΢�?�m�u���L]�0�4o� �b�#�V�� `��ҋR,�t��	nr��J�F�1Do���	4�2HL ۯ���=�)@�O�O=K^��O�Y���`ET:,�]���21~ޗGV�f���a���V��/�O<��^C�0=�s䱌zud�X>�V�{�/���tj�	S��.る�w�.!�D�%ogJ�����Y�c�vC�	J��L:[[~{*�RED1�'�m�t7��̠���ɏ��mE%YJ����qo�!�o�>m�z�~�ՠuO�Y�C�����'#��.͛NY)��ro00�f�'�s!�*-�o>%��*-+j�~�弆�a�������E�&��/���������pJ���rb����K�����n�)j���R��������'�LF�le��y�x2���ə9���'{Z���צ��xXʇ��u1S��u������{�KJD��X3�<l����u�*���Tʖq�9��,�ӟ����.�u���1���u��n���Ԭ���)kU`?B0U�'�-2�RwN��`��G[��ͱ��!i+�oDи�L�x�թ6'g�]k��ga���B$GG�|�q�Ѡk��v����>\��5�#���8̼7�FTc��I�X��V�S=�.ue��HC�c��������(����*����-�����;x�s�Nb��>�l�.94���~a���@�d��	D�i|�+u3�D�a��蓎g]��z[��G2�Thu�"g]�{�7�p�r'�s��'��1������543�?�W��%�{M��E�q	/�+=wX�&�;�t�%�>�J�ۤ����$�Ó�-�I�P'�6���S��!i��0βꈬ|�m{�/��R�?>F��y�k���ϊ e9"�,ǈ��v=�q��u�4�����5 �YT��ʡ�$��V98���
.$�$��Q 3/��Ѿ��M�c�I����g�bW�V��8ZL.�� N ��	�_:V��]�ŋ]����=�z�t��Z6�aE*�o��o��H}=U��\X]���z'˓Y�31�I0��,xs���$��/K	�yS�?@Y4�`��Z�=�����"!q�g�n��ݽ���DB@�=�.+�b,��a?%�3�y��.�-�^a��@jo_��~A>a?����A){1��y�RK��K!�C�Y�m7���^��_������t��Uk&E�0y��[e���1��$ �ˍM�x'��xp��F����4�&��x��A�~�A�Ĳ]�w�1�Q�%ĕ�o�]C�Ĭ��9�,r�ď�S�o�Rw���|�?��8�'�%�I��>/J�VߨP3���B��P#���E#[���*�뷑�j�;��a������W���S�����@>MV�Cv���/{ֲ����5�"T	Į�.���>���	���H��q�r�Z2нܜp�X_}0'2�e� �,�o!"`)�0V���QJ
{H�of� n��r4jHy�
��{��rQ���W�'�D�Ki�A�Ç�/6�5���#�M���k�Wu`7�7�x,�-xpd-[�?�Y� bh�B����%���2H��@��dkkg	����߳^������K�:��W�[5��G�����~F�G�E׻��^�|_����f��`4�Ld��;kŸCp9�}�$�)��m?s`�V��[����1�����t0@z��ff��vv���ыǜ��6���ѣQ � 1�=J����QZ�K,[�W��݀5�����7�Ƣ��N!�	����[%����r����-�7;~l�"��]�}WxǀA��/�� k��#0����4���{-��g*JV�F�R	��3X�Q4�U��scv=v�'�lD�{�W=�ju�D��D�\|�nd�P}YBh�|�f����C���jA>,ta��	ߤ�r���U�~�N;4%��k�]�� ��N��6R-����aHT6�7��r�`��$�LK�2n���QAw��d{�E�P�,�w���2ց��̍6��]�n��-&��ՊT<:B���B�|"�'��G�ω� E�00�D�[=J�&�@��gAj��cY�U&�s<�k.�4�O!�L��R��")^"���E�<"�U'͓��B�9(��E�|{ɗ�hjJ�ܞ��{�mԦ��2f��+m�D�@D������[*���|~A' �`�6e1�Y�as�Kh�L�'�:\�fx,59'��ׯش�+hݠ����|?c~��xm4��Q��sj�
W{W	PaǱ�vݣ�#c�:<� 3}ϼ!m�ػ��5���
�pO�*�d紞�[J/5�`����������p-ؗ�%gJuRvI�g.�����a��r ���.��n	��PP��� ߷4Z,�r����d�5AVY���`,	f�-�	"��G'\�d�Laނ��a��1�X/Io���So��W,B��;�Aj,) &�\4m��@Ȍ����aW{�/7�X� �Bb�=��7��TA�^#p^�֛rXr?�L]����nA�a��l��1�\�����9y�z�
4���a��� SM1�(V���VX;(p6��@��S!��`��Jv[ȑ�ԛ �
E���N���E8YGH`�%/�s�h��ݑ?�6X/�Gl�|mS��Ny��M!rGE���6nO��03�͍�)���3����DLV�<M�Ƿ���Ӫd���*7�� m*��\�|���,L�H�B ��BE��C�U�I�xst�$�\�?��m<,�6���~���/���*؝�D%���}'��I�g]���A���f��RSL��w�w*�JU�����Z�|N����)���EQ��m7�e�գ�<ëe���3�.����n-�|S���`�F��PٚsD�~�'��a��˶���� �%YQ�bm`�L 24Z�1��`���/r@Ko�+nK���Ĭ�Cs���c���
�z��/�W�S�?A�u ک��$���#ș�AN9�\����G4�efJ�K�j�eKZ�{�Xn����Iz���8��P��ܛ�C�`�Bz�5p ���(����ܮ<g�Q1|�A�,r���I��@O��W���U�>閇V+42"�d�`E���Ѳ�#���rD��Z�rⰹaBX��&|��&�𬵎��nQ,<?'BVϖ����z�G4(�х��l:��:�ψ�E=��{���`�"��ퟮ��qF6�r�dw��<��S	)qO#J��-���x��=.a
m^
߮(O��:@��۴�6R��������ih��U;~�Ƌ�y����09�̐�)#j�#��-a����%	zF�~�/䰍��� 6�֥ϕ[Њ�Pϵ��9`QOL܃\>{�E$�b���z�������E1?j�3Aq�/s�U{k#1�i��{�Wj��V�.�z	� 1���$�n����!Ke��E�ɇ��F�hk%���M����6&�r̘N\�X��_5��M���>1fΒ��_�~�h)����i�/��� �V���]B^Z1�����>�䒀�/�G,�!m���~O��<��M��>�J,�A!�Fmg�Hn�jG�$*���P�� �y�0�9������b��%Q4J�{���l���m�6����z�5p�pnVv1q�+��L�� �$܌S�x��i ����1[NG��hQ���d��a�#�Jw��fc��p�ң9��;�
�������>�  ��	t��{d��}f�T��d@�JGI���1�]l�?.-(6�uN}#? i��`��h������E�騤����~疭�� �[��1��h��������f뒲"s�0�:��ϳ��Lˮ�:���K���/0\�(��0u/�s7��4E��1��qvAQ_�'�1B�M~oώU�C+s��'5�MY�`,-5V�=���a�操Z�,4t@��ޢ�r>����������GЇd��y���u93F�Y�����~%�8CV�}�p�-x��(mW���,��1����&�f� ��:����8n;_I/a�,�c�d?�	#��F����)1��}�L���߀�6{(s������R�]Σ#��c�o����6A�o�m{�S��Yr�R.�0�/�|c�I��+��ie�����V�f��7VAk����!�k�q[��ri���:?���LX�
�yS�,2�F�~6�'7���>�o�.��R䐋���+�\�=���zd������;��ǬR���l����{
�(V�r҉��t���:�3�@�A�:x��#cbU����ݪ�����cu����`96G���:��a�{DT��!^+�������ۣ�X��<*��Wp7���ֲt9� ��n`���B�V�q�b�������p�%"s|�k֜Ra��+@����WC�-��Z�Y:R\K�˝o���
>SF[�gg�p����,^7b�����z�&W���w�,������q��,���Տ>FҢ圾I6+����6�����$2���}.E9��K���{{����S��Ε}�Vo���H���tE��%�=b1��2~x�>I��h��y�W�U�ZTݣ�5��O������7�*ǡ>���~nGS�/M�I�
������;�Q6֏�U��߼Qa1pq�����fDS�_8m��=@�4�!��rXg8��Wt�̛�6:U*�K��8b�F�b��V�*����g5�z!�U�� qb];��Rk�qy�ZS���/;��j ����`�2�<�)F�%c|�j���oV.T	�Je�mH�}Î��,�y�*�/������&�mfāHzh 3����>�fjH=���[bQ L�e�sE�+6�?Q�y"��7�HJ$��*����0,4:-�S�_��@
fz/jɡרVƊԞ ��F5IUz&O?�H���)���m��Z�z�QS1 ��s�79
u�ަ)&��!�>I�
���!�i�^^��߿��^�b|�=�c�s
�Z��E� ]��zC��U/�MZ#��<�y���
��݄?k��ǹ�L�n��eE
�xS3b.������
u�^��Ԇ@�\TMq�7�k���9b�R�r�=�_LBU��=at��D�
H;��yJ�t߻x�<�v֙�Ze_0��پʡ��R�D�c�?wb��Q���ŗ�����>�ƌ�`�-~Ȗ�(��F;cS�zD	�n��$�g�9?��0�9r�P���|-Ge�	+Ht�%a.D���J���q�z^42+��x�5���������&�/�;&���M£U�c�7�R�o]o��oT T���|�� ���C��ۂ	#��ώ�Y<�+[+�G�3�"A��w�:����ꫦ�B���T�z�i�����G[�|����.V��f�N�"�-���6�-Τx�ޞhAm���m���X]��@^�~�d�����rW4W��%1���J�v�$ƅ��;�VfKF�ʄ(ҫ)_���F�fB7�s��6���ۤ��SK�?��'���)2���2z�k3�P2}8��� �\	sb*8,N���\��s��|۳��>���FLE��u+2!��I*V˽�͟IX�%׀Q0Yo�Y���c<>�Oqs��;Kouա(zp�ko�D��pپ�Tc<č�b[�塴:D�V��11̺���d�<����7�k}(>k�n�p܇,�W	�*�K H�oK#ȲЦ����	��r1ᢍ<!D�f����en,E3��d���V�T���*Zyy�n�̦31�?�����3��?Q��@����1I�5���[(�Fz*ٌ�V}��^IxO�c9�����6�̊��ꢍ��"�UY���n9�j�p��˄�\�'2�ݑ	>�F�Qb-H��ŢL;S�&s�Ӭб�j��q%��FI���&_؝)�;����_�bn(��#FF����cb��
Y���x���F��J8�䎱��ˑ�!󰟀R:���j;��?'Ņ;~}��5��P�t�b�G�	R��9��LF����~M"u^�{�z���5cU�9_%��?�K"�Ll�`��
 �Z(��.L��g�)�A��h 71�s'�B>~���G��^��PE�����r�D�G�!�C��l�Bl\H�qIqٯ{4a��H���k�e1c�����<c7�Z�&1Fוj�ʯE)�"��_���@�E����m4���%�0��v�A�:��������腺���I(��>���t� �s��r�o�_�mD]����7��Y؎�u=��b�CB\gمI����7�Wv�\�*�7�X�8g�4(��PnO�����|���r��ϷC�*}ڇ<��Y�hq���hsWO��J�%g��5b�p�i�;SU�a��p��+�:?	��H�:��y��]\"��/��j�#����/?���i�;N!K�yl�ª�)k
��d��c����c4)L�x#^�LH����]�a�Y��|�*z"�n�A2��29G�
��O�>� �U�Q�3�ۗnjr�9h�V#���~@�tE�y�@7t
%ŢQ�:i��~"��j/�A��z��`*.<`t�W���%�x3_�'G/N��7�����z�8z�F^f�-9�	u ���4�������m5b�����R鍦�%�vO���CW"�|E}f�J�����+y�H$	LYTe/3廃ȯ�ta�o�`�������2�],<�!8����/_�L'}oBKߎ#�)�\`t�I1��A�g�[X�(}�ڪ<B��p�lS��nW>���6
��_h�F���sRkzs%+C�JU���n�^����&��V�f��-�9��9Bj�uU�^Erc�6����gr�u��U�Yxk�c��Vj�D��������I��>�'x!�m�
�g�'�l�aGܣ�:�K�є9�pY�i!�qx �{�_��Z����I�phgOl6��@�o��l,�,Ğ�i�*��>�K]�!t�Zݦ���߼� ΐ��R��]�6�ө>�d�F펜'(�I�69�c�B�71ʑs���#�h�g��UM��z��i���A�x����A�G9_���SU^XӪ����C��e̠�,곹/�"���q^#���N:�85	�}�'���y`�*h��O��HC��X>s�`��v'=�6R�n���Л��Xۡ�,C���"����`��-�s�En��=���26�`�Z`|�M�їD��(�%�z�
њ�>[+��E͛9i�"�Tﳾ)3s�Ʌ7U��y�X�jb�3Dv�v�)eୄ�c݁��B�vV/|�D�0c��GCA[a�Q�펷��jT.�d��O��汏��Y��ƹ��ɉS�����'�˴$�o�y�V���,���Z�n����jɛ}Y����&�BlU�p�TB�5���>�����׶�+\���\Qb�n�<jI̬��w��6�X��%E���V�t&Rj�ܯm�A�,T�-Ng�y�8����R��LV.�#��G`�]� �?(���ٚ*)�;�Nc�pi�yx��㩭(���� ���c�z�$1�S{B��1�C����A�
:��<_��^�N���gugux~f��g8��#=���H(�Q�,��Ÿ��ĸ�b?���E�;P�ыG���C_d]�_��SP�X9�Sj�����Wh_i��@�$e� {�z��̓�^k��
W�������<�s&��?���s�ٲ1*M��z�.��S�2bơ!�ĥ$���/I��bLg��4��qʤm�C�f��l��_M�Q8�zwxB���ZK���K`����ǰq1�ԗ������������G�<I�<�ş(���6��kt070�
�@{�9�Yg��Vĳ�Sy�P�ã4�A�ۯ��������!H��K/���~�QSeby�g�_�wP+�q_j�V�kê8�'\�EZ�6���sN�W]��'��0�b�6cf�D\2�U?�8c}��wqL���<���JX���*�-�"��ݼ\��N+�8����B�b`o�_&�s�����yZ¢���i�����g�";:�O�v�'��:`��B
wU���=�)��(��>s^I��`;�}�vݘ�F�wը����WԸ4\=+���2E2Zȕ]��8�^�bU�C���~P���y�X���:��%�_�:	��Y/�V3	�uW�&����\����~x�)ђcm��j�u��ZLD�'u�����;>V���w�]��,}���e6I>zCm�d�"�,RI�P�-������r�<r�<m��B �^���M��t%*O�"v����ٟ��	�=�\��~	N$˯:��i��wə����a@�N��,2��%������~����-\�lI�
�m�j+[{e��p��������5�L`��ۢ�q����K�G�	\�����4;����.����>f�NC����\�eb2К��zA�;g<,"k:��-/��S'w�H�]`y���R��>>}`�3�����h�Mx�[G��}�0ga¾B��.���<�����*�0�̵gW/�)%��\ڴlUǞb�6����T��*6\�+v��ُd���ς(��a�K_d.z�m\�i�FN*%�|&�[1F�ұ��p؀	�:�����c���%��ƪ���_���q�2� !�uԺ��T0pc�UZ˱�c��� �B('�፦\s���hU�S��Lzz�^B��
�Me)�E_��-Y�s��U�n�8H�U��2EG�z���wSL���G�7�<��&~��¤Խ�c�m�9ƙ�hW�Y>�jG���y��N��u~?��?#ސL���v+�EX�=-Obx#�#Gr	�w�й���|�_ �g�xk���U�|� FRUɱ�J���̚��
��w�9,q}r��i������BXnpu��]�}̵�	�����!?��0E�Y6�y��m\��V*��E����"x| y�m�oJ�y���wl��V�6A�u�ը��a8��foꍎ8��7�d�	���
�K�&ժq�^��D�{�oo��jX�xp\;ރ�np;�J�CMe�W��q���Ԥ|���3�%b���࠸~w9���⏉b�������ye'k�z
�֣ɾ���w�L)޳q�2|:��x{I��e9��3^Ig�Ĉ�6��8��l�+��P�.�N��͋ش�+v\�L/M�P�����Y�=:k6}���HnD��\������w6��ž����t �+<�ԜKH���R��qꖌ�W���lh�v�!?�j2%���uKkމ�KA�9X���|R�= ��*C�]'N���5SZ3�$��k�p��--86�|�sv�*E1�Fd�x���%��J`�
��/C$��Rt\_u��R͒��V#�3�(�0AA?N6�ۛkA^�=t�Н�^^�Dƛ��|ܭq�	���c��3��vg���~л��Y�mw�f0�8#A'��#a�7��J��nW�2�_�$,��iS��`�ώeq�1-YdA�]I��{��>�JNV���."��}ΐ����l��9�:1ݟg3 q��[�
4�v`@敪t�!��ˏ��GeD��- 0�&&�V�B�*���MF��8��?�����|�d-(��{/7�=jEm� ��C�����8�5w��n��9�1�a�v�5�h�4	 jS�O��n��;�� ;W�)�S�4#�<�*�y��x����Q��迤�S%\�����Ͽj OM^]0o�K3f�7�СFc��|ޯgr��z?pzhj�]}>���P�Dp��j݈�L��;b^L}��M���Q��f�" �-{��l+���|��]�.��uc2ү�}"�4�k}�<	DS50�7H�o���ܗ�#��`�����%i;�zU^!X�ښ�4:��q(�@dgX���R1�s�y����dHt�*�̮34���Jɿ��m��*m�F;�P���<�,�|\4`�A����Ld�uYN�{A���x���MJ�T���Ʈ X���G%��$���cO��#��'2�VS�|P�~d�� ���S ��Ϫ�7[2��}���L5�;kr�j�`����JiE']��Ii�`l�k�T$1M� 2`��K�z)#|�3�ʼf�^�98AXc_-���̷ͺ4����Ĕ�l��oL-8�U�7��R��V�#���S+Q��A��f{8Kg���7�Id�]�d���W�p~�����^�Ib�}`��%W��˿]��$�먬mڽxb�5�w
,	c��t�n�t9��<؞�I��1�t!.���	��ac#���w㦙I��~�1߄e��\6��)Q��A�~��6c:�Y:�����������ǙD��Rb3_�B�$��K�V|h)_*=Ϟ,V�������4= �)׋ve�@�
��G��kj?R�4S;����XV�Db�тB�� ��Vk��3�z2���{��i\i�G���S�Tm���2�=������턍C&�b	�H��}rՙ��;c�����PǍ�W�Q�߻$z�<��ﰇٝ�����Ă�S�;���iO-߀�H�x��Z�*x��Ԟ�k٥��wf�b:���N�97����CI�A��H�WWيv :�,7'|;F�"���Z+{l�,蜙�����R)�D�Y�oJh�ߥ���JM��T������k��  
�G��Sr���>eE����7���tÁ)�H�i6eI�WC.�%u�i.p;i2wPn��\��RQ��>�����c"�����KE"����\R�6��s�ak���bMq˗B�J����D���u{�?I�Z��F2�$Q��(y��P.Һ�TEnh
}K����QI,�r�ėw�d�kg7��Le�*;���܋,�L�g��Y��7'ִ�<��5�9B9D$%?7�l��;B_'$�ӆ�t����!g_����tU�)O`a�,|�
�no�y�ӓ'��x�L��|ۥ7��ݒi�h�g�=-���"�!��G�ݥz` �a���81h�$I���*�|�h�&����蒂hg��g�?/D���4 ���;��ٌ�\����bFR	n�����L&�b�(t�
+dqgݨ��h���10��=7\i��P-VqC�aQ��.�[��A0/���jv���?��`�B�����4��ùO��]�pQ��ސֺ�[�'�m��-��йRĺ��d톿�Kg/݀_L�E�Ԩ]s	�#Q��ѭHD#���ߚ҈���R��'�L�t�S��/��iD�=�&��4|?�\�2jQ����_��*�ĩ���T4��2����o�J���,vZ����"�W��ZRDR��1gU�UXܲh�='O�r��/�ɲCh��Elɝ@�{�}-�e�t;�l����0�[����˙O2F�e�=�
�C;�puN��Lg'���
Ea���1�1��<A�KD:�-Bţ�E����:�D�����_��h��j|En��|����={QN��l�����+���w��:T��}�-о8B���4�����&��[��z��@>5�H^ X��Lg<~{6����Uǥ4��b�8�U�,E��d�Z���xW2Q�WT�x��f�A�&�����H�s��	$�ƏQzw5c�Ep%2ϒ�`�T�@�L��03
��Kv���;�qm�͙m��<uK�B?�K���"U��`B
����c@Z܆2�����x&~(8��r��ໆ�A')6i.���ǐ�S�ݥ(]�"�����%�َ+�h$�ј���ouk�}h��0�VwW ����2$@ �U"��<�|���%Y5P)��8�	i�%�|�!�Nx�F��5�rf�ɪO�ml�I�?�-���/K�X?�����~5	���t����3�=�L�eVc�,f�{�˽Y*�A^y�Ե~�@�����_��4�Ȫ{m���Ѥj��Y�3y3�rUѝ;Pۇ�lHMu�=�M�WA-Q�S�τ��l'����?iˊ�A��l�Q���»;a�hs'Ɉ���ˬ_?�T3�l�5䯋�m	�qn�iX���%9�z}�SpJ-7q3_�Y�����TL�, U4`h-��{O!J��O����=O��U�̋��1o�\K:�I��	��'�uH(3
'��0O�~B��k�.IF[Ѱ�]���c�0�Vr�a RSݏC#]��G:�K7U�ze��Z���	z�#�{����L����!���!.�b^������Kf@y�J�#��'�k�}���c���"Mq�/�T�;�Y�s���� �.�yף&wcu>,9�	�?�d.;}E�k|F��Tz�T#�od5��.�.�0��[\���U�:H�g5�5QK�����N�V��H�������W��؄Շ�\0��O�{-��!�"�f�.+�i�V�,�	��0���Ha^]���Cd�G�/��f�Xu+H���~�CҸBp��d*2�:m��3���{���+ʒ��o �S�X��R��N1��p��|�����
;Br^�6�J���SG�lx�!4��stc�G|c1�y�p1Gy$4	� � \���h�B���Ȳ�#��Qgd60~F[�a����"��h��B����E���$�������z�x��@9��<�F+���,�B�[�� �ŚG���?��$Ѽ\�W�8n�h��&�C!/��̐�����	�[�'����WT��u<�H<��� 7�3>�-q9�\r`���j�(�F�GW'��������%������:��@��W�)Ed[\��Rd�Z���or���# EB	��Sΰ���ŷ�=���U:z�^�� �1�?��%c1 ��߲U����$�[{K4��Rn��EHb|��e��]��JrM�-���C�ДI+>����5;�s�r����2o�z8�"��lP0�ܬ���:���������\��@(C}r���P�	�]$�f�M�g�gB��=dp1;$� %s��;��[��P�pkO×�i%�6��%@,�ؐ���ۜyp�A��hXT��Iy?�{?��}(�Y���~"�if��2K��झg���U�J5�N��� 
qf#�6�L?���	e���:�Q~��K<���IQ�sZ��u\�}(֡\o�f�����"`x4e�EP�^�����4�q��*�_	���\�3�-. �AͲ��kUe!(�CL�|{���p|���H�5�.��2L9� �����CO!�� mβj�F�P�Ӿ7����!�H�9rW�\,R�yT��-�/T�	KO��ۯ�#e��B�J(2�G��n3�Å&)���'WX�ډe�M��s�aԙ���檤6tQYʏ޴ ���G�MŒ�w��0�[�&��| ")c�p�!6?�^���:K�W������=Ā��Rdb�Z&�]�vEb�V�_���2�f���Y)�i��'u�o�`��B[���lJr�μ%�z��X�� I�ϖ��FqTC�9��~���9�Cwj�h@��|�1���4�n�S��}�#���:�T��9������QF��u���G����>m���wL�x4����EN�4��Q�=L�����ƿ���̧;d  �Q@���w���H������&`#��h�Jk�L�~�x���{��"���
5����Ks�s�f^O���LEbC�y�ƣ[��l��*�_��l��@�A�_ �'�8�F!�s_1�Չ��?Y���=��Hl��+�����pZ�..���P�ߋ���wmF����l遰XQ`�1i�7}c	�E���!��0c�C��aܾ:��P��5&��9!�I�c,@���V	#�n�*(�㈖�?��=g.��)'�|�O��[���s�����pgeW)�'��n��6�#I� ����R��G�:�\���O �ޛ@/�R߁��s�/~5d1���-cy��ʈ �ҾU�-�XE�q�X�����PH�B
<6�L/�U/=3ep�%A6	���?���՘���X�6H/�~�����s�Pf(/f���C~����<٬���V��s[L�$U!ۮ֥�a*���ך��0��o��`��6�sO�v���j���׊(T�� w�'.�g�CZ�%��?I��P1ef� t\���$.<=;�>w7Ў�7],x��,D��&Y;S�;4c��P�4�CdP��-�_��D�G�p0Z�*R߰W�9T���4�xj�9����u�ak���<�e�pE-�[d��&m����T�����D�]��=���P���C�&�[�\��heJ�#mz'X�����8���<?���B�lk)>�?jE�?l2����Y~Ј:O$L*@է���u���a� �#Q9�/v�!ۮ_�����ӭWts`�E�	`n�J*�/��Y}t̷o���(h��V}���5���9��l���� ʅY�zҙ��d�w#���&=ZN��UQC1�-�9z� e$����}a	� �r��[`T�Ca����������RR	��kGkK��Ry|�a�A���a�`�-Y���1��rp�~*g�����>�d�+�\����:�����gA��8�VVOI��cQ�Nے��sñ[K�Ȼ g �e�E�����Uj5ξPO��Aw�ML[�"�=
rں0���N
�ɘ�%���7WA����Y�5��]C�ͫ��:��s 52I
��|M
������%���p�����8���	���2�5�, �3����
��*kӬ��%	(�:�_���v��4%��e,�-��)��{�����>��5��4~�]^a�&�*��/RE���z��,E�K'"�=���1I���%ܮ;�4!+{,~��6PŐq�s։?ֱf��i��5�;��Q�?Jհ�X"]Σ;�Jc�`��tg�����O�N� ���iK(@��gtM9+�._6.��5-sR�-Ŵ0���Q�ץ�q�����߼�j4��$�T��c7��@��A(8��W��1���T'+;� 2
x&:�2"���iHI�Z�r�鑤7N˝2\dʪ�	鷐;u���H�G�+
�Zd�4��^�ܳ`�E�5oa{M��3ZK�����L=���ՈfЅ��5�����RT�� ֦s]�<t��F�A�V��8�^��6�̀}B?�ʂ��(:��RO��.SŒ�j4�<��.�=)I|~�\�A���z�Q�F~�Èo�[ h[��^��%��N��+��\�!Io(~��Im����2ED�;]Ĩ��9���lv�I�#���NJ��*�:�^�r#�37<-Qh)����~�+��4�>�l��
_[L!�Q[���qq 9�7���3.���Z��F,Z��Y*�15�Ȋ^�xP1o.Fp�cN���'t ���±��0��!��OO��۳j��o-s��Y�����por^����ԅ�2��G�ńw�3;�?jH����)��ނ�����:�e&�0t������[�����F���ǓƢu�b�nń/�&$յ�`Iai��ys!�cI�t��drc-,i1R��U�Ap�3?�:��/�_��W�j�3,�?f�	/mM�����L�5㋾�Eh�;�����V��ѸQ�����.G]1�����{4���VA4fX��b����/��1X\n��Χ���i {w��<@sT�X��FE<��"Ma�*�%b B���P����ùfq�+6T3*�"�������7��F%�>�Y3Х�<�����N���C�2ѷ4E8�,2桒���D��t�4�@�+�L*��wI��������\iI0�Ss��9�`�ʇ���@<j}
���73J������]��~{���%X�_$���4������a�7ۑ�	��M��8�����љ��r�6���3|���CS3�D��cMG
�o�S�\�jp��^�Ϣ��; }�H���B�'F`S�����#��nA@�v �W��<e��ƈYü���(
c��,]No��'LO�^�� ��7�rt�v��atX�DI�΍�t��7�/�j|�>&�<��,!��ulu�UB� 
���	q��c2JI���,������0��`�4;�Y9��8=6��c>�1���R`�1�̯��Jݒ�:��`���cϝ��Z�7l7o72Bh��JS���5S	˯E�I��U��6
Y�� />�js�~�PbvF�c��x���j��p7@��0sϑ��^���qx��U�{R-��`��
9ED��\���8j��	m!�x�n��W�໋����9��$u{���7~�
���E���������z�X���aZpy�~kö#KfN��:��x5j.�^R�k+0��4u���$��2��}����h�#�(����#���XL.}�h��Z�h2��e��\��o��e�|��w5���Z�Ş���XD�۩����s���׃Tq&�^�ՎyW���Yp�V{S����c�>v��.��`���o׵���u�F[�;x���(�_*���mv��ܚm�6�I9[�[Q쨉��#���Z<�I�?U,�T���9�ٝ��p���Q�G<!^��
������`�:}�G��O&F?�Tfg�ƫ��I�y��V��C�����9|�%�V�}��wgo'(��}��;����Rf;�- ]�bcڬ��)�2a\ߏe曞_���ˊ�~�JB�M7H� �F�V���!��uP�9���;���{B"?�Wl�� ��2+86���Ub:cB@��Re�cl�����E��'0�� ���v�D �{���U�N_�G��σ�csK����f�r���,S�70���NA�X`��C���:F	U鼸>�_r��c����]�#Ž-�\��D��{\��ڏ���#��NV�/�9��k���d�+�R�O�Q�4��H�X���0TP����Ɛk~MYH#��s���Q�]���ǵ��r���ؑ|i���RB�l�i����Et!;�!�/Ǵ*�����-������.��F��}��<E&
�
��"G�w\w��3_�)_�#�G�>:6T|U(��[��(��f�!#0�	TK~̱�%�B�pb�r���v��Fq�l7�㢐^�%�Ck�\�5�m+�Y�e��|ձ=�~���P�|��An��d	��5�������eS|L\��gyi�D��1"�#�#JT�c�*�:Fg���1���̴�^�q�D�(j��f��
�2y*:HH[O�g5�h��]�V_*"]R�d�dѳ�J\R4�<�Q�`���;V�Z�L�\�o�躦 �U��-��*�p7N?��&��Z>�a�q�Qe��ph�c�4L�_� ��0��s[(��Y��r+d=�-�C~�0�a��{bf��[����1�!<�{�><����RZh���:�ȏ�g(3ȱG�C�PH�O_:}7���
��(����\P�#�w�2c�c���DJ>��\�r-s���P�2?48I�Vnw<ZQ��^��{i�Z��#ҡB�O[R^�v��s��8�@i)=��c���=6�z-�S�Jd�f�.�l������o�"ZN�C
���39�U8ok���(S�b�C��x�.������>�pt�o�v>
���M����P���/�*
�7���n[��H}�i�,�`�R�녧����F'$@��Ԧ%���:	L�X\>W��,�cJ�~)�{k9#[�#�m,�Z�3<�N�k{3j���Fl�6�ajMT���8���z��I�s�x�8��.��gL���.�Y��t@�'��9͖)�_ɟ�2{�#,]ύざ��ݜ�'	Y�;��E|�М�aO�����=�&iM�:�+Bʎy�l#h�oq��`��4�D
�J��pg����ι�4Q���X�u��ïΨ����A�CR�๜�9𥷯�CM����o2�89�����P��%Q�&��%�z����|>E�M������,zÃ�d��LyG��is[�CQy��t;e��%�N�VC�DSj�u
�f���^h�"D������;$�wQ��-����7s�JL�<��-��e�lF��V�D=W�CeaO����Sft���.'��;!C�@�߮xJ�.�'r1j�c��1d@9��*12�h4��2]U���ɑ��XrAy��H��D� ��2��4����x03������&(�*���*h��|M�|'�� 6�f���Qr#����� ��9��R�ڄS��-Ff��Spة��B�����1[d� W��9>����1���p;�鯗���c_�p�S���X5}i}?�����7I�������{�l�Cſv�d�]8R��:i�Q!z�f����$�ك�Jv�7�{�A�Z�Kh�rA8]W����=��BB��):��8d�9�����Bj����R��P�� �����|��k��7"��j�U��[p�Q=  �Z��ܤ�����`P��W�+?��[��˛L��� �������t���*B�0�|:���I��@�S��G_��;WDR��� }]���^�5�U�y?Z�iutbd?�E�ŇMx��o������C����ߠ�1o)�4����{N��)8o�)'H����rYDy4��:i�����'Һ^~��+о��q�"*�z�~��Po���\N�yjb�b�B����(-�����V*� �|��6K�F��d��ь|���S�o���}E8������߭bVB�,�休q���6�?��Yh�<�-�v]��T�z�Xpm�QJx}�3�WV�<
�w=S���Uy �4A���iw4�o{y/aU�=?%��%*i�x	��]1{"35���,=�ҁ���9��~|:���T��>"�������- s��'F;�|Z����9`�[Dw,^~t&fD��1x�a�|e��A�.�1�"� ��Kf'�[K�t�r�r��^�Փ��Rv�Ƕ.�=��.:�p��P�-x�o;���-��v�g��W����� ���#�X,��ЦXs��f�~��(ưn�����6(���}.!g�3�B���Rw�*k���ҝ^�a�n�F��4���I�$Q�F��� ��k
2-ji��������6����8q�. �"c�q�ƣ���+��٘OrR��N� G-D�-'���L�혐��q���K�oZ�}O�j�p!fd�bRL�'J��0wgrGݘ?��~Y�v5�0?��֎�N���Έ���q�\��U�D�@�C6F�����zQ=���]����{b<��4=�J+a��9�Saԗ�KU��s��V	&XD/cG��)z;��k��[��V���7�t �6��\>gd
'^V�pm��g{����l>/^h���e2�@Ս?���L�����`�2�Cf�;+�����&��CG?q���]��G��*�a��Ԥ$�l�)�M���\�u��h��i�ں��l�yC�P@7k�ɄЪ�+�UwF��=���Ru'��C�XWK8�jӍQ��v ��Dm~qA�(�*Ƃ1�7�-����ߤ���`ux��.X��LH/����g#D�;]��G�IH}Y7�*θ�E���~�\��������r�=J��%`�����H�R�ҧjk�.JT��[;�P�
Ev�����Fͼfjӊ�a�A��=���܉��r͟d9���u�'�t�O�|�T�U�h�Քc���6M�3׼�mݯp8�3��(�|����u,q��%N���F�){mBI9j�lO���Xr�ڢ*ql{!� ��<�I�߶���e6�����!��Ͷ����<�o���̒|��o�JY�a�akF�6G4��+�]����	jR�6$�20/aͰ0���c��D߅H0y|)�3�gE\HĞ���Єv��.�Ҧ]>O�e���E�4�� �sT16*��
���M	lb�x�>{~�E���w}��IZ
�}�k͊\��/�xDu�ױP׭�1U�9M�e����J��Q,!F��=�(H��&Ar��;�A�b�@4�ER�t�ˤ��t�^�~E���9���I��n��b}��h�}'���i��d��'��t�,;�Ȟ�P����Ѐ�8�WU��'&yv#�%���W��VUhÒZ���
-2#T�յ���1��r�M1�E�)yL��Jq"A��i�F��} l�א���g�q9L3l�� ��|j�an��*`�m~�B�L�;Њ��'�YY#�j���>�-������qv�uy7�YӺ�P�Q�u��A'P��#X�\�b���*�޳�Tx�$�gjZWq���,�~%��]W)�e��7S�X0w+�>Cӵ��p��3Q	���:e6;S)�XzE7�#�T>z�׆Ӌ3��\�$c���5d[�zq<�s���2��38��L̩�V��{�����yPPd"����Qu63d�[�XKeZ�$�Y����	���D�<Y�r���}���$h΀ze&���
��t?�n�K�L��^;x�8q:U:�����&�Kk�!�.F�up3��3W��b�U%6�s�U��I�*[5�H���� 9N�}pW��;w�$Wl_�|���G^���p7�FkUn�4�)S �ՠ��pf��=����AP����&ؘ�_�ë�%�E�0��nD)^{�u��^�D�z�2y��%L2)�K��]D���]�A��
�4�L�i+�tE�y�!&������H�ww�o�/j��kR���pu��PS� ���^o��i��~ŊD^<�X�!|��?�k%����8��i�����i6B,�����T"��7�me�;Qn��&��R�����2��� �.���g�o�;��"һlIn������g�3�a�_2p2|B�:���y,Ӏ����͸�����p�I!tD�L1��E�>l$���FXW<jc<)2���Sl׿�¸ Vv�N�?��6GK�_���Kԧ�s������7����aQ�Y',>�U�]ߌ\�@}$�P�0����f����?tՒ�I!���$�q2��]ą�!w1�����2��L�E�+�|c\ʄ��~I�w��1>Β����E�E6go�DI����)�3���я/��(s/Vk�МgA�&7gR�;����s �	Z��f���nL�Ơk/�J�_p�K��D,qp�^�'��@�����h")�1b�F��԰�_�п2�{5�+�z4"���{���&�W�$��ǩ�@��"m��6��'{/��f���)�����W�C_z��s��jt��yB@��r�d+3�`�p�2�b���J{'m��[x�qm�Ϫ3���ܗm[m��y>��=x���.���`0�^# �HAyKyfj�Z�q.�6ݡ^|��\.B�V�{u���Ny�w�
`n!m���6��D��@ȫq	����F~�bu����%~8ᡴ����	��Y�����QVp�B6�*���x[6�T&���z�B͗g��M�Uu��
���/I�$H��J4�m�&s�0
x>��I�=/;�;f�U�%�DYp���{�B���N0��VRC�����L�L�C���[���_���*&����$~AHv����z���	�I�����?�ƫ㄂�UY�b��f
x�o��c��}{ڠ7^�C����"�5U�r"�ʕї�ˣF��ب2U&�8��Ց�
��F=]�*n�9�&��r�R!�����N���z̛���Z��ٶ�6C!Ʀf;��W�V�g7M�zf�1"��Dl��ԝ�:G�D������qv���8��:�,�����:��H<��Sｆ�?���=�Vk!tw:@h��<�Y}e��/-C� 0��ژP�(����ۥ;*P�rB)�L=l�Ʒdd���G��|���d�Nź�3�X�+�/�jŖm$plf��v85x�7^�0�ȯuwSveG���Ro�>�̀�� ��P�V�8�F`�VkY९!�ET�׌<R^q�
c&~���_��	�]=�I��(��K�B�Q�����*�-3�
}ost/e��X�%2�I4��qz誨�o��pR0�1�V��]�~Km��FA��&C�mQّ���}S>"��
�X.�$}�����V�+2*O�i�48,�	���'�nodädr�-g|S�er9Z8���!c4/���чGP����ln���/��s: :��4���EH)N����l�F�QǊ��˂H�U
�}%�)�>�o@��	��m�3QGJn�x���7}q����#�/W2��b�/�ܯ�1,����iT'ONy�>J0E�~���oa{ce���w���@�ʭ��-����n��j��P�G���C���&ٶ#�"%;�3�����v�v��<�\/̎��օx<
dǽ'�̴��"���SYC����-L��!%tśt� fʏS���yz��L/s�:у'����B�H՛�ξ哠��ڊ�:�O+lV����n���?��2�xR�31Ҷ�2-�N���_�̖Ն����]�B@���t��).�����#]��~��CF���,�H�5Nn�9B�Փ��@U�;��J�̜���Ս	�4dB)��̄��B*)�z���,�)���!W�r��5q��R?�����ap H����_R��7#�-�z��}�D �B&0fa2��BH�
����%�>ZQ�B����I{�ʸ���W}$탘CSX �F4������H3�$'f�_@�wl�6��]�s�2q����#f?d2�ܘe�Cb#�A	�_��\ڋ�_�>15��1�r��%�1�UU]=���?2��R�~Pk$���C4:A����_�m�\�#���s��m��#`��/z��{ٸ��S�WY
7w�P4�ϙ����&�rK�8�[���Y�#�%cҿ�V����7���A-dj��`=�����E�^M��D;��ZY|,n��B��5rރ�ww�*~�2�	95D��������$+��8����W� ��v�9��U�߇/$W�Vw����{����Ԣ�4,��	b��qz�[sI�	�~�~���2��gב����MP��oZM�gi�vIV!:턢lf��;��r���X��o�?�����Ag���A�R7�LC��V ��X�6��^�ڻa�S�V��
%>߾�zG���"�o�B����> �����F���8�l���N�5��*ʬm���c:K��mL��sp5�Ah���m��iI(w.J�>�1�W������F��W��ۿt����3����߉;O�WD%���c��O�R<x�U�78L���>����q�08)=�<�YĻ/<,�zX1.J��?_aFaf�c-*�W�JJ��+6��N�p�3IMKm���G؁�獢^Ff*g�'	œ&|*�ͱъ	Z�
�
��F��uBq��\�'�y�/�G�{4ΗeXm�\l}nh��}�k��U��A�bS��]��������M����w��w2zƖ,�,�YQ�kM\<`�h�k�<v���b泶5) ;t	,V�"�qP(�������`L
Rr�p_��V���P���w�/�<ɷ�<���9������^�VT0冞���E�7�QSf��;*K����,A5���Ej�K��S�&��ǍUs�����'��z�M$�(�:�N�Z�3[��?T��~�Ē��ݘ�y;	���!��7�§
>�ڢ����P���,?g޳�<�{�T1�0�>@���|v�i���Q�:�'ܱ��?��l"��v)M��P�,&�Lo�;C%�.L�6j�����ۡ��`���N+���־jI�*2��L������t:�͎>m�vD����&C#��z���u��3f��iC���^pi<as��G�X��o�O�K<�%�������Rwfb
j��.���x�a>�����g���Z��G|����7r[�7g�H�un�^�-�wi��ַ�vޕ@K�9ټ�SԌ��x�Q��ݨ�ߵ�t��r)2��R�,�r�=!�p��!����zZ"ƪ�bP�ϗ�����N�F���ݫ�|SE��Cm�G�X���*��vC�(�)�U����u6��w*I�VW�����h�Y�za�3k�+�<p��t��ǀ
|�9D�PY�?�!8�9"����%��F��#uNT٭�B���Œ9sQf��WC?
�V�'�Ĳg��-7�M.���\H��6��������+���dYa�L�r9�!���Z����/V<I
D�U^����oU_�q�4�������XŜ�������r4��q;�i�`,������TR����O��5J,P����D�ϥƙ�����!?`��<��l�nĴ���W�o���f]p���JS�����z��)��F"S~����� 38�E�C?�J"ߐKO�0!��?��͜����D �c�0�\|
K��$9�?����f�P���h1��?	y�?k���t{YGx���fw$�6_�ID���Z�"� ���W���Uyt����
�|����w��GpzG9V]�'�_u�y�(fU�5嵑.���U�
�~�붛},{:릵�˩�BM��kWs^{P�,h��D�+Y�C��!��mb�B��|���#�œ��x�*�Xn����$�ɉ��5���lU�5�g�p�u�!ҋ�4����m�jJu�<�����V<��y�lL��e�C5(�
"�Ԍ\R�O=�1��"�$��ĜM�=&�F���]n��q��Z�Nr�J�O�M���%N�XA�x��������'JwB�l(��!��#՛F<j�t���(�(gTѴ9سug&+P�)�q���Q�b6۞W�4i�ge��ʐ��tx�7����e�ҹ��`Ik�F%����N�������g���`�Vp$zE[r�Pe^��>k�������p-�g��X5�q1!�w4sܝ�e�����({@�gmD.�(��/�8?"��S�l�6x�},{v�����-X@	�ZOϦ�
��ߟ>n3!���r��`�gpX-������
16��0w݉_�o��M���#�u�R���N�YVh�w�9s���Q�@P�X�;a�O��9N�^��g�Bڠ����h=��)x�7j+Gk��c
�Yzj�%�p����ʏer�p8��,yj�`�-���5��j7V�	E�����
���'�7G�V	=+0~k#i=i <~����Y��?(fN�����t����p�� �����'@�>�&��5�l���=3��Ф,M=�h��9u?���O}��$ur����M�L4����2
��͙�Gh�=[)����r�C�C���Qx�<��ޚ�`��i���D	�y!�.�<{S�FK�~AWO@���Ie�{;&��ws]��6��oG��'��C���M�T�ptH�n�B�nL����8�@�
�$6G��*ħ�c��'n�!*1���0�T��UKZЉ!�k�\eI7�S��?�6���JG��M��jO�Ck3:Z+("�URGhUx��-���M&J�|��f ��d�q�fBQ�4����XϿ�p&n�]"������d�Y�� 6���/B�`so� �!cj�kh��%o���9k�����ݖ���sd�C���<;���)�>�?���iy���n��	�.�17Ȥ��`RrYs���X8A6$�E4;7���V�Zp��A=0����s�4D�˪$��s��4ah ��vK�U�)�1 rG�0E�N�=G/
V�����5�TG�����,zC�y���.�J}�,�
E��J�/I�Ƒ�87R)}��W�fFܑRd��
��\L���F0L<嗜q�_v�x����.����46�s� #�1]���/��?[�7����]����e`�ô���t��
�%��e�Ġ}�4�]5��@Y_.۰1o>�=��-����
��j��ֳ���<�u^P����M0�ღt�a��PJ��s�e����OH��D�@A������i��û��r��(���w  2 �a�YT[rv�hLf=-�!��G�R�o��+��d���e��`���X��TNmd��>2�ϞT��i��~}Fdz�h�'E�k�7���P8�z�	��pw1kǍQ��ak�y�;K��{[$���J\���8�;9��R;}�pt�^��.��<����>�����S3���}��1���<������W?T��e����曺K5��b#���L��>�nH�h���7�$�mM2�!�k�a�rA@Vv#��O�_�tYI׻iO��n�(2P"���86��ձ]��s��t���UbD��Ӹ����\	�Wh���k�{1���֦�ݲb��ߗo_��({إ�������HU-��\C+�i!���FhM!c4�=�/��$�{�u�d�A4�}[��������U6=�����ec�U8��C]A�L�UR��A�H��=�yA��z�yS&���w�=���k˼-�)��r��\P� �^RL�u�������i����2���gn���?�(5�J��
�G���?렕kg���+�S�kp[`Pd�ӆzC��:�X� l����)������]�B�y:�n����Y�Hjƈ2)Q�J���~��{�1T�
���7|1ܧ��a��N�u8�-�rb�`Ze�VQ� DW<I_�XK���g�;��b����h�
=(��3�qu��
A�n�"E-�{j�LF�--�GR� �e�Q�_�����!���3�Y�^��q_��d�B���C�;�\�[C�X3�T#x�Qqw<�*[�D�}������t����Jr���A��%�a���&��c+�1H�M9l<�ʡ���϶>^�~�P���}r�� ���%Y��U�׉�@��`(b�p�C����"�����(�����T�����n� ��u�vD�Jpm���Ns��]*K:�[B:�����	��j�n�$뛔�e�CP�b�%JB'Q[��w����ͫ�_�'P��\�NfKtjCd�̈́&ˣ�ʟ��~��Tp�}�(E�\R�p�Z���!��
�P=/C|ݹ�xei�QT#Ҁtm�O��H�`*�W�s`��Ih����?�̖�I��K����L��^	�H���{��]�P����?��ZA �h'S=Ńm�iG�PQkE��������CXA+�nǓh�D:p�v��.����n�G�c���������6�pП��Yt��ȒNʤ��!���W��}>�N�P�����sr����Y�T;��{Xe-8l�;����
� 	G�o!j�)\a^&F�,%�;W���tZ�f��t3R�3��9�k����l��w���Z��uD]��P�ߴ� <����B�dt�pd7�hm:���t�d�w�&�>RVw��ߋ��Γ?��O�Ǩ�,mU�	�7�\�L�U��ԭIA-��NF]f"=�N�Ƶ��k����n�'X������&���B�X��ڹ�;�>wH������d�
c?�Ф�D�!��/�����I�ڇ��X��U��af�W��17|Tdj�>A��ohZ�:n���RI}BRpת�@(q3�����O7��e�9�X~����� �$XM:�+�/�HfP��x��2|��b}B�Q< }��"J���������������|�T��9 ��c��!S�>��-��=LH��!cЎ���bj?�NO�Q4�:۵��J�����) �5�yl �Bj'		yC�c���ҕ[Tt��B�B>e&ڢJ޻ 7>�J�����?`۠)��
ӭc���%�^9upz�;n��������.�(�-򗻜��Z�a=�c����q�Ex��x��S��$1YΕ:l������Br!�)�=�����Km[�+C4Rw �i�En�[u�{D$7�'��'����Ao�{���zKF:R��k��Yn��G
ْ��@���w�T�s����5%��*����3
��f�UZg�Z�c$�g�w�S���D�)�8��"����?���᠎)�0+(�5	�%ߋ���+����Ʊe�ׂ�W�i��K���ƮgQ� f�A��('�jԌ�ZHm⇧j��
�U����o�Y�I,��":��p4��%�p��;��ϳk��;�4�i^�^x;�:#%Վ��ĄZ5p�M�����e��*���_W93��O���}�E�T�n�/x����o?���RZ5PE�������W��f�/!��l]�Kn���#E��|r�`�"K"�ܡMR�i9���⊠s ��`i$I:�Cwf����]l�7�����pËEG'Ek �n������K�:�}Ʉ����h3&�YL�5S4�Ŋ���
/nd��Ѿ�y:�N�3��ze*\q�����o�k�dm5��D��i[�2�#
�j���q�I�T}�j���h$.�ٕޥ��uzA�מ����=���8c�l]!p$Y/Gi�**%t�)�oJ�in0o�V����q���;a���&�(�č�����'3D�fE:!l,*ʜ�C��[�/���M�MC?l��d�xH�Nhʉ���"9���B�Ї	���͔$a�))TS˫n3��;uZoR��U4�����ȋ�#��#�l�8�oВ-83��g�ő���4T��<��!k�ȏ6�����;�\���8_���wrοݳԃ�r�_���G#�t�#*j�Z��pɯ�e�>�T	���Qİ��/��!���d��~��������aKٔ���a?d���5����%ٳ�� �XK�6�֑ o	�&��0��K�d��������D;����Г�]+<�6]�!��΂F�sH�1G�E�H��f���/8�^,��c���XS�{��4�3��ƫ���T�-*�������Z��Z1��i���#{�h��ç�Env\��kG�P����T!���������3\���i*
3��a���䲫�Ȇ�J����+�0cn��NO���k&|��b#d8Z xV�d^|�7O5����w��!���ME��u�A���ܛ�_��;.��w�	��<ޥy'��S�)-Z�P$�.�-�:�A�myZ$�6E��S&w�϶$t.YG���5m��w��	�Euqt�5���mp�F�E�� �}q?���ҵx.���¼��{�M�:
�)��O�nuM1O�L�������T��2��:A�O ɢ�q"ȱ��0�I��g!���7l��a�r����6y�����Z!�u(����&$�471��/�vk?�NїY���p�{P��2�k�G�:��9/�|:��� ^T��	��M�R�R���R:��
c�O��!#�����Dg��V�cY�|P*^��Z�`��"y���k��ֹކ��H�x-ڞ���mV��:i���LL(��ßv���[���M6� ��)��ݏ-��p4��h�Zu�
�	7��M>�X��d@��?E
�@j`��VP����ԁ#��i������:7�c���G��bvw�6�@��2L���lG��A�_/=uD��4v�4'�G왢w��F�R������&X��a���;r�{l��~=\Jka��^��~/\�i4כl���P�����t���VM#��/���aJ��w�\W�J�Mt��?������;KȐ����?�^������F�����I����?q�:�^Q�����������b��G�]D��N��~��^�r���C)�Cض3lR���#UH�P��	�ު����%���q�ɀ|�$J!�}أ�EU�Y`�~�|֟�ǄRŁM�9�@Bĸ���Nc�)-�����p�<_G�l����_��憆��BDYT���ZZ�յ��W��)���YȺ]�t���.̨�<⚀��y��7��Vʬ#\����$��2ӿ�HP�Wm��_à�-8�ٵ̸�rc��p������a�Q�b� H+�0�x%�����ovt�_<I=��l��Q������X�Ǩ� ��y��]�h�{@����Gt\}i�FDA�6����/ȹ��g���(���$�����<!9�͑�tݮ|Y��
Z��~d۾򽒜&/�ү/0d�v�P�o����@L�"|���w�7+���C��_C{
�Aj](���B`�9�u�;8Z�hY��w�����e�
����d8��f},֚+r�|��O):j~�0�=����wD����I8z�L�h����)���e�5�=��o�]��������a��h7� Jڂc���QZ�ω�6�/nzg_H�:2^#� ���H�+�QA�P=w�0�UC�_D
l�����+�3�Ø���f�9�e`��_<p��}�v#�(��1��Yҫ�,QQrz�J�{�Z����A�`l�=d��kʑ�+N����V�}D���1!���}�Lm����Ᏺ����^��c	����WQr��	݀9D<����{K&n���}��6����n���lj��Iቐ�Ei��0g���׭�-�P��H����. J��N�q�b8^a�����|�F�An���[�n4Zk}1�D C'B�I�Fm�u-j����"^�d2u�db8`����"�摹�=i�tr^xWű�:�
q:�7�&��r�i��e!u	fS�LTs��\1��(d%�	�:�*tK_�)�|=�M�P\��k1������"��Yh��q2��ڵ��� ��g�F1����à���ֈ�]=�eq3�MwT���`�u���P/������^ѣ�O���R *ʄ����9�*Cu���r��d��M}�C�d��\j�?��T�ݫ������0 ��#�\ǢZ��:��^ve��v%J}�(t�#��W��}�9�v?�c�Ȼ&���OI�87F6;�����;C���'�r�JG�zh�z:+�iLA@@>�J(3��  J���Js��ZE�K{�x������r�ZI`����#�*�hm��A��q#�����-{4��B���2��oM)�$�z�ΒdHR]k�J���D�m��I>�������,�Z��OT��9̺��۹fvv���j'�,
k�8\Wߪ�]N&�#|V�<">�1����$Ub��B�')Cb.P�;�	�[n�?�C�*��n�l��׳`�2������������gU���|���E�[Y�Iq��L
��0�w
h�[��v�����hPӶl.��M��$�/:ؐx)L\��"םD�L�4�.OB�hX#��C�����-��jW�z�y9W��ɑa7��5sѓ��r!�d�b��_�� 㻈{�1��w�̄�%�P�+�����(������8�N� d뗒	�(7�c�	ĖɊ�{�gv��9�z��!���xe��O"�h�V��L��m��s����J��h��.��u��9�32s,�F+�՜jP-l
)('ǌc��'�I�I�|J�d?s�e�]�EAׁM�9�㞶z23���x���S�H�̺{L���|Ȋ=�3w;)a#��=���h�X�=��i���ƗpG��Ŏ.w3�ƚ�:|�*���D8�5[W�� 3��y{�%@������_�"�z����
�T������ą������"�z [l�8���9a�+R{��w�����C�uE�� ����ߢ�A�?9�Q�