��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l�JR��� `��	JXK�?I��`�/t�t�稪�-JP��1^ώ='b���|��W��ouj@�&����8�Dm�)���S�������ʥ��O��#V����'Z1���㎶p���Q�Ӫ��fwv�yݻ'\�3�,��{9K��GG򂄺3�@�L\�<���6�΢Rΰ���릃����sΞ��]��w0i��]苦�����k&EP��.��՛*���mh��Ђ�v'���O|c�ZI�-����У}����)�D�-�	Q���;���A�FI���hrͯp�����L�6z~R����Г��N��t�n�"2�]��p��^9�NrG7?�	�cA�]/'�#{��̋x��,�q�i��E�w�_ȱ�����L��c���	��{T��L�4����_�:�b(x� Hx�E���..�����_!&��7(�y����h,l�c�{��
2�N�G} ��}�Z���"Q�v�d��ߤ`9��@�Y!�=����N_�@ƦK����%�q��zr��.��<�濸*�Vm�T�J�+Zo�[�|P�5jS�܀���!L�4&i��lH�U�/'
׽�x�!�7z�2;S��/�E��Hyb�+��ߤj[�7v���s'I^��w[��EY��4
��Ǡ��ф�5�a��aڬs-Y���j���fg�I�Cp N�k�X�Њ��/?�ELX���@t���V� 4C���A�)����I��R�(PL4���`D���i��{��lٖ����0��?nM{�Il��zx%;o�)W{ ��
b�l�i���Fb���\�1f��h�c���@w%����Jk������]dg_�6ry�܅]�N���-���N�\���^k��P]M����-�ק�h��i �ð���z����)�j�[�������͑����-�	��~5� �ϭ����dc
�S�Dȁ̓/x�$=&)�&�}�C���'8�8=C��%Vz����
&nI�ښT��Uv��^	:���c����ޅ?� pA=>���N�3����K���$��4ކ>
�p�x��w֖$�����DЋ����ō�Fx{g������P���6R�R@��n�]]b�(�\ >��(�	�-��,6h�����K�����5Qn�8a|U���@��Z�n�,��������t�C
HO�~�\��rx���}/�	��<��x��V߂�@��US��8�Y��!a�p���������� �U#������z���R��^,���/�e��n�Y�z)ۙ�x��~;����<�:}����1�y#�{���b��>%�c1�I�[32�@>w�2r'rVl���OI!<zk�w�&�t���|�V���/3��4�\!��̅�`�� �8-��@9+j"¡,�뮵��P۷��Z�	�I,]�w��̜��Eh�0b������E�}>����V�l��m�Ë5E
�I�����6푖Q���l�K� *lp�;ߌ���RU�K��'�Ϩe�C��Nv%�!J1�E~G��`7�k��O�)`�R�>��5i��mO0]���.%��/�":H��G�\m��!�YR���}϶�
� �<h�Q<�s��6?37�Qd%q Y��^|֫�1;$|�:؇tC�9s�o-���y�T�QǱߖj�ٷ���Oq�V��[��1�S����؉��-5�pA�߁(���3ɰ�0���oF~�rn�]��u��`�>�Cy;P�Q�"��K�ڻ�y���a�0�Ȁ�L�]�i\#l���g�,�rY�r����?\a֚Q('; k��.��b|��V�]e H���Ja��B�YUAএ�(�� V�;��N��Nk�C}���E�����Đ�}�4��]�9Q� 4�B��q�4�{��!�œa�U�篇�*N��������Rʑpi^�P藽i���o"\�&��;gM�*�șǂA1��GH�q�[۵	�HG!��{�]���A�B+wO]�
�폓�ݢ&BD~I
�ժ�I��5�6��#�r� z�9�$ib�P�L])�k��
�ZQ�g��ƈBV��K�������f��ow��d�3���8U�%��o��F�������)ݷ�W�{��b縮7i O���+�mS�)l�1F�(�͓�~�Z<?�^���EW��K&�@k8pl�L�e�Sa��Xc"��^?Gy�f�O��(��l.���8*$�F L(�p�����z�&)����Ʉ�Ĵ;Ņ��=�_b����NҶ�����M\:�`�6�Y����9ϖe�,H��]Hu���zFH�:Hsի�ucE�+׻TE�2ۜ.M"��
^޹@E���6-���='L�	�Gg�u����$�{#��>�L�%��>��B��*'��9�l����QK߰7P�������O~���u��Rs#8>�v��{G����IH�����F�N��'��0��5ak�h��cr��E���!Lľ�3����C�2�� -h������V�N =������0Yq�X�1�Hp*����%.�8�e5\���L�2L������
u9N#	
zJ��M���ֹc�@6�y���Q��7�f�&i�m�-1?)S�U�l��Y:�R��Fz���FD3�9����_���%U�H�W$Ky�J��2;��lU�~��	
9!t>��)Κq�ܷ�b�了�KL_6Ʃo��嵐T���~�b��Y��s��J'$�����LR���>�	QP���?�*����c�z���h�Ka��1�6H�b���ɮ.w���ET��fG��^̦���8O��O5�6�n�S���75�I��j�^�a�l�����1��������W�(���ț�?�8x��1]�@|c1�U�	���|�d�Q�D����Wϰ�M��#!�M��pR�H���#ѶZ�H��]}��QAFlN�m*�	Apyy���uKK�8~�dB���+��Ͼ6�wP��\?
��2(_�5�����b��(��9�4b�VG*͟)r��c�I��K^��F���:��R�g�G��8��*������ W�������s��t�Hf���a̗�j�H�r����|`J�����B٥	�r/��!������&�o'�I_�'^��.W�t<J;�~zJQY���d5!�b�j���s��忬��T�l8;ߎ�����Fax��)�R|�p�f�)���\f�8s��5���)3]9�E�A�1-�����҈�L�/G�3���11�Ǳo�,��@�<��3w��m��,a�vĻL�I����.�W�sT7�ΰo)�׼O�,�%8r4�Tqj���,����B������c�f$��W8!W�S�����]'#��ϊ`6������Ox��M;� ;n��1��$��N�x�g�:���l%e���3"J]��o��!Yy��%	`�/�:W^�e���2�R&�M7�F�U9����&��>���N�p=�I�a^�+�t5�z�B��u?c-�\�߾��(�<��F)�ׇ�$,�ց��� K�D	�>���D�f�N#(4��ڜƆ��%���Qo^��"�/zE<Ѐ�#�%j��@��*��z�^hE +�8�[0��d��r�#AѤ��������w��hQ���&�N��(7|W�/q\�?�y�0�t���d��փk��s�Z쵦�5}����fU���u|ٗ�.!C�&'w�ʬsh�3g��ғ��*�罩������p��kk?��c�U�۪����KU=����A��4u���'ܯ��S�q�X��ڌ,��s̎��FO�(j��y���g
���9"�K��mmSբ���i����K�"�ן�'be.!-��,��Ĭ�^y�G��HL�w�"�`�던��@�H�MH��J�#�K�8�<?90��|�0�=Xs�5c�6�BFU6����I�Ո��"ЍAH��v��
������	�z�7u��F��R�I��ļ�K��Ju�9�v�׈J�!	k�� ������M���5���_X
�R��k����RU��8)l���Ҍ㈑��Y��o��}�	0��tFM��.��"G��渳̞�;ʝO���
o���|)C  <ѷ̻(H<�	QJ&��1��z�v�w�~�c�n;ο/fe��#1؋���v�%�*���ם�sA�o���\A�)�7��c�k���8^N�橽i��J��$��)>*�7�8b $-���[Y�ɗ�v����	"P��ʺpN���`>��+��@���4��9yۮ��/��x��Ki5��k�����T-~���ު�x����O��?������t��}���|���{���~���׮�Љ��wiM�xbU�kz�����xcv�|~MXO�=��ck�����<1�9H%F��I"5�QB��#*�Ӂ@c2�ɟ��fLQ]�f�4�o�D�(�~�����)��B=U���yE8����p=봁��%��(�)��e���M�$���Luʸ�u&kҿ� t���AlN��6�_3� r-�ˠ'y��bY�3u�5& ��~R�pN��i'!����:rmE[���[�Fw�<`Ro�,�<�V�$g��ww���=�*"���w�U��w
��Zl�i����	o �r�V���7�3����Oz�Y�Ͳ}�׵�R�_�����qQ4�
+�[T��V��E�Ф)�}`L�n�n��K��LNP}ﲡH.���ۤ�6�=N��d�!B!I����.�4�;4����cb)�7��ZԺ5e��KzR����1f�B6��䓋��<��Ͷ���!vR�;�h�,P��Q�k�N��0��