��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K��y�rIg[��?���������.�%75�N��1"{;�3�=�������"-9N�!o�C-��`����ܩ.�95�4����e�s'����T�*Ճ}�ܘ�zt+�m5Y�Ov3�\6�S�-�Wj�����b��a�d��e xGp`�q,����6��&����J�(2Z�! �-��=�fX�T�\�-ƕ}��Йo�V6gE�|5a�x�)��2��+�Q!�Y�2�Ը5��� rҊ"c�/b7�u�u��&8�[y���*Z��#:i��s��s3�5�s���g֞���\��T�������W��V�q��8�do��8���/֞�9T?� zN�ڠ*"_5��)mW�@$�I��-�����åZ�k��qԫG���r� �9~SqV-�C�KP��q9t��b2���-���S5�' Fo�M~�L�+G�����p��mn`q,	e�P��5���@���a�[>"3DzǋP�òB�e}9}��mv5D�ħ�y�ݹ�� ��1���t��}
��oSwe�׭t��F�c�rq��d}~@�ު��}]����D1�;>��ۋg%��># P\��|4qEK�'�(9vF���
Ѭ��&�όVg�k[3����nK���	���X�R?�0�sQ�)��?/͌��rw~T�����]�{-���[)$nc�z��g����F@&���|.��>���p}E�)M�q�d"y�B� r�C�fT+��mV%�տӚ.�n:�ބ΄�ʞ��@��� h;���D��gFz�$���mr����{^�<�V�����w�ȁ���^68
�b�b�OqG;S�9�}�w��}Y(��u�	\�ږҷ}J���Y�L�y�FΦ=GH/� qQ���Hju�,�TSq*}-��$����	�Օ�6q���<���o�7��΅ʂFی�^ټ��	���D�����%�抗�
ݨ>]>���Fec��I��z)Քo���%�ˢ�����B$ޟ���������Έϊ1�S���:LU}��Pms_E=68�.��Ԍ�%]A3��
qƗq�B���������̚�}ɂ��G�s������1�pfK���X���$	:jV�.}����DM��)ܳR��?�ȴ�����?�`�m7W��V'>����G��>t̔*,]]��tG`!���]����'��>B�Ԇ�wuC��ؑ�����%�AR?�NT��&eY��l�ȴ-���Ur@5G[�uM"�u��PѰ�t�ۖ��:HB�7���$�}�V�%�	ZN�̓`�D�T8�p,pp~�«A�g�N��"~�1�M��TZ-�?�J��ca}!�-�^c�j�
��fm���d���9s>M�a�b6����P��� 0V G%���ќl�m%C�5wOa]
�����h��x�.��9�Ы�O�l$�Ξ�4�+�����s��b���Ƒ\uR�oq�*_�2=3�Ɠ�MU0�f<vx�E4<D|�}S�U�^�l��͎���H�v��ЖF����!��������a$�l���Te!�5	��d�y̨����Y4i�y
��M����ҚM������uѵU�p���m��&�Z�h,�^��W�lb
��1[<����_�?�3���Q�qJ<]�<M�tij]��#���2�yB9H���r��3S�.u�1>��<6ۑ�f��W����b�A��J�墁��CQ�zb%��H��6(�r^c������u��x."�p�Û��}�[�����D��<{�'c7)�+�XMk�A������L[���0)8�Չ�o�7���D��F�aa�Uy{,@��0Ey�����Z���x?׀�)�j�R�ch��Ż�  �V�6�qKB�Q�x�� b;�Y'�a��!�EV5�8\�x��9Ը��/=y6.������	-���р����R�j�;^-���cA������1e�����	
(�Y+��-�	���~+A�:-_�*-�P�+��LF`Ou�w_nS�BP��E�УA+n ��x�8���H����0�;iMS��;����hH�D��Q�ʦ�����8�Z�VSe�@��ΰ��P}XY�K��K$�9��b6f����]�=���L�a�0�]x=�
�����l��1��Py�m�Ɂ	78�<{V[�؜���*kayJ/���\�:ڷ�6D4m��Wz��$�n��S�7qPe-mM����R��v����xgH�j�S����8�[��9��C��P�FG�_������L5D�|��(���7��1�,TBz��=����7p _4�I,L ��嚸��w��1���X��q����V3P�'>AIĻ�3�M+ּ9�-��� �桦��!�{��PU��5�k:`�&��=u���D�B�r��{Y�!��w�C�2cr��x,Ζ�O���kp��������Vi��y�MF�P">J��-Ѧ�O/؏�{� ~�/	�ψ
�2YӢK��ԎD��0�~+��i'q��X�%0#EN�ૺ�zM̹�fXN&�n<?=f.�@_�#��YQ]7>KDWM�|��\���b�s� �;�o��H�]��r�Q����[p|������1�K��|��Bme6�_�e��� �5�t>M]J<�#ʞ��ڬ3+��a�F�U���x��Be�,6���Ô&��GE��.xΐR���7d�J�\?�&)3ΆZ��:5*k:�GV��9���,N��Ro�R�w[�1��ҼR_
$R����r���W�,���E>�h|^�{�㰰�8	�<�\�ц�]Y˘�N�n����	��çN���"�o���*��h� J�� �h�l�@>d��j��H�TO��82�,�T�~����|��^��8���ϝ�$PcᑟUl��z�r����w`�e���yi�߭�4~g
����_eߒ����?I��1�C�gY�뜀̙�<�A�wFO�*T�δw�@h��vM��{��Л*���AQp�-z���wɢg�C��t������Ae`����]�,;&��?ޣ�%�!�Xɯ}%�B^�2H�u����H�Kf�����X�p�`�w�fA	�F�c����Y����Ľҿ�Nrk��G*b�
?����*�B�5�f�y���[w�&1KNC�Vi�� v�Z
�	��?�=�oԠe���I�09Ń ���Mf$2���1�:�*�}Z�|�p~�����>�� $���7�������J�Ľ�N�����3�GAz�Ʌ鲉-e	Cl�v]
��r�R*rXX���C3�b�xO�7�j`�]��ؔ��W�)�7� #���0�g�.R|;Шj��9Tz�V�ڞ|]�Ө�oF:ks|�.�̠OҒUS��?