��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���۰X�cr��	ɹ�U�����60=�ܱ2��-utTXfϕ,��r�ҍIz/k�T"̴�2��o>�a���1�.��n�~�ZIc��\�2��,���Vj
-�NU��&�m�T��剤��&(?\�i��V�ӌ@�I4���vd�����,if�Q��3|�]tw��7(��zzݮ�CO{�դ�L�h;8،�ֿg�v����ӄ�9R�*�R5_2pw?�_���{rf�V)�2�;p1�Z�Ŗ ��T�ߧ3}_� ��O��I#�m��o�O��kxv��ި��3���ӡz^�-$Ǟ�ʶ�皘�u0t$����z��jSU�J=t��8�cF�.��\�4�Q1���Iv|%����e��	��g@��2yb��+�k�+>��PπjtMܥ�Ξ�$�	�����*��.�g7��V�R�N���3W��'��Ga�5��u@�e�D�v��.���5�΢�ˮ"�$WՃ��k�B|�����ל��WbR�= �d�_��W���Ii{�ed򊗿NQ��kP�����_e_콆Jc�T���,�ب&��AS�8����y%��v�7�|0�ێA�
�J����μ �A��F��8���Wb1�=n58�O�ep�F	��\��'Nҥ@�&G�� ���{SzQ3▸��ce����ɖ� wKhRX��m�I)���8���
a�1�z���դc3� sC���������؋�ՉΞ=E��њY��g�}%�ܷ�Әo��o����H ��4����u��G��J��&�]�]��>Wm@b՘�:@~�l��ݟ~�eq�	��TRw��,��a��^9�gr���!�j7��;V;I1(����֐�������5x�0)k����1$���<��CHI��gq����v<�a�Ly1�㈰v;ٔ�v-�bT��)[@����@�dfz ��2�� �����d��PgM�nͽ�#'�k^�oJ{��)���O�Nۍ[�n���ٴ��?�e&+��֤��s�M��?�/�!��z��X}���:Y(U�S�Y@�S :k�2Č�rN�-���:���X�f�`�!�����72�Y�&ܱ��J���D=��C����T������s���`Kx�f���/p�����S�jE��z�*��*��c�3�h�B�p�q��=��ᢵy��i9H�+c¼KlV��}�%Q��F ���ٞ��׋@�ֹ^m�\���^�ǱGn�QBP�
ma�l-:��,�5��r���\���q~v	#br`!�d�){ E���1b$J�˪6!<�|XfL
�WSE��	>Eo�\����G�3�1@ƴ	�)q�-$�����(����3��Y�`:�f��f�	�c��e�G�����IX�>Rz7�T[���C�ms�k����H�����n.����2�#��,������V:#Z�ڕI�g�5�n��%0qY�)��mI��$A�l�-9HU�<�(u6a7N>�[QCr(�EX+����eP�_K2����=#ic�}}�g�q�x>lSNl�o��9V�j�/'���� �-i"C�F3c�of�d�|)��<^H�TXS����?,eL�
N!l�vGf��T̶���!�>ye��'��p��6;��ap|_��]�B]��
4�~�J9�b��9V���O���:�5@��D+��h�k!Mٌ��9�>�R�߂N�aR��#~�Kj�ƥ����)4x��4c��o�:J�_��<�=���u�q���h�BS�<<93���K�����Z�p��2Ru�hPb�7W���H��d*���:10��qv(P�ڪU�j|���H/���!̌���c���",�>L�`Q(A��UnöF�H �c��`̓�w\��w���n�.�!��-�`�T��}]_��_}�4���I����.�3F�F�׷���
΢�����](UԷ�yRn�*�¥�Rsq��*l�tem���;}V��I\@�&5<�d�ɐtI�J_F`�f�RL]|���JrWO��P1B����=�=���S���m+�8>���
	�b�k�q��G���$�7�e�P�W����-�nR"D���Jz��qZ��
!*IpzG4�P'
u�(��&��_�λ�ޑV�%�<�~�V�e��"�!r��f�r��м��ǒq�������a��x��F>��	J)���ڛɸ%N=}�+����-J�n�:ɷ�mN0���Vi�%#g����J�ֲ�|�g�����W��K{{ ����7m,�Qy�M�[��k*��b�����E�=����g�WR��`cx�`

���ҍ m~�b�p5�O�I��Aj�s�;e�kz��"@��;�k�{�cP?�jLuf�hn�&�?B��yk�=g�cd�6�u�JF�׊��ԩ]J�n�q��,&D՘�.OpΔ�j�{D�M��u�f�r2�LB�Q�Z�<�z�:'��UQ�HL1�Ҍ x�'5�u���sunD���|�%���x��&�:�<�eo�����V�:S��|��X�x�}B_�����|hsy_=�V:��u!�Y~�[P��! V�<��A�X*&���hFp�H0��]�F0b�_〴rF��]�2�K�&i�N:k��C���v����5A+�W��h'sA�!4��X�a�`��J�uHI�YI�A%��Th�@���DK>.���p5蟓�ЮÔ(��Z�Ŵ=j�2���@5V�>�����Lږ�{g�Η�����ȴ�њ�$��(/W��X)�&Z" �����,Y�`����-T�qĤ>�ysȧ����Wu�'���JHV���@�$�f8�T�� �T0-L�bW�������E�O^��Df�T�	�Yj�.��^l�/P�)����{A��/����&�z���	K�-sJ�BP6KnL
|Ƽ�S� �Kj�M�j���a�JR��aR̕�����/�g����㻈@����D�N� �\���/�ͳ�����ʓ�	DV(G�N��~{5�_���MYh���܅�z%��sԦ6��ꙿy<�;��e�]�����1��Dߌ?'����L��7<Ah*�ܡ��H�
�$�\�M&_�%S�☩[��3A��g��V�D�d�y�d;����WwZ{X:6p��|��h��'����&T����H���*�]� q)rh������;,��Ǥ%��
�v��Xbȓ��6wh�u>�M�]����Tft���LS�<���[�Ӎ�0�����/�S,Q���/�L0�U������j0�T.�`DE�O~>�b�����p�p2/@�R uX��u|w��0�b��xS��qDD�����7�?�vQw��6��'�"r��l�
b��P�ŗ���ݲlQ��0����}��4�j��v�g1j���O>���H����@;y͗���1�1q82�v;+�S��b2�4�Tl�f;�ϯhG�~̄Sy��
�/��,�,���5U�K�_؄���}؁�A4��Pl��=�<n"�6
K�vUbUA�#������?k2�T��<)�J�=�"�M#�.��y��i�-�����s��\if��0�*���6 +}��_Ȏ���_u-���?�g���י@SSL�>��=6q 9v��^.<��//%�
�u�r�;8~�7G)E�f�N��/��J�غS|7�,�ݥ�# �R�thQ�ZA�G�]��������^Y.��K�	�0��,>+�5{�6'[�_3��e�z�;.�֊?�n!d�Z��`�HAuظ�D�����s`�4��ur䥆��<Q5�-H��t���"�Й��r��by������Y4�u��h`	�5�e�P��و���	�����Z��Ep'���N�}�k5r��K�g� �?dlZ���.[�:�k
�c=tR�u!�hO0� jCSʵ�����{h�����kv�/�1�
x�r�Fȫ$��E\i�"�4ϾjBV�R��|yp5��ùT��R+Rm�c�>%нe��؝�����O��p�mOFJ��})�&'8���P��3�0���@�."����q\�o�@���#��:֨ۂ{@R@����/Wː=��1�؝�PD^c���LR��o�%�\�q��٣��J���r�yà#�m��'�{zR�����!0�~� �s��4�r�-n�%a�����|�:�$�I6l�UQ�Lۺk�z)��5������-��ӳ�,��d��)�A�NC%4��}�����u�J� �HЅ;�G٥!o����^aY�X�;�͖PwV6[��=
"Zj<�S���x�RP;_lf��m�}�+�_��C��G�;Z ���[M����[MT��*�����1:i�)�<��ѷ����x'�'R��*������ ȫ-������.�	r�č*�	���D��g)%|�������eӄ�!�#Z$��q��\{�ae��Ԉ��L�1c��YD�/�/�������:�XWuA�9c��?��<�a_�6��ޡΊRڈ I��!� ���H��"���_��6!ܶ�k~�<�QF��9h���ˋb��
^�r�:y9yZ��_Ӑ�����~O)��ȫ�ʪ�"�m-V*� MpC����r���!.����_���̍�+�V��$pO�L�A��WX�Zv��s�p���O��"�ƅ :�.���#��rBCɳ���>����헆���n?ը�I�W�Ӳۉk1@7�j��A��~';
w�Yʿ���P��J󺽆<���l7X�����PߪD����޲3��tB?��w^C`Ym��8�C�d�X�{�而oʉ&Y�H��Jp��(�����~�R�p���L\�;�W�sa~��w]�b�1'��C��b�_�a%�P�tՁ{��4Ep�Ə!��S�,�v��~G�X˒ah��N�Ńş%n����5[-=�q̯���6��SG����"���w���g���H��E�����qpe�@$�n���@���)��Dz+3ɵ.�̗jK*c��΀&Y0~�j�>b�� � D	��2]�T�"=	�Jhl�M�^}�4"iJ;)e(��o<��<��j���c5;��tOc�I���j�e��L�C�x�<�&Ķq�N��9+�@�}L�_�H��M�h ��"�͊�����9����z�}�m]e��鄴1�ue�w������UG�7���`�Г��y@�T�~�vYn���/���۟(��rt�d��R���&
�:�6�>��T���n5��r�"?)KV����j���ۭg0]���ͼPs`��hP
wJ0�V��h��l�}��P~�[���MZ�!t4t�J�f���P˝;<�J&�m�e:��o[%M���f�۟�6Q���ns��n��yܝ�����\�y��7�i.����
���>���y��Ou�%�q�<n�R~�7�osI�_b�!`��$�L&]��o���k@�kA�FN:?л�>�Ǧ����T7M��j(Pb����&�>�zk�9��~+�B_t���BK�v�]�Z̟!�2��A�i����g��e8�D<t�Fy�َ3:��8y�w�Q��Ԓl�{��9���T�YU��w�O��Gw�����z��Ɛ��Ҡ#�d�S]$W�d����R'�A�����;�A?JWQ�:�PC��F�'����G�c�+O�.���� �H��M���,ȾPw� �N���YE�&R�7�G�_�fW`񷕗��p��R0���x�IRM�F�EYa5ֲ�P�1��?����m:����3���#3M�+��[�5r�D�`�_Y����x�� T?���|�A�f�ɚ�����h%r��'u���Cƒ�3���w�ըG|�7�IY�kB��n�ʲ�"�NA�����gv��*�@��J�����t�B�5�z���[b�_�J`�ެ�����`ێ���Ί��Ҟ��P�A�m���I��Ḿ�[�v�T**E���,]��8vU
�g^(�1O���@��qjJ��5���K�*���f@ʏl�F��D�\-�od�I]l���	E����- �Wh�f-�Y#�I�b<U�e��/a�8I[�I��!��O%WJG=�nxЉ��x����e����8���O
��J��V��y���6����Es@EXL
οX��'��I�����6����$'\O�l#�P �+����f�M;�/���H]�7B|����k���SԮ��Q��j�v�7LLZ[�����d�gNo@��e���w/��^�ʃĊ���"�O4c����z��Sqv���^G%���V�\Y�����$�������r��^,�'l/F�� ,�K��fvw�����3��K�8F
H��r�
8��$Q�Q�bn����;��� '[Tk�{��!J��B�]Z�f,�Zb"<ZI���R�2�T�DKOHC�	�#�� X���>ZY[iFs˶�I�|��<�v��t���tO��*
�J��.�*!1��"�Я�R�t�����*�*�jk�x"B�
�C��`�[��q,�F��I�$cGAr��:}!�/���ZК��઺E�`+��A}I�9�,n�$�0����0�#�����d9���R�mp)5w��G5Ys�T��Q����
�ߨ��M���!��;2���W��ە�����f(H�必s>|�g^?Կ�x��k�W�m�毓�����sQn��T��7�Py��w�XCX&�����r0Na�V-��]�,�~��͆V���,zB�_!B�{�V���ߟ�Č�طA�����RǉXs��,=��
���9����Q�Ŷ?�~�U@� �l�GX;��=J!\��PS��LW�����).u���O�K�C�u��v��J}��8-��^�I2싿�_r�̞F�1<���;^-@F�Ņ��S�D ?�.񗝕��I�Jc%��mܸ�c흏G0�k?sH��C8��W�q�\7��I�"�l5d�-Y<�պe�?{|Y-]�����nP��3԰!d^��Q,Yj�G�- ��?{���3w�*��X0R����tf
��|���2�yi"�3Qz�y�Ͽ�%��L�c���ř��_�s�b�P�^"�ȯa�@5�{�CO+��g��,Ǘ)=�R�.x4�]�������=Ht�<�)�����O�:�­�_��a���E���h5������� �ճ��9ۈC߉�숰�V�~��fC�m��w��-����,ԳN�(���b;+\ڃ@�%�u��x.%�x|�����5�*����Ƣ_��w�n{=�Pˮ(������%�8.���1�r�0�y�I�,kӊ���B�έvH�pP�����#���4���NdL쓇������
ݫr���xac�X�P�1T�zW�����F�ЪQz��v����Q�_����"rݷ?��?�b��}<<��>�-)�R�1�P�6�폡�����1����a��lU-W;�~i�6l�"�%�ޕ�r۬}��6y��*E���!�C�����)��Ɍ�L���Ϻ�u�zY�}q����y#�Mo?N.��ĕ�$o#��,�Ì�u�S��I��J��1p#���[ŪR'����z�G?G�_�z\�o�N�ڗ��7b�h�����������	�*���V�7��Oi?�m&I�����Q�6�	����E�W����k�
>u�����Aњ�U#}���Y��t_�U� �by��J��qú#x���]�J����AE�|ʬ�CK-ԭ���J@�9���4�����Xh��H��� ���D�(�M1 ����(ק߽�'�����,�<�Eف&�cU}[@��R�����el%Q�� ~�co��:|�OS_H��YM��6viUeT��Y������W�s
��js-~� #sU)QovS��d�.re��)���^����zӋ�I��Q�Kvc��Cn�&�:r\gD䘨%F�������x�ه��ye����:r��U!l��M5�8X��2�q>Թ����E����~��M�b�R�y%-��ɠ�����5~c���=�e �M"��@�ԄMg:r��*R��j	���$�s��U>Z�� �G�8�bL�����/�b�ǆ�;}c��� 7*r�Yc��*�5h7s)�9P�3�}�������]�{������Q.��ͤ��aB� â�	��E?;9�e`[��4*;���b�S��H�D�0d�F��~��m�\�@�K"_�F����%_��H�=��d�����'�'�=p��;'�y8�����u��)L� ��6d���]t����(�V��~��Ε'�|�^_|Z�K�����a���lmnz|!�D��������W֘O����{A�׾�I�ɱ�5����	]�6���ƌR����Y���vw������Aq?tI�����E�%�?5gd���G�'B̓�����N]�s�MzJ�`x>���⼱*}ْ�w<8%֊�]+���8�y-�L��Wv�ݠ��l���#�lCW�lR��)�L���5_^�&����M�c]� v;�`��;�����ךK��ĕ��6}@x�%J�*��^`�)[�Giv_��WQ���1��V��Lc��-p|V+��G:�[CJZ�%����f�;�f���W�ٶK#����:
���eK� s�P�^��m- �G��P��qZg?!iY;�M}����4.���8���<�λ���^�]k	���뢖����M=�=�҂:c��K<��/'�bv���������"vE��cSS��ܓ�TQG�U�+sbK�`"��KȀ����g7��>H8�z5��F��1�Հ��3Z;j�^/��PS�p�����z�%� ����0�P_j�]�I9��),�B���$�����I!��'����~�2�b��h�$���DSn7Ĭ�PU�����9^�\Z��#N�����������V��Xv��U�s���鳄���O�D8R�{�2���s��(o ahR����)�f�|�j�y�ZB���sh��^�0�m'H�^̬Pa<ݮ�f�"�/6ʶ�R���	,z��HӕF��?���7V�:�;U/N��'RP��XM���Aw�	R�9?rw�">J|�Tටq����?#��צʷi�tJ��ےW���,5*m�u�o,:�*����\}0�j$N��W�e*}�[i��=��$���l:���7S5�Nވ�,}Y��C�mR�@�YON�Z��MD$��Dx�ɚ����WIT
��?���,�uM���2ա8�����2ܘF	��-H��
�)���PT+�IxCw`ZVk���^���b�Q
�֚D��m���QR� �8x�ŕЮ��T���l��9�P,���P�Z0@�&G'>�	Ôg��gN&4U�������~(
��ϒ��zժ�ڕ��U��b�u9�J9� �=c��g-�M�7(]�)���6��L m���m�MLҴ��MY<5@�h����uN� S�#~Sy�U��������k36��"�o�wE��Vvk���V%��j���F�M)9��E�ʩa8�E��m�g����䞷l���"]\�iB���̌��r�E���)Y��(潥4�>��:"�-˥D���w�b��,m`���]M}�B�1���D��Z�?��K�!���e���$�-�lQCB5�͠"3(Z��J�-_s)�T(F�7Ϭn9z������o����~17��!����z��3���j;��33R��֭V|�Ce�9 -4����r�J�c�!;�O�T.��;�o��°�#W'��7_��^i�q̮N�u�U_颲L2�����c]�3b�Ͼ�}�k�8�rr
N���T�,>�_ Kv�4�ۈh�J�5��w�m�q��?� {��!�B.���(\G��X-�ff1@���a��0�M��{�4_R8������m𙭃>]߄��
t/�$7�s3��d��Mm�է�O�&��&�c�fbE�Z
��_v�\�
jP�.e�gyR�c�$��D����.��n��Q�+�ЈȈ9Y�p�?`�s�6�A��d� �^Ԫ��K4Us�ۄk4���9k���\�M��C�}R��osĠ<ic�V$�����ʬ�I���!N��ƁE�L�Y�<k=�bx�S�I���8%�U�����+.r�~����/��_�fd��Ax�!��D�k�V��06��[�Qˊ�]�8,�A.(� ��j����aKYD��_t[zHe�a�a�Ps�n%�L\HCT��m��}B2��v�D"�g����Vp�MC�I�9H[(�|��8�E���meRMo�E�$�֌bu��D�����x-�=�>B��P��v��y�j�ҎM-�p�y�;��G��^8��܄�Z(�F£>������O��1n�`��4��6�eQw{�.�]�Yg�Fe(eN�
�������/�O��O�,^�^;���a.��4�P=G��ǫ�� 19�-E�4(#o����N��H�}� ��:����Z*\8���P��g\.��χ��4�	�voU	�·�>%�7��㡼ǣ~WJ�ƞ�J&��\Y�@*����4�e�%�8�s���_=�M�σ��-�,�iS//n<u$c~�d��-�+�S�,>U[,�x�=�E�N� xe����I��P$��&�(嵍3���Y�u)BN@P�������,{�҈D�?�y���R�1�� �T��="N%U�鷓7̮�d���KI�j�����MW2��޲�<���H\q��ٕǉ�/%�z�$���X)C^J�
��ȍx'c�`:�6�f}�
LK�u�������PMU���G�b���Jpy9�6D��>ښYrJ�Dl��t�k9�Ģ��ۋ�\{!��8�`�Cyv����܍�T~��K�߇��,n6�d���|cы��
�D����Ay�o����"�8(s��v��P����זZa�4-������#��{��1�g6	L����n�|�@D3�Zc����|>�2���)K��ڞ}>/��b��\���7����4n��`�8��hbTJ��9R��>[�IP���bV�'�cO��^� qqۊ�����Q�k�ɝ����3��i��h�TKP !�� ?��V0"�]�v��������T����z_-��gI���Z$�Y�N�/%n�FE:-d��@���gn|K������!7�_n�I�u|�S5s�P����D���E�<}�**�Rj�=L�~�$���!�6������+|-TeoA=ʦ��~ܫȧ ��j=~���)����O�W�d��\����?f�M�aq0\P{vV�˵���Bc*$�V�?:K u�m�1I؃]7#d~�9�A>'A�ƨ��t�̚�$a��17�X��c��s����v��F�p����@j�{�nV�9e�RUD�|h�Y=[N�� 9ެ{ә�n��e
 &SL�Hd�@��lR��jc�E���0I��:_�Z̖�%�q�v�����8s���Ǿ6i�~��e-�+��Q���'@�<R'<I����T��ko�D�`h�o���_�}�{�rMk�.m�WPk$�EP��,�WsM.�l�,ezn��TJ�
 �t�^R��Zr�ĜP_^����o�4)�=Y��%��8�wQ�ɪ� �Xd��x;��p�(��v��������֞7R sɚl�8���G[Jߡ.4���Ė�A�T���ܟO\��^d- @�r`�ec��&�N��_��� �%9������YC�C
SRI,b9����i�.���5*L�2r�^�]�g�$��]	��M}�`�x��#�����UZa�0C���b(�C�峈��}N�vbZ��)f�2��С[�>��~c�Sdg����Xє�@[>eB�[���k�r�ly�^Z���c���UY2ɉȺ�l�UO���!�_O����bfu���*���\<�;�k{�1�3ωf��:��8��7a�dϕ����m�$��'�����0u���K�%�ҔBמݻNpT�m�
4�0�LOC3?��������c�`h�2.Z��↎�9H[����.w���j0�.�x�YI��y���O���W��/V$`������K�o�Se'���$�rĖ�Y����Bi)�P�)���qZ�C9f[S,���<��+S�X�uv��Q�1Hs�k�w�&���O��(-�a���4�7}�V�.M�۬(@�q�$dBJ�a�dJ{x�>����BVp;4��a���N!�NZ���6S���ްD $E�l�3�p�[S�Gs\I]��U'��+�ش �9�U��P��R8h�m���Z��=�n�臟B�e��Ĭy��SN��T����1��Q	�����ĂS�}n$m�����l�4���� ��UQ�Z��ep�4��%���c�6�������rĿ�b��yxE�ё�����M��;���]��D|���\Qk+6�L���a��]y��Iw�T����Ǚ������1)���!�m6L5q'S�5�˫P���_�������j0ak��|��w�p�>�yӜ�Oe)�F�lh���'�c����f3�8�'�e�T>�ى�Df{�U�s���CۘW���o����r7�B©�c+������ �	��v�l��?�AT%g�U֛�1� @�,����W�e]�_J����O����ip���!>����푍��@��������z�30���u8v���T���2���2�7�zS���c��k�m����[�x����v\CM�����ܦL+NX�3�ڕR�!^$S!)�#'�tl���m9��^7 �]v������ ��ڍ�m���Y�8ِ���;�Tb�����m	.m���a(8#�ӆ4ǁ�}�fx��h�WvR�-�V�U�'	(�V�wB�s���*>t�%g�n�݌��5{��&���p#.��ļ����	ybFz��I�~�L��>]lEo�e$P�t�1�.�d��:۟��+��8�_�- `U�kI�yo��ʸ�L`�H��t�G!��e�����c���o��ps����GȂ=����Z��L�W�`X���v�+��,e�E��;p �"��2kH��>�rk�U�;��7�20��(���k�~��y ��@h���fT'��Ւ4�X���*�yDT����-��@�mc�=|���l�lE�sC� �ØP=�+4v��;�*׬\���ye:84����@����%U�,f*I0ˑ4Q;���"��n}��_��^i�U���VF��/�;\����Um����1B��90��o��ru���\KF/9=G�D칮iz��!"��4}=�a���7zA�d��9�$�ME�}�����JjuM�o! �H�^��G�<-� *�y'�u�rc��*�7�`�����sK���n�ji���qcԗ�r�X��߶��x�m:��)�����ƻ��uzmcC�{�U}.��`3@�S&z��s����9������H��`v&������xD�F�ꨢy5br���]d4!�$*�t��W���A��6bm����p����W�
j���wn�0*/-�(\�NC7*@����o��
P^���% p5�{{	j2��ؼ��$X�R�Jš����a�����
���ifB`��'�w�wV7�q�Rp��V\"񿾑�(-}�E5�Q���-���u���wi��=l��N)��a��y�J�e�[�"�18�>|���In�?�&�(��Ѽ��0z�;B���e�?�CH��(�/z��l��ת���*�?�>1�B֜9��";(M�-P��)����ȇ;���7ԫT��N�䟲�P�����P��$PHO^��1lYN��R!g}�pi�%*�bI7t�*�s�X/����a�F���O*��bT������u���"j����52ј4h�&n�Iu���*��c+���\ZN�?��%�&�ᨳp��n�
S^PX_`x���b��?q̃���dr�Fwӥ(:��Ɉ����Gv\zǍ`����[�|ԝ0G���r��por�.�@PP�b`�o��� ���SW�&L�����p���ӪuA�y�n���@��&=ˀ<�� �	0z��AQr�P1;o$�򓯺��jk�2bB����OZ&cO����Z
��S�'�hL��n��a�e�>c&w�c�����%1��#�d�&�<r�#���{�-�Fd>���e�z�3|��X�hz���'��m���gnL\z��&��굼E-fJ��Ia�t���l��9��=C�P��jI(#�qQ�·3��C ��)�a��;�� ?��~z8s5x����{˚��g��m����y�خ�����aQ$�~k�W�&���~%c���VN/i)����?6iQ�Q�n8��q���L�^�"��<��Km�K���%����_�?��#�^�c�;i�ɸ��t���A.�$�`�:�,��4S�?�.U�+]e5��XF���16���!\B�N�ʿ2��2�|���i1<���(��Ðr��i0��f;��k���dt�&$�(վy��^��تJJ(�	�'��t�v�� �y�ȸ�˦��wH^���( �-�o���	9�E�p�@=���<ĕ�8Y�+��{����k�����wd��e�\�����3G�����v�.d��-�z{aѕE�NY(˱=@��h!��LBj�!z���:T۩��=V�4�۫D=]mUƲ�b]�!�tY���=ZE�R uK0lR��o9�
2���%��9����q+�e��~ Қ�yԏ�e����eJ��[��̒����T"n,a�c �$i�I��Ǎ�P�w=���&c	`��c`�{X9I �{<�XY��sO m@$�3�B�퐰�z���j�����I��lܡ�r��N�X�Բ;��5Á[{3�>�\�FQH��oZ_0�'.�<� (Nȵsc�OZ�N�M��P{{���V�23��:�OL� Ơ���;%'w�`·5��� A<�=xv;�V���w�-�P�Y��ai���c��s0�V��|��%�e���:����ն��Z<�/3���4b�ŗ��۬��iq�o�u�����V�sF�rM^�Z�` B*��_�f����(�C���a9w�|8۾�O9@����
�>���w�#q����3���,/�	���+���������]A��&�S��o�+N��W�? �"�(.k����YQ�p���%Rn���	�x�.�Љ����E�Y���jˏ���"��N7ܴ��%����9s��G#��CgR~"A0������1U�7��(Q��e�GWؽ.s�<�� �mi3��]Yyl�I��M!���B�s�f��o<~S�`qA`�Ƨ�i^���i�
����`�T��I�� �٩�`g��T��׸��򟩉X(�0�@[��Qd<�<pi��*�n�*$:�x����$��ʹT����1� �,��$f�C�B��9hu�^K����N�����М���<�Z�f���iE��<�֏f���/�Q'�H`�?t��:���q�3��:~��7ϋ47e{ۮT��$7�D���h�-<y�&��>x
�d��%����k�~3����s��ŷ�-��oΥ����X�����8�"���q{6 �Q?�ܣ0�f�i9j����8=��0�y�D[ tq�)Y����}5��~CWB��Ш�̡�:��V����[9z(��Eߚ�u0zųG�j���ЈL�����$�!T�pB*���8�M���a�f�vu�[�b���B�ǻM��oC74�O�|[�$\SB�'�XS>����d��V�6C�J&��yADf���a�<J%�@e.��g��c�u�T�CWhG,i��!���H���{��l�%��'V�[p�W���r�ݘG�-�N�*��8h�O|��ԡ�u`���p�Os�V�a�����:�_�g�X��.�A�#!2��JIet���VNo����0<f��7�fc����¢���H�@^��
["�s����/����w}��:W�MmB�eC�����^~����W�7|=d�+�d,�TR�pk���mg5|ϗ��Sm���A�[U�ڦ&F���cA�7ı��*��'�����`�@�XbWb�	C�V�b��j(���~n��bRe��P��#��[p6�̃��?ٽM�����,����Q�!>���c)�Y��Oq%��.k��m�2�%V$����d�,G�_\"{�~��ab|���^��|*׀Wӆ�f^a3�邨DZ<�.(J����a	'�(�>��;�QD��u��-�Bvj؁���"	�u��Z?����(Rwcjcx��@h�T�|k"�O�m��f­����)L�[����8opr�D��d�!�i-����⚣��k(6��Z
��9y����}�a��z�%ڈ㖬��-1�v�#)>�P�/G�Ұ�2�x�9U�R��M��hY����qh�˞7��9��/<�0T
S�ar�hn���q������_u(wy;���<�WPDC�����ΘL⤩�dߦ>���ZI�8W��ɹQ���!����j�P����X�K+J��<�oG��ˏ�x�J�ז�#���
C��1!��ۻH#�c?��IM�. o�dݒ���p��jG2��dU|ow���q&�Ͻ��y<���-�m߃B���{M	��~��PV�s
�+��&�.(^���;h\Z�j��-P����D٘�T*��z�'��ЍV5$�E�*h����K $�C�|EY�3���'_��d�Tq��&���m��m43>i����uJ����6�Na$#�8s����S�Y��FP�A���new F�9�|���jl�	��	zR���|���4��e@[��Ӡ��>+��{��'Z\ϕ鴟��&)z�] ggt	ə�:3@ӝ@ۏ�q���AIN�l���.uT3t��{>�g��E�<b�*��M���\b8éI�cݤD�תza7��>�oZ���=پǅ�b�G�W�%/�ҙ�>$pS����_v����2�{9��~g�A)��R�ğ^=G|�J���S�ȫ8]\�k�T
F��4D�r�s{Ҷ}��Ϫ�����E��kv�)�YG?�˱���B���Tb�`BQ��Ԝ�E�Twu���wKӰ�+F9^I�ب+��N̺>�U�|�$��>�*T�=��wlΓ�<��R&��('-a�3�^]�s�/T�s�<��M�C1�3$�D��E�$�8ƺQո΢��o��7f��D-�����H�n�3̖�)R�$�)|�����w�8=��H�oq�k��G���
Y����-�Í$�m3ɶ�����%����H��)|<�y�A�ᛍ"f��9'�����4���(^�aAh�F�UD (U�xve|$=#�01;Æ!]�F%��z����&�{�HZ�n�R��aRrN��bc�� ��9B/�!P^hd��]g,{�2ʘGx���>�[6_td5�pm��yA�E�}��A�w�$�>c�G���O��n�gY�哀�̖�Vρ�*1A�p�5�o5��5+AZ# �a�,GW�?�x��4��Wli�Jo��M�6��$H��Qgḱ�xi�U�����t�J54ZI��>y�:�0� o׎� +ȳ<2T��l��j?�]���O�JF1Ź-blz��7� ��	D���$0v��.#A9;��r���똌Uu/.N`����<LT�`�����;���X����x�vz���I��t.-��_��^\��|���v��Q���g+:�����bs��)��	ʱo(	M�!6�4�j�̍����^_@B��}�L��e�m��Zs/P��6�EI��[�]Nt)��	4�r�����M�Ͱ�������
����A�Xn��t�Z���N��iwe+`�DX�h	@����etǶR�NCCҁ������l3!�������ޓ'Q����"!�0�K"scg�G�OX�JX�##��q����?��H��������y�z�FNn�SH�_S���)�6��孢�*}v����qR�T#j:q߈��*�lVD�O���ݱ�E�D-hP�`���T�&y�FLH�Y|7Q�dqͱ����4NЈ��0���Dx ���϶�/�>v���i֫�%
bN�FdnM���O�� ��hM�fo!;�ug�^u�a#������^i'�m����0��K�?��� ���\��fj�~)�Z��_�q��l�*'����;Ϫ�&�����G�,��!�)]{E�ƹ��J ��)���u�Cʠg��;>=�䧷������
�K��*�k��̤/8���7��^�;*����/O�f�Y���h�>T��e��*_~���:R{�\ɸC�U��������У�6F�q�ҿ�V𺈌��HY�Lͺ��]�����z']{�+���8H�	Nq3��8�
V#{qY��E��kej1h������v�l}�LT?�? �q�̚�_�3�T�O	��ؔrР�^�k���b魤>��ӿ�b,������X�vx���!�#�.k�(�#n0g�3뛫�y�qN~Ơc+��,�C��/�E4b�TEP��yT=N���G����V>�R�Mی�.�躿Q��0��B�{*���D+$�&X'1�ĚRX��Kp;����ߚ��	5�'Y�1fb�z�3�7�����d�i��y��������%�`�8�<8�Z�MX}�؊<m�`<�$pp�D��4����/�_W�|��>�	c�.$��9����@F��A9�A�
^�`b�������g����l.AG��p�BI����>�֓
���/y��:>-������e5��]���!�����>��]/�I0���Fv�EɁC�۾��1g;5���}�9��[k�|�VA��SY�o��T��`L�z�v�<��PO�,��0��`ι!KȆ/���r��EZ�BmZ��}>,#@B�pf�:���fuY�^����L?�L	��yQ��	��-Ac�+X�V�ˮ�EȥtF�ޒ-b���'��XZ��0f{$�o��gCV����6
���
va�/4o��J�6�<w���t�b/�2�[��P�M`�7$f��6up��퇐��bčy]�f~~1��L<�}��d/�.��BF���Wޗ(�?v��/���x�������Ԝ��N�Ss����t�mT�^��y;"�{%x�ÿ"�*����K�Q��M@U��Vi�[�m��ߺ;��";�+�q\�K�9:n�f�x�T��c\w�����$+��ontO�� ��;�\P���ض]�FZ�y6��Fo9���#�,~�����)"�df@������.�=G�6onS����}�����l~����a�Z�{�
���R�V��	���fqN�����G�4(�\����;	#C��h�7��U�~U���X�ا�8�Fڴ]�9%���R�4|��)#t�jG��
�=���q	��Bf���}��N&�u�t�(�*�_
<�#�Cy-��
C�� 똔!����Gq2�{�8CR��٨����O�wʣr䨾$� ��9�Ѕe�_w���6�V�(>~���O���Ü��v��g�M�������G��ڛ�~���df]�3�y�N�������[w�т(C�Q2ϟ���SJ �K��Î�i}n��I�_�D��$���+�b�N�9@!օ����dkLQ5�(��#	��KC���;�>Fo/YE�RW0g՜dB�ηtم:bN���G��mJ?\�73���kކ�E"H����G�_��Oۑ��WnV�n������P��g����H]PL��� /~�h�K����t��;��H�y���?+8v0#~��ʥOx۠��}C�Q���1둦��c�:�\�!ĝFNL�61�s7��$J���~����SP��×11�XV�e��*g\ɫEz�(@O��̤OB~~$�Sn���'��"53�Pa��,����X
��#𠕏��d��4�!ù�H�)'������������:�$��5��`-������Ս