��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]�������|iW��WJ5��`�����"�x�� X��Ȑ�)2�F�Mߛ���8w���ӵ	dQ��y0���Jea۾z�M�@�vyJ̞�O� ��&��Hg�Н�����$9y��������e�9p��+�B[�heBwM�r��������b���t�#}���m�[0=�'��ղ���k�>7l<�t�����3���eP�l/n1�C�Ic�z.�kĤ���Uf�:=��FRN����S;ŧ���i:���Mh�b8i���db�V˺�Q��?ҵ��	Z(mr�U[�)�B��L�/��z�K=R�(߅3�h�������w���q[�����^ޓ2I�6}��^9=���Bk
�O���rl��;�U&H�2w� �#j�8@��Jg0k�tD|��\8$"	2��F\��h�u��T0`/.���)a�qb��ԏ$�]�Ǡq1T�:Q�E #�V��Ά�{����@v8��[c��d0�U��^�Ce]t�@���\���!��UHϊ��,pT�\cp��~��	����,>�iɷ���$sW�m���ڸ����l�nf��R�R� =��V�pǿ�^U�����_*�q��}O�eT��I-:;��r/��Syٱ��,_���q`���sô���F�,^;͞8~yѪ���;��g%������͢�vt-�x0bS�|��m$��I1�ǂ�,CMf/j'0[;��c�R��Ae7��N�,�T���l�0PT�7NB����1�>$�v��"!8~a��j�%c��� �\Þ]�:M�T�E����AxV؈�ڋ��~D����!,G�=���J�hl<P	�V�DF��K�QS33���4�P��_��;�!+1�*uk��P��y�2c����v7Q7=��Jsj�@��ake��<״Bmv��ԷS�|V���.�9�}�({�k.�1�ǽ���d�؃-�p���N��.K����Y���
��{m[L�h��]^�!0n֨���~gz�����>NWW��e�����s�my,�@��;^#�7�j��߅[E^�S�,�o(����=7s���A��˞��BI�3g���t��Rl{��1��p����x��)�b�(�����NgH�:�����vC�b���*����3�]v�����������o"�Lݲ�ql�x�8�E��n���ܻ�)��p�U����(��X4l{�N����}�K[�M���W�ܨ$GX�W�O��̀���XFN�����(�Ψ�̝�MZ�$��`[ k�u���
l#�b��]���q��.�g�R�]."����L��)�y��h�!�#���鐃�FqY}�-���_�\�ǈa�.�ƨ}V		l!���U�D�Jً�D���"��,֣g������ ���b��\S�{ǒ$:x��@T�#��cR��l��~����Wl�3M=͌�}�#���+��k�:�x�"���ֻׅ�Z4cN+Ԁݳ y�����Дk����W	��9^���H�Z�A���~c"�$Po� �$d�Y��[��[1��)d��"����P[�F�����Dg��q.��Q|v�ߦ��)͛ U��o��EC�%�.�)��<��L�aq����< f6��p�;S�G(�ׄ2����t����͍ӿu+U|Yh^I�!���,�^������N���aV��.q1:	�i�v]2���ߖ�$�u�L�O�!Cq9�mZĆ�;��@��-d3碚�M�@����}���'7��C�耽ƞ��j��?*� �`�H�h	�ն$�5�7@bkU��H�7��C�.�r��l��_��0�O[�;x�X�&��H��'z�:�3b����8ؖ�� m����_���9�k�Fŝ1�ڬ=&آ-�,}T?����j�JG����Gh�C��}	�R�<�'�\��I�	/NPjAP�閨`�*�床Q-�p�����7X�/�'�}�v���7�V��'�QY��RY�W�GW��a�LR9C�o{ʅZ]B(ڢs�5�~��
e��)i;��Wn.���U�wt;*_RAd"� ;�0�x�k�>�r�Ҿ�h��w�Q6c��o��e|є	4�����B^�J�Z���ԍ��0�rɬL�N��"ۀϰ$E��P2Ǭ�P�]�lї�|QРy��!�����Т�ol
|B��#=B����rK�)`�"�B�ۑw%Q�����E��5۟1�c��Ȭ��g�9�;��p�诶�r��<)�b�u��/#0~� L7�!��뒑W��y�1����K��ӷK�����jx��	�ѭ�x��fD�y���82�����$�	��.9/`��w�s%����aDE��Ȓ��S��&a`��q�mP�Z=DCmrs�w���U��֚�I:x�\i4)<�[,���=s0,K�h:�O�n��5�P����v�*��`k.R��"��ĳOPl_���ĸ�C���-�	<[ΛH��R��,�����T�|�g	y/���n����.����L���c�*�D��r;�ĭ��*�<��G���[��m���+��/Er���e�Ȁ{s1J$aQK�,A�%�U�v�i������o���!|�l:P[o7���/����(X���$�OՎ��C�G���w��M��;�z�!Rsrs���&<�8�S㼤�^G|�^Q=��|�m��$$< �On�N1���n�e8I#�9G6��7 ߩ����\�r�3�m�l�����ؼA0��`.�<tf�I�^�)�t'���X���ؠ�RSM�eY���y:UV��	��B˖�t1����7!`6`샃��ʢS��ts��cHV<��s��S&����-�L� ��m��3Ƕ��O]���H��K2��Y+�̰ ��L�uF��5�:\V؍<J�͇�!��Ԥ;?߉]�:�i�D������8�ZL�&���D��ѵ�Esn�e�_��v͋u��͹�����skg��DѦ�s %AW�%�pçX�b�R�p�N~���q���������U��4���e����L���.|���3��*L�A��N߿���N�<�S���҆�#�������ϏZ~K�Um�����X���&�ǁ�j��[[��z���PL��i-8Yw���#D��=�<��_Sc� ��6���_Wk�
�T �r���]xm՛�M7b
����-�t���d�T�35�sw �rL?p��`0/������*��ոR0�1U�&=NV�{Bc����.?�U����dbB<�z���9���-��j?�{2�^�ţ�]ao$O�NE�!�8s���w�J��]��y�ͨ��_���ha�r[�f������N�K1���Ȝ$�'�tw�O�(}�M����;�5!!�{�jĂOn4#(����ו�X^l�����\B�F� q���Twɡ�>C��&�CE�Ugt;��a�M��
�k��hf���Pk��)oZv��fO�MR2+�vֈ���0��l�5�%�g$co�!u�-�`p��f٧�;�YCÕ��Q-�����	/D�(ÿ��鉪�����vOi��-�����<�jnߦQ�o�E4w�^=�