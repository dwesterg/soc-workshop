��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��P6��%ܕɒ����[�Z!Jt�oZ�)���C>��G--ƄV�H�4 ��
 � )���o�X��[rLo� �G:����� ]��N����`�k3O4H]�}ݔ�<��dV|��+}���&��F��Pa�[�FstH�8 �Qi1r����fd�E�,�C�bi��ȃ{D ��y��5Y2��A�xs3�I<L9	�(�`�B�#��	��w��#�zE��Z@�kh�� ���o�	M�2���|���#�G6ש�����_�����J���g�⧼�V�V[� � ���A���x�"Ix��}ݤ礹�����BS�W��
A�IE�Dn�*�^�{��+3�@��|��,�����|��v�ZDI��o�,�T�h�C�Ja�K��k'��/d���s���@���ǿ�Ŷ�
�C@��HÈ&t�V�)��Ly?����7��erlbh���ɫX�>����1L��i�f���m�I&DJ��Y]Ө�s��=�M,�EIo�;/j��b� ���A��$Sb�j���I2�d'�x��,#^�9@mO�)�����EZfP�8�-�y�з4}.�r��8��	ZܻW���-�;�ǘ�((��-~1���N�Ip�ߕ����U�߮��Ç�"^�bc�eZ2L"(� !��0�E8q�e�#+��D���&��fT�����5�b�5k��#�֚�CZ�)�=в�
�\��xť1��$xH	�@�nS�4I� �X�1ז`)8���^n�	ݜ~�s��c����~�ͮt ��bz:�w�tYF \�ɷ�,n��㲝�X���Hm�g������v�;R��?�u,~�`����n��t��4��.�>+�gd�8�����m�4�	+ګ�IF}����!��#'�xM��P5&T �e#6׀���aL9Jh��Q/�$wSԯʻ���0��u9�V-�O��6lJpI���׷N��tTŢ���g
4Lݣ��������`Q�٪B���Ɯ�ek��Ir:A6\���\�1��^��G�A���Ed4���UNj*A� TW�8��h3��*Ԇ���c0�|�dg�h����L���8gs,��qlC� B�ɭ"�w�x|f ��%�M��$iDf;ek�󙋽\��l���W�9du�h�U%�+��ulK^�>���vZ����:6�I�41��B�pa���q+�S�E�
�b���˥r�N �*�w^�s�����}8
�f�Ek��T@n�y���t`8���!;��.$T�ڪT�&7�����R5��Pqp�8�
�nd��e��%d}MVP�4�\