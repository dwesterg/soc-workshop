��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ�Bq���F����9��	X�\|(�-��:j��ۏ�,���$��,�Y
��c��9r�?�1���\G��L�T���|Q�CN�0���cJ�H.��3`�H�:sz�+�+�:	r9r+AY�[����9'�|�]�wy�WX6>���S��:O�0��fӭ��ҍ֞���gUbo�����`"�jyᛁ����Qy�J�k� a�q^���;��u|���܃Dq�� t��֨P�����<w?%X��̮T�\��i�n#�3̓g�`DcP��J�*M�*R̺	�+',C#�ڎ�>Pm����gE�Zқ84ud��Z��LmQ_+�f��sW��|�7��rX�\J�'q���v)-�0�t��Z|~3����~$���}����,�\IW'����X`��#�l�bJ�h�U�MͽӟVӎ6�Jg\��y���3��`t5w��?.�����~�Q�D�Oϭ�x�fZ;{��ǔ�J�	���;e�e����e���X���m�p�H�<�-�OBo)�<�P�X�m��ט��}�ƃ�V� ���k{������:΍�Ɗv`_�pQ���?K�z9�\��N�����p�_R��F��X�>DZ���B�{�7<ȁ�F��L�=��QI����e/mf�sW؊�H�s����4�#7��}V�w���,�x�#�ꅤ7�����0�7k+�~�O�8�Ry̶�C���M��kd��E��1�'�E/K|Μ�Ty������U�$�߉��LO#U�y�s�qdg�r�Ȫj�q|F2O��y�3kHo$\QЋe�t�D�F���%��.��>x;��F��F1mDڗ�f��Ma�O�_���P�M#�����3͉�I�P�������ݪADv�?�jԤ�͝��7���!Na(��u9�68$�����\�q �f8�YZ��3Մ��|7͌H�()���©(�?�������qW��bա���Iަ���c1&�oSKj_������Vy�b���]����ĬY�Ə�B�����FG�~�!�pJ)i�^ė��=;���m�ۂ�NV�Wʷ�z���=l����5q�E2��.N�����[�/o9��Sm�� 2S� ��I�+�U1e�NL�k��� )�:S���5�v)�dFs�9��[!+��ѱ���ؘx*i�%�
�l��hHmu-y]�tO��P�9$��|�͒�\5zuG~����7��P�`�v=p����nҏ�"�`���J����<���HDk�ޗ��<��mΞ8��_��}�bw`��A���*�b���o��g�u(�?3�U�װ�����+܇Y��l3c�n��L���jR����aI{�4�߭5��l3���;
\Dp� v{ۍ~�ٸ�L^K>�0�5+L����x�gn�1a��0i�O��=��K8⇆nG�����v`A��L�C:[�^����ID%d���J�i��������@Mx�H��ۮ������"B�./�I�[��
�{&&�J�U*�������t����(f�z�Wwt#�\��9���Rb�B������䁡����.օq3p�»T�n7���?`�s�ȷ\V�oO�����
Q��f��fr����a��a,ￗ_�G�+�{ՇI�-Z��cr�p�+�����,�n�Z�>G��0>�b��,�C��`)[�I)�q&w��fNx;�󸬠@��JOY���U@�x��a�s��f�G�R>��d��2|Ҥp�}-��+��HTC�Q�#�;�t�bk �o,�(HO2��b�_��ն�*�D�I8|da;���}��3���@y�����H�)�:� ��3�hv-��)�j0K1ptLhPXABL���n)5^L)�m��2"�!$"�YC�`ѧ�1�B���o-?,ı�Q,D9����yH �D���DK#�Ń�x9L�(�V}��*WpÆ�����Ӛc6��
�P�(O2�݋�Gu{��a0�����,�]��g��}�-8
v�_Z�u�����MjL��n��|�n��:�D���%�ųA���p���y�ㅐ�����D�a��ڷZ+p��s)Z+����֋���^r�d5)(N9�?�����#���:N������t����x��lݩ�I��m�O�2wK/EL'�Hc����O���� ��K��H�'2���u�dɘ�G�y5O;)��n72�� ��U�_q�S.�u�$9GUo^T�$�����[A�&~V.{u	�k/k��;-�Q�X�pLm8�<k�����^-5�E�A_u,1�i�5@3��>z:WH�,�5u+Ns�N�l.aE3��\���E��Hi�\X�ד��u��m��K��ŶO
�&����%o��aY�x입v�
Ub~E�>R+�γF�
Z��+���^�'�TM���_�i�tC���z�1��޽�a���b�*�*R42�Sj5���?v�V�r�sFDx[z�R�J���[���\gu�c��`�u��x��m0:AΗ�������,l�,��A&H|�Z*n��q�2�؞���yו�7��.GKސ
v�d��Zl4&�AⒾlbS]l�Pa�
�,G�'����k`G��-fmRgD0�ȑG�C�ZXP�Ǟ� +f7�S"�ϋ�r[4XD�%�d#�޷x N��ۯ�Yr�Ӄ �f��Fk���t�@���K9�������񻜤k
���b��DTs����~�M�������UFFZKpԾt��q��V]_��H�7�W�Z6x��'�J��maO�)�m@ j"GW\3�7]]cpU���o.θ��О�LP�R�$I�:W�ѩ��MO���6�u�Q��ں�# H�O>H�+����O}���v�Q�@�P)��;�w �1�x�>c��]E�􇎘k�Զ^H��A�#��VM�?RTڡ��j�F��E�����b[<�-�]ht��)z^-�y'LY��\� ���՚�]��Gg��9z���`��I��lf�oE/gv]:����\�׍�TX����&"m��g�jթ�1���n�#��C
J�ʫ=/�d^��B�@�n�yX�_ln��N{/}�FI�4�Ԧ��O��
2߇��0��\�����]�߄}.Ϭv�����44���k�����M��n<򅱛t�ķOT9�lG-�xj�Sf�	�D\�z_�W��^���;��j��r�!Af <�7���!�hT������޼R�����ra˭�[�����*9ڤ�3�!,��~��h|Y���.x�z��E+s C$16~[�Y�{�"�H��;(n>+��G�V��4���K�\p-���$�d����_Q2�"����./t�Z�c�j)����ɶ'�gE�E@\�㊼�����ۭ.��3�)�L�V�(j`'�u�b���Z[��驢9 ��$���?ަ�]b�^{-�	�|ù"?��&�ѐ��⯰	E~���o�Oq�Ӓ*�~bG6�R.�9fR];�j�� >��i��]�|k���{�L�&=<�DS���V��9Cp�Œ1��M����%���{6ӱ�˂�?(U�aAm�k�Ik��+g���Q6�C�=�vH����C2��[|���f�y���`3��_�,тK<i�7�Dy�:J��1 ���kѺ{�U����bh|���M�%�DO�L�$�M��N$�8FRn�x a"�Hqy�[�H����������N�����S�j2��S����nm�zH������%I��6T1;Y�2���W�����ϲ ���C!.އ�	d�Θ��+��>�Ĭl�q��!���'�{�a��M��kJR#=��J�U0	�v(f�(a��$�{�<�(3� K޼;G��1v�񢄱@3b��4sG0����@�X:sQ �_f��E�ǫ���!�$~�u�sy|ǌ����N�]ͬ����?���
'�퓠�J���9_���	·��T��}�D��׵�wo��%���0oZ�|i���"�^��*��R����&�
[�S�t.�H��a��x��=�Hu8�.ۉ�,ݧQ��,t˩�f����ag��z)�>�dU�GM��_�������;B٨���z�%�D������[g����G��g�����1��K������bS��V�Sq�{]?���\�@Afz�����ώP!�K�.��	����}M��m@�_��:��~-Hdn"��%��2����t�ۙ6�De_�\C�m�|`�~0D�^!�N�҃9�m��= ^v ƁQ��d�]uÐ� v:�3���٢�4s��0,g/��TeC��n
�q�	B�.���]�ޮh�lB䈀�-v����.���(cE4s]r���G�`G�i�
o��_1�����&o$cQC����`��$��2yֹ�-�}��L���%�LV�D4w>��8= ���	Kc���uhk��] ��}:%%fip�0�㖗���Ã�_{��n>I������RY����m��|�F��y1��*�2�rS4�q Z��h�TҼZJ�o8�g�Ftj��ء�EE�\�Ax��o4��'J�1�l��J�%^O���6~�3��O\���\	� 苷&��$��w�~>k��SuE�|�Ǎ3�8�'?�,��@�~ߊ�(��T�]�}�A�ak��6F�R~��)}r�g_y(�|�
B�y����R�����0�y�̞O!w���f����u:���e�@}���]��l�M�k?�/E�����2��J1L�$��5�|��4W�W��F�Ù��G��+�A����h����5p2�f�K?�D�öt���;*����| �����&�H�ktH���,/�7���^$� sb�;k�]�I�8Rz�R��.�"ᔈe��\$zD�i�&2�RPF�}5�z �k��JwN��X� �ݐ�����:������(�2.�L ����є�I*��:|���m����'j�8)
~�����A�����%Z\�0����׵ɲ��%k s�ylU�l���� �̳0!CyAu3�IBFk8�Nd�P�/H��u��hgO-!Aj�C�Ë�,�X?�E�_!�m�ŐRו��E]�aG�19��6J��{.��Ulֽ�Y)�-�i���
�O87Ҭ�;E�oC�p9�2s� d6\M�PUnwI�:��To'���8�r�$��^��\ ʐ��IgF�t	Ķ��<�.z�cd�hW�%���8ƕ1��?���Y0�W'�#�ik��eP���;5�`F3�����Ѷ�H���x���ΣSD�ȑt��UR(&��
b�l����dŢ��[�>>�6%^W�4�f��bo����G��;z;U���!p�+N!��Xi��!�axjZ�瑑�~�6��2&l�L��B�9��(��&��̴�'"�!λ����e'���,;�^fë4_��܇�d1X�eˋ�4�9�)��	�4�.	qgt�����Ӈ_��ke�=��+��k@]i��R9�Of�/6aϯ��5�@���#IpQ��@&�Y��s�!�����T'���܅����ogx�^�tG�[�g��f���c�z��@(fp�r�38U�Я�V�GVYB"��ElE��?�ȪfUi7ux�!�++��V��W��	�l&VX�	�ƽR����yI��]��F����D���£�To������!�a���÷Z�� O�y��N�/���'�!�ˑ�Bg::�@�n�bn��%:U����;j���fV#l��9����BcW+(��K*���TE"�l.���s\T��X�)'i̏�Ѿ���w����M[�ι6�Hrp��]��d��z#��qx���[���&��n:[�ɂ�/�����`EPV�2���U0��t�j;b�M�`�y�̑E��J]�h��������LW"��qf�k���ZO!�N�7��}�^��w.��u���U��b����&$���U `��>�
w��q�9��>Y���H�J�����@��P�g��_KJ�^��*���nes�RM��v9k��E#��ؙ U_T���lϥ�� �5�᱖��7Z�o���AU��{�f��;�~ ��,��0�/���~�`^ʌ�a�]_wb�C��F���	�N8�	����� ڭ<�%!����b�T���G����?`I����֘�#��C�X�u������g)`�w��2b;�y��KA-��s�xu��v9�SŨ|O�S�>&�h�����٫J����2{c'�I���4��H���7E�)}HO���L%��p����6��(Qx���'
F;�H/��o6�@&bH���кK��|� ����3���e)/vf	QWz>�=m��j�6<��I�3/�+Q��.<�L�~My�.��b��&�������/iD��Ot�[݊�	bTԴ�9��X��4ms���{i����4��h�=ɜk�t ����k2�z!�AF�D	��\��.�� C�{WĨ�9r�w�S/�ۋu�%J�)"���G�H��5d��m�L�����C# �������玶οC$(��������RN��"���	h�;�ץ�iV,Q��h�ʴQ��B^���l�{�M�E(j�b��V[ĉ= r,5^�L!¦5}�ԍ{f��Z��SĒԵ�D��@aG�/�6��bQ�s�E�u)7�&� �!¢mu�,i�<��Z����|qk	:����E�ȟ��_�^��4ՙ�����p�:��(�3�E���9g���l�\$�B�#��f�6(��E�I/��_(v�O��;7g5�+��+����;VP[�
��W�R�mմ���25�X��m=K����hi��1�q*^~? �÷I�=F����DKD�T�Y�!aq3S?��v���Ya� �OT���SXs|�l���f��|����GP�N���G��G�!�&~��P��W�F�[�tn�ޤg�.��q�mu�{��/Q��(�,�ga��9����ԗ;� A�2�  %cկ�R�O�V��Z��� ��Ie:�]_-c�� 8���@sV�GT�K�6�a�,+nC#T��Z�ˑ_�h�i������J4DS�|�qk�e�^�$�OxMț�(JAŷ+��Eg�YSْu*���U2�����i���W1-��U�;���}>"��H�ғ���g�VeT���ZfA�->'�`?���(ҌA�1��b�Кǃܟ]xM9���o�y��&��_����D��� V�ǄD�����j�a��U�v���`SK�o-I?s�]~l�!�x���ͬ��{ܤ���w������+��P�.�H�YQ�鶽T:�&
8.1g�Ḥ�IL��P�qL-�\5��?�OA~��=�C���Yy�GX�m������/&�~a�3h�ܲ�����3��NBk���AĈ���Z ��iC�E�=�{QP\��k���|xY��L��X"�\��C��7�]ߋJP
[f:e0_��kc?=���9e[�n�h�ؠMb��:����]O9�#c�awxB��8�������e6�vsb e"�5����̈́Xi�+�T���]�m7�Іֲ����L��8i��K�tGa�C��V�~C�|�f�B�����e�}��Aj�m�jv�n� +40�����55�Rd�ɟ���EנVn�H��^v`�٭�VU=~��H�^}�9��}K��XGN�\�P��ٔʷD�6���$�m�o�i6��Z�Ѭ}��Wks��T�E%Rzݦf��f�Q-���9~��%+EG�?>��h�(��NșA?�hT4o��T�[�1��۬!M]{������8O��j��+gv��nH�� b	���+�&�Z�T�,���QE��� tma�1��)HJp�N��Zx��\2�h*@�1�d�{��*[<Ӯ���=�"�x�!m,�I2�+����Q��� k��S1��所��`:���8r"WG�)�H���#�UF.a�������B)�S-�k��/��r�9�dh|�|��a�d��-�6j������U���m0N�� �^g�@���w�W�^�k�Ьٟ��J��܌�$�0c���m߿�0��p�^&��c�^��ZN&�n^���$ �Z���Q:�NW������$���H`ž�!S�Ϛ�W�)N j3S,@�~��IP�T
���SI�KYLQ��R���M�Yq��>��wuh�{����C*Q�0���	���)m)Py$,��7�W��4)]�;Ǎ�u�W�^��/�ϨA��D��B�1x��D����I�%&O�� ����}�����?woDIB����٥rjIv���	e.��1�2�TQ�5*�~D6{:��e�����1��U��=}�'�~���י�D�W�gsr���PW!Q�|o/�%7��w�R�s�Y^�7 c���� ���f��y'X��阑�ti1𻑡��%a�$Bky׏�B��/~"��!�ۻ �UX_� ���[�W	6�	.Mv �䶂�1���qK�
�{���X*ء�?Q��.<_ee;��*F���p�H�eei��0ݰ�>�c�ĥ�N��#�aAY�x�8�@�`�n�3!��H����YC���,9g�B��/$M��;*w<���׭/V&T�rj �kv�1���y��8ѽ���<��L_2;���jw'�@�Z�o�Q9F'w�Lf�ҫ\��yh��t�6q��{i������2w�
�u2�ArR�}|�PQtђ�&�*�ŝ�<�R4,j��{8E�b�&NWh�p��Y��/Sp�?