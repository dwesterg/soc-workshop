��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��/E���3Vʅ�����v���p��A�̠m}������"�|7g�f 9�����9y�ކ�������M�罘O�{j[_Qg>�1�89Q��v4ac�ʋ�Ȍ�b\8����W������K����R����s��i�vrr���ܴ�<%5�s'Y�G�ӣ>�$s����
�נ��{�%&����d����m�kB8^9�ҏ��R�nL'qn4N_�����l�C��l����l�J�>�Qv���|V y�e��݇�ъ%�=!; $K�/Q�]w��{�<�r�$fC�=&	��@DKd� ̮wu���#l�>��������jY�Y�y?�FD�U|��͗��7CAO&ϯ�<h�!�s��~�^���n�V�\��.�R��8��s�9�����͸m�W�,��l�C��o��Y��?��C͆<@�VA%Go�����룮{���>� �cH�٠�����r�1ѫf���#W)'����C}v��Nh�,?���ۑ��_+�%p��kF�92�g�W��r%��Z�"��&���(���jr���ń0r�N�6H43�E"}��@̷kF}X@[os���E����Cs03=2�y�x�W�&��/ �A^u�G��l;�7�kB#ȗ�J��ѥ�+�����a�Њ�����[VC��ʱ�ڦ��Xj��i�4�	��7H�ŝ�°E6�����=���c&�z��%_İx@�HE���*CC��]r�)�ixk7ʣ���if����t�U8:Ѻr�*H�F+���0�ñ^rm:jU���0T�߯�y#�����GO��E�Q_�d���3f��c�K�#ޠX�?��-C�H�0P�c�]���4�j>@�=P�鰗���\��K݁T�NH����������/����H6�$f5H~d�jA]������S�.,����掗V����n׋�6�1��j�i[��_��5J�(��2Ù#T�s��i��ĜY/����߻}�{��#�
?�'ϡkC%��bнeP�2+v�����ҵ�v������]{!�v��*D��ܚ��UGo�Ȼ���aR̘�%-��d[4��1�7�̽r�)|��b�a8����b!�tI�3݋|[��s����'pG+{�C1�!��EJ�r/WK�p̏�����_ʧ?�{�������U7'�'�H�N��qW����(.7_@+r�a���(��Ϧ\m�\ 2�)�́��7�f�C���xS�����(*����{�7�;�t��-4o����N���Yޚ��6������,���C�� �WVj����!v����C� (���ƅR>� ���b��h���>\�����Ɩr�܏�UQ��\uΧL��?ɼU-&o�ȵ���u����W_���2,?6���A�"�~�[!�}��@�Ċ;v�T�.�<�24y9���$��nꝑAq*j����az������V��z^�.3��*zN��ۍ�����wWD�=ǎ�'� �`�,Svǅ��,��v�����|
���H�����ՙ���Gh5\g�>t����<Pk�:�H��}����N�P��I}��P��aS%_Q��Lgfi*Cu�0�̸",��l0����a$MBa�譂���o7���=o�� �Ug(�Oy�*�YlG��N�N+��ш.:2���(�U\�K�����?VX=D��t x�`�h|���)��V�s�ŴZou1<�O��SJ��^ݗ[��!u�p�T�̢^KN��\w]�oO���(��M�>�av�#�Pɶ�%9qTGw��e��)�ګڡ
6
�D*Ս�[���0M|!T���V�C1d���(�B%�+J�đ׫|��1.8�*��Y"�D6wh6!ڶ�W��&8�ح�4o?:�쎟p~�孃	//��B����$�Ъ���X���"5
��3�]�UMh����ȡ֙�6���&Ȧ�aOtS�A�������?��
+cC�:w��P���)^F��_�L^��l��1F��dC�3���Ul�7rȺ�v��fe	� ?�f���AV� �~�^Px>�vl7H!8�t���P��'��G���b|n�g5��<�`��sJ�U��@���ԥ����H�`��&��ߡe��%QH�VcE�Y��*Q��#^��Yk�:dO�W�n'n\Z͘ps���7�����A3>�T1 �Eӫ_!�	�P�T�2	%��Î��VR�dFt1��֘>�Lfl�?�wN���>2f��B���t��GTq��Z�pG�V��l_�-V��	�����o��2)1���dي��m�.9�5ǀV{����ii��yf�>Ӊ]�>���&w�!B_h���ErO��샋&�r
E���X��B)4�� ����}��IyuO�0&��o-�"t��t=��"�����.�t�ީ/T�,3�s�}Ф
���E�u�k�F ��댚`ߒ���Z�j� �89����~�+����\C��d���Ki�걅���r��v�����u�Gԟ l�h�;
`S�����J�edد��\�l�U������{��^%BG]4��o��GW��>�1�����v-�o�hyd��g����_�ֆ�ЊZi\5ݿ��&�,�Z��MUϓ�a[�[��'Э��o2�����\�����o�])��T����q�+t)���w-5"��'�>�4m�:�(o@���ơ����'4yW��d�5����a?}v�.{�~���h�J��Q�?�5���K��Y�����>^�莻�l&<Е:00�C��}��X�+����e$1�.�+S��[�[h��a�+E�����a22�_ݴ������X��i&�#�!�tW�g�Ǳ�!*X�F� ,m���z����v�� ������01c���uaf�����5+FNQ��	;�3�n)���D�u����B{r�72�a����z���L{� L;��p��=z�/�b��Ldx$fI"xN��_�q�ƀ���A�����/�G�߆�D(vvaKsB�|"�%�Crd:ΐX�"��ZZ싇�X�yᷭ3D���[�׻_���yߥak� �(33	��&^�D�\7��%e��Q2�[�=b;�E�ߚ�"����N��bJ��imQ�x4��{+�p�;jż�m��k7��S���ٺ�2����\�a��
��?,aS�g���~�4,șP�����-p���&h+5�ś`�/@��zZw�ď�O$G�D����[����K�K�ƫѓK%��a��8�Z��,��i;Q�?�@�e+�m��:�0��Y�rl�g��x�_h� ,Cp�)����(�4T��7 ?>ԋ�=T�l(oٕ���2/�|S�n�{�0�{�z��i��O��W"�)4i�6�L�G%�ޜS��5����F`��-�>�e��AJ��8�IA��7�)��'���>���|0�X�9��$�I����������I˪�a�v϶:?���i:
�����w�3���ճ�ϛ��GJu���}�Q�U��#U0׍����N�2|��H�kmݤe4�¶��׸��@D|5g@��@��/��˔�k�u�R��;��&A��V������a o�D�å�+y�d}�7k�1���f���
Gl{��X�G::8o�k�~�������;�Fb�q#�'|B��>p��gfS0��*����h����l)W�eղ�$k�S(ƃ!�����ŧ�P��z�)��^�=�i�c0���G�/��KQ{D�ףz9����Y;ك��;�ₛॽ�gr�ֻ��A��}�<�,i��-���Ę� ��)�.��!-����g�_B����2NÈ��\W�n���=y�`�$k F��rG�[*9�se��
�ڒFΚw#�E=:4�L!*�ȄRS�ܐ2��T~�H����ؔ��Ic�}f����|~`C����J�)gI�e�7�&Ua��L#�.9	�\�fS0��E�һ�M՗+'CN Up.N��"��(@���.�nم�0c*���DX��=�KLH�q'N���x�٨	��)�1h��B]7�[L"�P��X$%{�,�"9�<�,�S��+�Ӥ���������Oݞ���b�!ֆ�l��]������81pXu��l��Rْ��5�#�3ħ�&`>�t�$�z2����o�E82�\֢�(�V�nox��E?����]����a�OA��rୋ�?�ȎY6nsOF���v�F������@R���} =l(L:�|̩1�_F�a&xT����G?}SF���1.m�,���aj�fAIg<��4?H�B���2�*a�'��Su�!�'��2�X~�o3r��D ��8�,���0].脲M��0�_O�0�eo$����H��U��1�g�V���I��5�V����7�y��R�p�l����0KuB�Ȓ�tLB�bK��	�e7qU�TT�:}& �l��|�37�̬}<�DCph�L�	���tX
M�*@�y�cu2%�j�j��4-=Y�w1󃚑wf�x:���/��/V㨵D�W�V�Țׅ���
/��bE��6 ��@����>��P/Z$�������.@Z<dQ�d���D�D��a��ވ�����bt��$�L��4����c
Y���:�B��R,�"������qa���
Y��@ȊE PK��h��	Y�ŏ�z���gѧBmN �^�H�}�S[�JJ~�v�f��>�E�&Oj9����u6| +ݢ�(Yz&f���uNW��׎�}|�*����)�'T�*��FM�c&/y^�^κJjIf�I)���'�v�EN����`x]����}��\��o ��@w<�L�0��p�e�H�	?�/���S���A~�Z��Y��L�ز�a��(���l��K�8U��Vg��fQ��"�s-��_��^t���1T�P��4��(���v=� �Q�h��3��T%>qk]�ֶ�i��R�ۂ�xV���4�9��7Z��w'ZIL�R	Ͼ��ﮎ^|�>|�-�2�؇��9��
W�:_��UK4�E��i�<�Ȓ�7|@1]r�키ť5���8ʮ�~� ��	��z�u�ӛ!�Q��s�ؗ|���	@H�\�����K�,�[V�nlH�1����q��Ѵ�Ze��F+�#�X@�3�\:1ʕ�~̫�;�.&��<��/~$.=F^����&�P��s:�S�Ok��c�&4;6�c�i���v����1Q+A[T���d�чe^+|ɢe�j��g=\d��K�$+D���b�}�$RȰo�R��ڹ���B��w����08�EJ"���)�ۙKl�{�o��J�~�����Ț�����^����:���9@ ��ny@�l�݈t�jVO��!�Y�����j3`h�m�%A��]����ĥ/�����i��eA�����D2��	øRw�� JCu�Ȁ��ߣ�n����a8f��u!#ř��g��8�AD`�;�>��-�
��Od,`�2L����~�?�kbL7�M��z=��R�xap�?KH+�� ?R
1!�y�p0��O<I3$�/Ղ�AbB���T���0���{��q�i��ko� 2�M�=K���kr��߰���ı]5�6�b�YX�Q;w�{�ޫ�h6+/����w��J�ˍYL,���Z3G��G丄�n-��!c�_�����i~)5r�~5�L�8� 3 �(��ݯ�kʂ]څ[�rb��1c�l�� ԫ�\.�t��I�6��0C���A˭;��e�'��gl��%t0������B��!��x��&DC)�e��:\�.j�]�8G�{���Pd3-�Kg��A��:!O��iKN�rr�����˾��R&+i�v�t����t�7���gL ����Da��<rJ�&�g��Ib0K���XY�#U�n�֓��QE��@�F��_�Z�H&<���b�:4����pG��ʹy�Nր�ܸ�t��M�������2�^�'.��&���oF����lOS���u�/.Ԕ�\�o��F��"�F"��Ԯ٭E�&g19�x�W��/<D:F~�*�1�A����<��h�k��N�Ӄ�lЭQ�a3bD��z2�uL�M �7�'XXՀ1� ���M �c]� �V*�?��RbѨO�{�]��[?��*Rη���T��ɍU1Z�g�m4HKha�gqC� k��v)�	%�0/K6V}^�P۩��7�,XG�^��H�y������R;/�}��ˇ�!Y���-�ka t�o�(Ⱥ�͚���ՐdD"S]b�	s:����;h '!��� `�B�x��|&��M�娒V��!vN�H����!�~D���[�5����b����.�6��_?�����6SU�lԚw�Qw���ќ:?�2|կ��ɷb�]jl��+�*�2��p��a\vw��Þ_��jG{��_���>���VM �B�ƞ$��7EKA��?��@�=eǿ�v�����R�f�@p��r=T�gn�����::�[d����N��z9B��IT5m�D4׬|c$���S�E�m�b��b����6�my����z�0]���M/���)���Ǽnm-�IO��B-�,�����׽��D���[軇?�fM��(���F�;�sk��'�xks���N�f��D��L V�5�'����%�T )�o�נX��5~�Q�4wƑGt���9 d�5�����w����E��[?04c\��(�]������8_����^�D��Gц/uY܀V����b��bn�G�������j� �!�����?�;�@���>$�<������d��_�u��֝��~[Ù	�ʂ�(���xX�@ՌųI��$����1�ڰ��� ����Ӑ�LE� �fJ
Άn����nm�'7�S�2ƃ�>C��*P�ȭr�I���W!c��DB�Lο7������g�3v�Ķ���o�*��:��(a���%��R��[x�R�=�*�X+�F���X�s5� ���Q_����魹��.F��������A�<U��3�l��k����	y2��A4��kj�,����E��ft‚�8f�4�1��*ڹk񊆅Y	��r��l�a����2�Ą�M��7L-�f9���/fIqI�@t�{s��v)	�е������Pd���x��6r�6�&�:����f
��]����BC��7��W:v��7����`�Q̇�'/�<��H̓���7���_Tu|rʑ�!��^	�8�m��dW���H�.��0�D.������v�D�e�TOE
CĲl@3�5�b�(��Ge�ο���y��n�C+��̣Mr?h#f��-�&x�\��ʔ`��c�C�&�h"�f'$��e�xc��XC_�O�ʀ��,n)3��<i߱y��nt@a�5�%�2��٥k���ɯSN�_i�����b �<K���� }�Sd`a����ҾU�Sі�6|�:��D��R1|��&����dDܵ9��=o�Q�Itl�F*l�"!��3z�vB�[h�/����m[w͉'"G����k��h:a���5	zP�V�N��l�=:���<����P�E��ĕ��R�!3Y���?=��k���y��{�7��TN��Kx�_���=W�4�Gq_C��b(��5C��.
�҅e�ql�O7}�Q�.�e#j���_b%<	UpkM	�G\7���D�@���A�<,�5������]����G������T����~ɎmLa�:�C�(��8ߥZ���8�DY��	ۖ�ɜTM�W,@�����	���Sb�E���W��\��"!Ԅ�3X39�����(bc�ZϤ3n.���˅��, ��ψw�0@k��P���!���Kb�[�O�nYA'A`���H���C)9�W����e����ȰO!d�0��}�/�j��Si���(ڒV"~�����98��b�@���P'�v|�e��	zB�����WMKldTȥ�y~��;��(t�����/<��+�B��V��8G��0O/��/Jm��v�/�� ��Bw�<�4�}W�z B�Kpi��G9U�E��w���q�4T��t�$�_UǄ��2������x�����;̞J&EKd����G�K�(0e^#�V[���Y��y�����5�_UR��\���;�����l�M��9@o���YMX�5o��Ku8���x��g����w��h�<wPi�a�=<]r�urq�1�"�\��/��+ÄU��Z��L·紐�J5�q�9�@�5���Gf���G�P�fjeJ͹n�>�w@�y���fY�U���� B �'�-ɾ[m9Z^Qpe�a(�7���,�q�l��ZMQ��1a�'�/6
i�b��߻��H�VO�R��h��[�~4ځ뒕��<������)��z�,���כ+��F�r�|��"\�?f�C!�O�l���Gz6�Z#ti�����:�����Yx�Q����:���́��F��R3���'[�ǟ�"�b��M�u��Ȃ��]�tᛟ�%��1A%f95�+��� b$����kp�3�s*��S��X��8��r��_d]F��r�S?�P��G���D铽Ѷ��S�8j�F$��hּ�ې��(���!�1�vtz�^ѝ�������U�<]��?0�X�d��e�� {�5r~a�?�����u��'��J��S{*� �Ie!$E�kck:�ð��]GKsn�D�S~i�Oӊ��ft|�lfJ�

�����@A�m/dC��%�S�zx�aqէ�;�A���H�/�BCǈ�O�4��Ϋ�� ���^&Sz����J��>+}��*S?��t ���S�mn�s��كwn�W�Q����,�-2�Q���C�IeVB�J���ɱc���P�7�j��ȔЄ8{�w����G�֝Sl�{�hs�B������}w]m�9����l�nxW���H��3�pEf�+G�K�9܀!�|
Rw�����wU�R����oڊu�i��V�#�q<�5ƭ��i �Q�H�ѷk�s�<�	���L:(r�GR3G�C�ݣ��\P/��DGk���J�8�,�r��&>��2|��[V���~����I5C��͗}���{ϊ�����<��f_2$���̪�����#�⧜�4QJh�6KDa��}�Uy��Y�@���ď�yo*�s!\'���U����X>�(�a;(���T2�o�Q���6����X���B��2z%T&  ^؂5(�S ]�^������tS�t�����u��f�,�����fX��.G������ae+{���RH�B�ƛ����$;ᨽ�"�
� z�H0=[� {m���w�A��W�*^o��n����Ӧ��)��u]���0R���D�)sl��!���XΗ��m���J[���i":�����k���
��$�7����£��0��Oo)�1'�������^�Å~Ǒ����Y}�ތ�g�j��G:�2/7- Oa�.�qy��E;wL��1����o~�C�Ry���Ӻ}��% z�p���>�ٳgi��w��fG�KW�a�d.O��bm�aێ���0�g�S��UАQA7V0j�F=ִl#��<M3=�&Ƭ�/�$��.ou�g�P�!���¶����|��������/)\�~���91}:!V�HC6�^#�Kuɽ<!U�2�k+�$�b����wf�T`��'���խ�i���,��-�޽�J2�9q��@���Ni!��>
�M��,���z�YmIj��G��EU�Kx���oe�FCU��H��;<�n�h2E�,B�A>�/�Ư��%y��ֆ����W1'~�FzX?���
��m�ux�h#�żj~ɋ@oFĜ �9w���n�Nm�
��O��5Q�j���2�n�NT
��k���R��@�\܊ ����A�ݶ�N�k@\y̮I���/Ն�gx��Ii+!�I��)�K�$j�����u�6�ք�M�Ǔ70J�n9�|g��,�f.[�mg�8壍���D���A�۱/���剦���S�/�9�A�8"U� !�W��sуg���*�8'�̛\#�h�<VZ�b��x����~)�}��ڐ�# ��x���OD;��;EX#�,���+��Y���r�e92�Yn���
Sl�Ѹ�3
�?�4
��$h��I�0�W�ࣲ9���C=�9�U��4��
d�԰VD��ѴK�95�=K��ܶ����ݯ��GBlo��d�Ӣa��V Íǖ�2(���y~֮;����T0}�X��b����5��v9�����W�w �`S�K]������uFD���!8�Kt��4l�	����=�[�B�ʛ �gx4}__����=z�R6�.ѡ�-6�"^[��z��u�(L�_���o� �*
�vr�Q5r0�	� ���կj�����]sT��7�N�hq6MHmu�(�-� n�1dSN\�V�M0O���p�`G/B8�#�o�\kb���	����J�t���P������>���y��H; �Hf�;�b?(n��Ff�٢��p7/��vV���1V�ZQն&2W}��LŋVQ9�r���l�7�ۀ�l��R�$�Y�R�U�~3�B��)��U����V9���'^����+�L��j�'��Ĭ3�9[K�8�3��?��^�A�X�YZ��EeWX��x�q���b�wf�F{K��-'���T����wl;��n�+���'��
t���V@6
Ph3E��v�K�I��m>Gi5�B��f�Ή�K[9V�#�wxao��L_ۅ��q�v=S���E��g@Aԕ��	��7f�p��E֪�*6����u��V:�Xi<U�xN��,m���^Duָ�:�5�9�&-�,t��\�V�L~�/ޢ09�т3<ݥNQ��z< %>�p(Y�r,�eɤ�H�vu1I_�; ����Gߋ���H�����:I�:Yӌ�8]ԕ~:h����n0�����^=cސ���S|K�O�����d��*�����J��/�L(��zy�0"Y=��xC�{�u����ܫ��k�7���IaE�{�*�*���@��v7��w����X@�m:N�����i	�bM�}��캋Q�
���lڭ7+��c`�jR3fP%��r�,����];�����Rjs�`e�;��Bq�	h�5u�~�5�~l��^܇%I���B�r�Fֹ-n|Z٤��ـ��� Q����s�����F&��rH-xh���޾�8<.̮2�(p�9ʱ��:/�9o�<3�=��`/MJ�`�O�����1�a_$Tzi���I��t�}�Z��51�@a���(]��+>t�MI��؃z�����2t$�6�g��%������Ŭ����9<��U�i�Go�d��_х����M*`'Ј�6��M�[6,Y�iA2P��u�oKPu~�w�=;�#��X�%Kt�q�����	���B�̖t ���{����L����S�Li�YO����Wj�Y\����+��͆p���.nY�����qTVM1ӟ��lm�w���!+a%!V�hQ�V .!'[
y(C�Be��[��d&�]�1*�~��pȋds(�$�+���d��w�����ϴ�