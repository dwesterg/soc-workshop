��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t�� ��R�}�m��|��\��A�ZA1+ ����$�ay��ї�ۇ�k��u�м�ad�r-z����4MnF�t��Q~��w�[���J@�K֊�}#��#�r>[I��0l@E��(���ΰr�ޫ�^[8��*�5QOq*z�]f/���d"�,�W�������2馩�)6v%B�U4Г>���^�$������6��ł�F��u/{�H�ѭ�f8k�������*E	U�$;�B��"��=k�����%vY�vr3V�B���Wz�m)�T�$�*Vj��o;���a�N�Y���\F1o��)�ɧ!���Vb��p=��ul����v�8���"����ge��CXuw{�c�y8	/��P~e��A!��ˮ��g����#�9a[{�"�����S����=���e>��[.�E���� �z0F�KͲ=�7�=�4���4�$�g�ì��f�$]�a.��u؉t�ׄ���.|�KAU�~L�xA�����9���c�Qv���c5�ɞ���H�6\�@����y�=��s�A�B߰�����(Q{'��	9���{Ru��"���iR<zS�qU�Oq���t��=P܄ȼ�2���i[2�.)輯�>(�is�h�3�5X;F��Q�Շ|�і�8�ģ�]n��{dkVz=.�h�i�)�V��Į�vRȁP9o`!vt٥�H�m�j�xͧ%N�J`-9����]�!�3�һ��x�'Gt7x��k�%�|am���2��.�,jf|"�	v�{��i�2��:�m�7��yְ=ї
��f榅Ԋ� ���H니d�Xw�PU<4�m�α�����a�T���Tԅ[>7�s���uh�<N֘lQ_��!T;�^}����r�62gdތ����i01q�v�4J�<PaiLZ��h��d��uTqlџ�G=kK�H��{����tYͪܚ�0�"�⬯Ǌ3��S!�?�����OI�/��]��[�h����[X�y�Z��Y�t�<o^������k��\a��iZ�+&�A�'7���se���|�߁-����됫���yu8��m�ʀ��"�6=��@Q��3j���^�E�V�w{Θ�k*��؞���O9�_$xyjE��S�$%��\<�Za;:���E�@�5�$��h�z�^!|X@U�M�yVxr��2K�37�# zo-�*i�Z@)����7����@I���|���<����j�X�0!z�&%�3V���O��Q�n�p����n<�[h�9F�G)�l��xVn�ƚ�1�lr�u�ٟs�$pM[������"$9��N��In[76���@9܆��:#�t
žu�S;FI1�j0�y`>3W? umggnv�ۼ��h�7#����9�j[��gS�/�	�p���V�;���+�xA����:	�ܮI]S�fb�F���[eȔJ'^]}�b~���d��V�攇k��2t�ʭ�\ҌPת��8�:���:��͞6������l3^@�f2��b�'����$�׃՝�wQT��"���%p+�T.��NM������R��vd���+�qi���ٞpi��9�d�[$���2�  �<�q-�E���z���+8Q�����;�F��l<�7����V���d�_d�Զ��l2A�G{3�G�����ʵ�y�,m����}yQ���[�9�`�@�#��B� f�Y����mпa�*ڵ��	��A���4ڌ�gE�r7.�%|{l�E�"j�z��4��1hc�6�N&.d^�g���O�����t���'L�@�����)x�A+P��5�@����##�~U{�W�ey���)/V���G V�.�R�D�����B��Ȫ�����礟fI$n�Yo�+*2y��
��>�:��9������9���F��_բ���Q
ȑdW���㰾?ϵ]���H-���)C�Iߙ�����F�Z�@I���v�t�%��%�ѐ�+�$R�y���YyE	M�Ze��2&岼�Qw,C�_�6Y������MY�vo� ��B��	�/��������������Ŵ��j{������u)�D;)QS�m�P��s,������)��d:k�G�|�	��6N�W��r� �ݑU�n�n�Q���<�AD�L�2�_5��DeN:���vY���O��8@�y���N�@�oWx�q!H%��"IO�.�o�yt�:3�ub�����҅����$�M	����/�fY͸�x�,�a���V���[�MS�>.>�7�u:��C�V'3)I�6�c�V'�ԳEr�p�T0iŻA�?�u���^��;�H����n�Q:�Jk҈~�A0
C�6K�_\<�8(����`y���^��j�F&��^�P�R�~��Z���9ϒ˔����خ�c�"�pY�����}��Zͽ��7:xTIvA㦷����"7𦎂�ت��fr�l���l�����[h�?9�C
�qO����5�Ɔ���X�o�F"v��G��D�|.����ٍ��X\�ekI\Ef`�=��k�H,�����lc�|��u�.�U��䐵UVJ�S$�ep<U�<������	�zVA{J��^�.O�.T�tFA���	vfi�E>��jO��Y���$�+�J���θp\�HDf��Zh_�Χ�(��*ɤx�*Z��+�����(��^Kxk���*��` ]t�r�iT���P�WP�B�'�͎�=����f�MoBQ^n�!6��H0��Q[�D��7R+hb�@~b܅�$ �M��_bZ�it+
'p���;���y�b����W��0��=E��D�.��9S�Udf
��ί��=>V�J��!NV�X[��SM4"5��T���*jӛ��t���Sc_���Ʃ�����oH�OXB��P��(eg):�� ��D_�P�n$2�8a,�-�<�+r-ϐl�;_�������[WL��
 7�Wc���"A䨃��t��$�#�2ف��r7�/(a}���x������2�w��r�W2�DoNs��xY�G��;o;Z�7T�(�\�i�b�̹�)�⃜n<�{�Zhӳ,���7�D����� ~3���_sX�D~Ɲ�
��/Ah�aW՟�	 �I$e�+^ܰ� �ȱ���#2!!�3��`�����@fF��0/1�	���1@Q_��K�0���A�D��]Iy���T�R�ȁ@��;e�~�d�Hr��_z�r���lԱyئa��%�uf�ɓfiKp���k�j#˧��� dw�_�F�[���}Tc��jXB�U��U��e�,X|$�Հ�������
n�Kt��a���C 6���x�J� >ot.�Կ�� ׺1o�y:h�"�*->�� �8 �2�	x
�ᱤ�x��z	���/p�\���#��i�g�����x���=���H>���$i�g�>̶��A���A�i�}Of�ؼn�i�yj�� �s4�t��a�Pka0k��O`-hln�.�����N��(��=�g�G��T��c� 3��q��(~0�*�1�f�g���R,�¤���L���.b��QMZ?V<�N����	U���:�W��� �܁�Ϛ�����_� ��0�z��t��rUA�\��	sFՀ�W0n�⎘�Z�*ў�G�o�л�R�|(�rh��������f��j{�Z'Kz��̓MHi&���L��ѯ�)��&Ѷa;�6XM��^�Я%V8C��}XE�_���%�+a��\��9Z�zg��֠-��yʖ"�"�BHC}�-΂���U���
��#M��ӿ� �>hZ�?��c�+���%��o]ܸ�� ��9d����0�]+
��.����NJ���j9	�{F�@�è�d(9�	��h5�rr����/nXX)�$4�g��a}=9�� N9��8b���)k��mU?�h�2f�|��wI�ID�`jJ����5����}�.�C�,+���lq�0��/�>ڼ��f![.�>�Q��钇���U $����D}W���������=,��+-Y2��9IY���@B�Hzb��p����8W<fy�Ej�ؖ���4-c�f�d�M�Yȍ>����:��xP��)$��.�q�ا��vp��^'�IkMR�t�6�j�M��q�U8��U��-7�%B�H����P�'4Yb����J�;{�~ط>9�YuiY~E���r�Gn�(/�������z��|(��C[xz�Ka�!�C}ܡ.���I��̣!��]�Ib5	ǈ� �v[�����������.�����7@1HlE���ԡ���>�.n|s5�\v
~4׏vI���
H��A��;�!�m�W�g�	���F?h���R��f0G�E��	�B�;��7����/���L���ϊ6V�{$��~?�W]\i��/��s�s�>q{��5t�;�(�8�Fp�#�zc�����{�{���ʑa�곧�\����B�gf�#!\�����2���癋�e�R�*q0�?]�S'dK� �5.�8�xY�E�S��5��V��<�f�F����z�hU��g `��ʗ;�=R'��h�t��w���ϬG�{�h.��t�`Y��BS���_���|
B�	��u���,~��G��	>�1T�·�F\�������ǔ�� �0C�rt��W�aSp�b%.g�T�ߜ��6���Uq��ch�;M�<���\�d��h"���b�k3�O���@=�P���/M���#��� �y�䘏��9%�T+v��$;7�$�n����2[�1i��وJ��} ��׊�Nd{y����v
�UmcGk����R�l��H�QhD�-N�&b^�E��qY]8�L"�
�@+7�����PL����&� ᣋ���\�8�� JR�3/i�/ί��ΌR��U�r�B�`Bԡ��~�3�y��|��Й#��`�ZEJ^�����SD��+ (8�3g4��>Xhe�<�)]J㌻�4.h�=S��;G2}�y�E+����I���mT�E��_�W��'��\Z�x(���h�OwJ6��m7sXId�ۓٚC�Z wEH������t���+�L9�Ą����h JL��AP%��	s?�p�d9��-���)Bqn��d�_C��O�L�˹k�u�kCodB��>шDa%M��.���7�d�P9C'�}���`S�E�9$��"�@'����>!T�W-�o����#��lR�8�񭙡��SzhQ��3(.��|b���֗���Lk��gK?jDe~z�_m}�$��	3ݮ6��+���4�E��T<2����"�탡�L�Ǽ�J���VUX��Z8!�e�e�c���Z*L!���?;���K,
�K��3`�,�KWfp�J���2�L��t�86�P��l��B/6�.���uL��JC��3
�'�$���P_^ngg��%�M�5N��As ��f��S�Ʀx�=����[J	�br��<��t�1�o���쓁�H��N�ID=���k�x���	�ů?��,�X��Um!?-	(~��A��؈���/��y�7�\�S�\q�.�\|���,gJ*�;CE'f���7c��nNI�����kw�a6Y"g��� ;'���-#�vԚOp��#�zX�!��ʖ�a�9���\P�����-NP�5�����*GqۂH�����%C:8�C�����Y�{fA�7�g!�۴mzh�N�I�K��g�˰u�4]�h����򯺛,Y��k� U.a�ˤ~m!O98_��c_��/����$��w�`��U�Ъ.�qk�@{�a-���Gxa*� 	�,(dW7��&G��u��@n����n�{�(�rˑ����{l%�i�Դ����짫��������E��)4�s�fҪ�F�'�B([��d�d��g����T赕"M���lh���g҂���[P�f�oM���fJ�߁��� 	�q;(aFc�PeU����*)��s�!�8��-�������,�8�]'��\��S�b&ڷ���֩�Cx���T�W�5��_â��6ۧ����5_}���V}�H��(0e�v���@�d˕�[�_��_+8}�-�W{�� �������ȋ�F���61�2�0��!��2U,|vh�Ң4ƪ�O�ڍX^���C���Ҿd���(���X�n�F�M$�,�����/�O�d�i�j1���&>�F�#���k0��[�����h�&Bs��9%�	zd�
���g�����[�;/� ���|VǑm���ЇB�"�Uki����L�Ĉs~]�ڼ��=E_��8
_u"}�V����ٴ�x{�J͚��=%�;���v��]<��5|"O���00�+9��kR�N�ިY�.��z,�����1����XQ}�a�CMHvL_����X�S���C���������O���#ƙ>�0V�H���(b�(5!�c��X'�p�W�AeMS�u�{,GT!� ����U�����i�>���M,�e4��en�o��D�����9>%�����v�[1H�u"U:>^�'EIN���&�ҧ%�}�^A�E������G�S�)�pԽ��2(��>�)�G��0��+�8��T���NSr��<��e�S¥G\i�ŵ/��1�p�u�ŋ��z�������g9����P2=��޳�2���f�;2y���8�vt�laZ��W���C��}!�> ��RN�C~F�-pV4:Y���f�Rk�����O�x��b�>ƶ¾GsPNp��0��&�&����+�yv�1G�z�ih{#,'��pKy*���,�R���@ݽ7��.�r֌Q'�D<��	GJ�������	�w��1Ƀ��_�-u�6�%�z*V"vY��k�DE	 �~�O ��Z@Z+�亂�e��H���<U�y{}���3��C��0���e���`�>��ߘ�c���-o݋�e)��[&L��N;�61��%��̀���S���e޲����l���{�3E�16>B�mN7�v�ת�Ӄ �r�U����v<Л�h}���v�π�ݵ��.WY��݅��c�B�\�BU�{��:�ɳO�H3�3�`b�mF�&z���l�M�iɏ4� x"��(L7/�^T_����c�b��X�d���3M���P<�3�-���0
yQ�t3�O D(�4т6x �'�'�Ӝ��v/����0�c��A���M0�C� J��D��6J�s�j���dJ�p�Q�I=�����]�9�0����]���҆�m��޿>�o�2[�&i����Yr����A�������7Ĭ@���r=�i�qy!�n�+������k�������L��e�,�=
����3;ni{�����JT�f-\8�Oe�M��X ���n?�Ys �:I�Y�l9jQ��ձ
S�Y�b�}yZ�ɑ��I��
�<��='j�۩24.�"i$<��-]��j�OY?�V�"Q�I1�XڍW4��𸁸+^:��'��4T8�5Qf�Ea��+ �w�HK�V�UUaz����e��s-E3���R�ζ��-��i!�"*"q����['B�C���$N��x�罻X�.�..��g$�py��vr�?��ݩF�H��Hj͒*�Ksyԗ^cG���\V��HW�@��b�fa �L/�~}�kL����R�o�ö0��<��q/[׿B�Y&�%����������*?G��pd2��H')~x{\�O���f9��"�z��oZ!B�z�69��8�E�c�A.����{ԴUHT����J.�'d�����'q`ں%�5S2w"�5�M�;�7*cX�Ԏ׳,w��J�,��n�o��[�0s�X*�Z �Xٰ&���ۗ!4ڌ^9T&Ԍ!�ݦ�^�b�.|];���>�U�,���zZ"U��>Gm'�О? �f���`#����u�u������ɳ>N�P��H���0f�\W��3QA0���j�Æ�3x*�uu ��)���Mwޒ]~K�V��1h�Ǣv3�Y%9�m�'�FԆ7��IU�����P�]�ww��L���X,LaP�7E����Hb�S�c�L`��� ��1�������e�n�� �z�����~0B��YbF �X�~WbZ��f�쾰��OΕ>jc��aѳ���[�O��sT�s�����h�%Q�
~z��~�x^�����0}�kZ��3v����E`a|����!e��SQIu���9tN��L	��C5���W���p�Ր���x�Q1G<�}5�U�t�����t���æ���m�*�'�_��^ ���~=�g��3�e�&F�,�OZ8�kϮF-'iʉ��pp�n��I�GD�	� �5j�#�=N�tPV �z}����]I��m(/��x���(z�^��sGm���V�}�:�?��)[�����~�=�!g�j5C����#���K�v����p��d�އ�'���J�-"��9��4Q^��[�9�LV��.���E�͡��Z*/g^��<�)AK?N=}����w��S��E���lv��;��u�E�O��h0or�t�w҅��q���e�G ���~�4,�P*�[����5:�aB�h��������^ypT������I��"#c���ς!]�c��
�3>N�"^{Q���t���܉H�	�z�
�8��dT��x�y?~ų�S������G�n���{����}���ԕ��4�����򆈬+��ɂ���^g��2L��+nhoT�b�.(����/r�,����\|uI�S��� �I��j��UYW�@�䓋"T��e��*�C݊,&�Wm�\H�� �o��_<�49�~���þ�W�c���`���yV��qgj?+�^R����5����c��|���1d���UE0_�P��#��&7^6OM|��W�u�*u�����B9,+�����;�)���
�òe5qq��6��P.��@�0ގ��-�U�`��:S=#�ښ>�k
|d�/�IA���Zk��,b�L�>�>]���xͳ7�+#̳�wG���vM��8u|T��m-�7�S[�l�f@���t���[��O�zcA��s�(���Uqw���ϳ��	��s*Ԩ��.���V��;ʺ�S��IcҬGn_C�T���o-�LJ#
��d!1�r��14}uoQ�q#��A�	��Y�fG���O�x��X3F����k���n勎�@r.�wiV��?kJ��]�����q9т1mEC@Ce� %&�mF|�O�������|i+A���.���k�����W9n?u!�#���ɞ沔��i /sv�������	LD ��c�n��C`�s���]���,��:5�)}sV�ѭE�\Dq|��3
|z�*DnO1iɘ�.�LNC�9z��nɀ�ĢQV�q��q9���4��}�w~�o��3Aus�L������k�L��R�<��	'3k�zKBgK.��p8�����������
Py;ڰ�f��f���Җ��Ģ��󬐯���{�Jk��a�ʲ8�_�+�|
C�B�Uվ������A+��2��XM���E4}�Gu+�Z�a�4m#�������^�d|�r��6�c�>�2����\� ���<6
K����s���L)�k6_a�r��"͞��%��^>>�֛$�hc�U<��k��t���4���a���i�ޭ����	|/���✭��%qP��g9��0�y��K�v��+h��5{>��{���.�\r���)�	<�Ȭaa�L�X��hM���=�%H�j���
|�C�"��S�#���c�s.W͠�i���꣯��mO|�@��e
�L,�B� �*��%��s��FS����Gͧ�����:Zmp�*i��k��ݷ�o8>W��B��f<M=h#a"��b(����c��`-c���0�������O%�z	���
{&��Bm���
�&��/�d�	���셆�i���S�7�ch��~�*���,!����m|��K�Yk7ϲrq�?���r!וv�[Um� |&�>���E��������/l�q�	-u��t�mS7!&~���� /+j��_�2/���v�,A����P�O�$I���K�>��!��3�7�=�d��zi�@�gF����q��&ݔjm�>���Q��#��i/!����s�M�2�V����{�QXt:�佞4�(�$�6f@$ʙ � 3�q����G^��l��ԓA��0��t�?�;�|F�Ǌ��e�K�� ����5`Ƣ�߹@:a	|��L�<�c��ܚ��e���<3mȋ���_�$�oB�ޓ�$�A�k!�/ƿٽA�0��F�qd�	#~0հ��ȦY�D�ƗX��. ��J.wu6�K,Y��������J�3�ΰ���Hwx&�����������VM�E�:��F��8X5�׀�7K�<��j��V���3�\�_��J�h���k�Ep�L�u3�m[S��	�����J3���B�͢ώ d����nc��kj |�?B����=/w����5��|[۫�u��.�"��I�L!�.p�V	��X�Js��;Yty6���洔�+��U��D40���|��_ N����6�,TOD�K���-�[�ZGV`�sh@���,�����3�EsA.%�9�������0��I�],��;�(aW��xP2d0Պwq�����qȗ�T��0�EB���b�9�5R��]�=��}�uL���8$�^�r�s��M�W>��M{v=���>}��_��R-��xV2+'�w�2G'7 �Z3c��� ���g?�-��$O�^�ۧ��*���.��B%
��>�ׁ;�����f�\�Zȼ�}�>bL���3�)6��H���bM�/e�קȂ"�MN����<�jm*��K?�@I�U�6G�}�z��aD�hg�R���Ӄ�!5(v;�p�������-�֝~��&�2D"�A�Q�F!Ň�^�6����?��lB+�Qq7������լ���]ָ�.�����u�v��5r_����7]�q���,�*Y��f~Ӛ��+�t�ZB��"-^�%�	���\ΰLlb����'�<e櫉G4������K���Bi+祐� ���U����w�)c�
&�Ȁ�����A��ҿ�՚�_�5�S����a4����rw�F����Z�ψ \-��q��b�6���h�f��|�!UkÄ�
M�+Qٮ��+w����<V������L+����YDe)�5�9J�,~�ٱ:h��`?/���v|���"\W��2�P�֭�eoI�x�;O=�PczsI��R='���3�I��6fɸƁKI�O[+��w(>O��7qb�t�_�x���(WG�X2�X��P+�_���q��-�~��������_��yF�Ge3u:��
s���]��2�щ7,^`wB�����rj�C�	�򌃏���%��se�`��tz"H��Ǹ�I���r�G��hX3�bYG49����i#�(�DNI#F�x��7��%3��>��^������$�X���ݕeW0n�A�.��W�8���m�ն3�KZ�w��%H=L��/<��G�����D[]b�+�=:��� ��C��>��v��{cY8���2BgY�/������9vDQ*�,Z���<��8�m�����3�v�Ȫ��a���#&8��n=~����t�
APOW�F���!@���4|'�	
"9|H��ghJ
i�u�Y��м��w�=��,�3U���Y���qYWf�?��^�����/��;���:����X܆W?(�/uD8�G!8�%x.��������az�֪�?���P��_%?���N��d=�zV����w)�室���;��P*��IV.�b�J�&��>?(�'ߜ�K�RC��b��zӎzlv�N��,i(�FƇ8�*���F�(�#�߼_�VZX��{^8��-�'�aV=�枎;U�Oz���ʥ�~�K5&�����U_7�]����R�.�_|�a=��R���H�6��t�ݝn�H���i��v���Ĵ`I@�#AjɈ���!����̫{�3/�z)kݫ�0v�I�ˢ�v�mHZ;�����L�3Ȉ��NR���Fc��q4l5�UVD%Œ��(�	����X�Oq��USVz2�8Pl��K�zB���Z���sù�^�d���u��gT�d	��EJ@�2���*L�	7���RU*l��)�w2w��S�ٱ���*���u�� ��Q=��uD��n*WJf���S�"x�Zb`�z�o������;�J��L��L}ʺcX�\�J�|I���L2���Ē�Y�S���Q�v�*O�4���A9��Z�T	�b�������������$�����C�K�����QE�L�ݚ.ܚsB	����^��e�m�:�;�OH�W|�xk}L{7F�8s�w�l�7ow�J�W%��H�� ��&��(Z���wuF�lc�h���T�b3n#&x���;��p��w�礔b��h�	��� X|Ro8u&�P�{��-hO�
���i�yliɧ�#x�9g�D�*�i+ն�J���B|Պ�w�6<���ܦ߫X۽���T@�P��E��7立�TQ[�]�� �t�ן�s�W���z9�Q�z�cX���#ht��-�u��" �M�q��a�h�V9�����r-�qP��k��2��v3Snwp�p�~A�cR0'�������H+�m�c��������MS���2����j� ��r���|X�i�ΎB}ԭ�.V����)t��-z���OrF:t�G(k
4p���h�׋.�<��x,E[o���P}h5���\bp��/2�=ɃH{
�˂�ߪI~V�n�ܧl�,v���ђ'J���r1bw���n�h:\�(�[>�� s�4`t�q�t���!�����X�_"P-������	ؐ[�.pM�'Q��mcM�Y�#��רʹ[5H�e�_������0�ھ��p�(+xn�*"���3C]���+q|߂6��6%������� �3Ň����)])A,���EF�k���-�n��u`���{�:Y�+�,.����p@Z��-Bl|���`7xg�fA^$е���MO�i~H��+���ʹ���잸-wB�$h�C,�rBNN�^����ȇ6�2��+�y? 9�-�.C�MG��L���!�x�O�����e����"r�yU��w�?\l���a-�VYS�KB	��j\�E� �P��@��Z�o�Y�xs�e�C���mH0�O����� ��W��' ����u��V(`�o(5%t��YcѪ2lm����G�⦓�9�Ku-R��ߌ2"B��V]}�������8�GAw����a;�YJ�Z���=U2�����Q2U�V��[t���@�DD<,�ɲ8$Ͳ���ea��a¨�ħw��J�ס�}R�����yŃa�@v�=�Rh�\��L��k�
lp�r9M��t5ъ��S�����g�����Tf���P/�<Ox���4�#�\����P��o)��0kᦏ��ɡ���"Kd���m��ӂJ�x�Y4��ˊ����%���2����u���ƠF�^�X�oXj㱶���D=L����nz
SrxX��J%�=ɥ�߽PS��	1���X �Z8\�7ź�Ӗ�}/��j�v�,�Q)�7�ᫍg�kw�9��!{J?�o)`Dyٳ��t��J  ���u-����1���N�C�m,��(�`�׉ݾ�� �Rӹ�����T��< P��A�e�����R����f)��,�4_;�r��g���	��D����+=B�K'{Kʤ�&����fѦ0F��e�z_�e��uZnP���-
�p.S�]��
IEhӢ��fT����9��\�� *�O)��3&���ǮBE���� �	 �(�
YFFJp1��j��'�fn��C�������#�����k�6�ߥ��f� \i�K�N��\+�c41��;K����Ã
�cJ�n�8����?u���he3qn�s�O=h�i���(~KQ�J��C����k��Usc�^�2�w�Ү�w��S_VTGF�����&x��U��QJ���w�"P �wXFT	�sPɮ�;�$����
����6���æ�C`?$�?�08R/��NoSv�:P�vp���A��h�|~Oj�6gT��a
~���凜X�O���}��a����%27\�Ӽ���RY��x�5Ѯ'�x���h��?�~pY���+<@��ڿ����5kЙ�(i�Rr8�����;> ���*2�����[ ��o��-�"��c:u0��hZ�D������e^��S���I	$�ؿ���pS*O'��x�� �
D�!���r�J��jJ��^Y�:B�
��	G�S�p �[��܍���4��5!gސN���L?�e`S�WJ��"�G2��j��X	M�P�\'i�V0��p���Q��|��`S=4��5��+&b��Q	x~
�w;KH���� �!=�r�}��emfm�jV�?�yc��^�/K��Bڴ���yS��	N�_JN�6߷�8]o�F���	AB̋��{ZNX�d&I����T�M�`9e��=�쭆$�>\��.��>T�Y��3X��[s�0����+�2=��/B��L���{����K��������cZI<X7Ob�Kf����Hr}��/`O)׉�����"���;�,c�p�� �\U�~���Ե�e .6�M^��6�ڶVq�ZN����d<�0�>@�NK��ω*��,��a���H���U�l@p�e�jDǚP�cS�2-,Y�Gr]rTp�T�Lׁ�4���8�?Ft���Å����x+Ȣ� �;{J�O���������]�p�v�<��o����U����.��>a�4�r��93K�k�͵t�A�9��և�BG��c����z��@�,���֑�C^#�9Ab�x�aV �j`�j���FfV�%����_j���A�������~F�)Kъ����2����A[�;�K�P��#��2� j��]���/�!_�5xt�2I�$0(V�ʋ��Ҷ�GP���M(���qm<[�0A�J�|gs&�㫗��B���8�Ap�/=�e���MUd2ޖK�ӓ��_�]�XM;Lq~�F<��Q�?T*��~{V��:á��~ux$�o2巴%R ���q�n!ik]L�5$�I]�&_��ˉP�axS��a�֤4��8���r��>r:�� W��S��a7�i��wC��<u跎��RճuL�g�l�|>��Dk�r�PCr<ܫ�\e��� �s��]1���m�����TPkK�Y�F�H@
�:>�.��}.���Y�}0�m�Ǌ�Ǽ�5x���[9��?`3���Ј�~���-�O������t�Aid��I��ܐB@�_�R3�k�vk�p�Lj�-4���-Jչ}65���^��+t�.q2���� %gE����A�.�E�Z5�����C���i�_�����]�y��˯|�	ś�Nq���e��#&*V5Z\������ڠ�����r]�h���m�[��C���݋�ŝ���>!C�?����R"����簁�j�cnkA�*~Y����J�Yf)�٣sҎ�N짓��|�Q�ڎ�Sȇ�Y'f0q�j�2;u��.g�'������<�m�J>�b��-ݍ!*�*Ut��_����s�2��ߴ
W(�	�:���ZM�P.�D�v����N.~����U<�[5�T-R��tD�^�f���m�z�a;RH>�Sk��9�anW ��9)D��M��}X1U%�.>&P?'�Ԥ.?}l?�:�d�I-��C9�+.������K?�f ^$��q������A���Ţ��U(��Cj/( Qwy�
����(��ijʑ�:bb
A�0$�6f�tY-;�7VC'=��A���D	JJi�A�It"���1�!���8�N��P2uh�~Z��+���9Ee��%�0MD�~Q{W�� �)�(X�s�������iT-y[����R��g�2�PS�t{"�5D�`(��=��!�=�$�hA|��Q	`�-Gkۭ�A�9��>!%�S�H)��&�78#I���+C��֗Խ<������3P ߊ ���lwP�;(.��fs��g��1�����&�ց�{�pw���/&9���&�yv��[�ቡNL�J��d��rë�6��;tˇ`Y/��Q7�0��ꧤ�Ǝ���[v�w����qko�2��`�2s���dlNxJ0����?T�#+;���8��7ч4Rq��VN���N94]D����ว���)R��j\�h��3�T���ϵ�]���"Z�������uEK�D�ڝ@�E^����N��ς �[^��}S�܇�ܸ�|�8	�YߐD5��|���
V��;��&���e���EjS�/ĝ��ʒ��hD�6��+�+e� �}���'�1Bo`#�;�`���26�''�}��G�TG�&Z3ݛ�G�=���m�2����#��@A98t�j��~���/3>��
�Y4�n�,��7$��;�Q;�$�i �yT�q*3m逃��7��/ !%�n]a76����0�rH�Ca��n�  ?���$��=Q��z�a�>� mR��$����{-Lq��T�g��%�i����$O��v�SN�83?t�7(�GͿ���#�j�Z���kQHZ�R[�=X)�{�j�N�wby��u���q�]ԿRQC����_
T9�t�����/����І,^�4�Ógr-�~�{�þ��U�"�S=�y�'�J������	�x8S�@�r�9��}µ��NZs��s�H��՞D@��5+�|�k��[s4���_^�jjwR����6>�,J���)*y��k9�?��61����= ����a�\<6��$���fmuq�r��_�/��ڱS�g��d�I��=dʎeh�{	�$6�MZ3b��B����Ge�Rՙa�z��~O�q5
Ǆ���?�W\���PR
�p�/�0��Z�Ҥ�� X�|Ug��P���D�op��j?o��&���M�G����Hō_f[������
���ER���P,���`\\�p��o5iC�2=��V�u�O�7�^u�r��t[�S�1�l��D�˗�4q������oqg�E�������9��:q@-i�s|��pk�.b`�g���O��V�y#.x�t�[�X��ATq���&�EoaZv�Y�H�,�+s���ݲSU��<đi\[�����$٠Ҷ5�N"<���.~�t->�5��s�f~�S+hN�TZ���^͂��U�d�D�eB̫XL��.h��0��N�x�'���q�;��,�p�A�F:��S �����A��G�g��[zk�;��lS� �R�5����̱N�9ߔ�DF���^��2�.�)�G�2�;Ⱥx���� YW�X��N��F�����$>~�:�$JR�Z$���M�[h�ݣt嘚M��R�\�O�����3ߌ"����E�.�ڴ%�ѻ�>��m�3�Ǐ��3��2����U�}p��F\���ǵ�6�s:��&_�#�x{E(�۪J�xc�@N6�<�$Mp���1B���R��Dl�*Q��B�G�3*�AQn�=|��Rz� (�n�1��x�����#aX��?�ˑpxC��׭,zz��ϒ�?���p��~:N�m�!�6(�Ae�.��1��`���l�$�����/Q×��Dhc�Cy����2�����7�n�{�~(��݂�A3U۴�̈́/�ױ���R��卖U �O0�ޒ�,�m(��O,x'��I��S�~5��X/���^k}�i%�f�b/�؎s�j[`����R�yj�E��N�^�'����! �[^�Q>�RG��+�s_�3Ɂfrނ��G�U�+��Ũ"K��[���
�n��Wȩ�-��勞$��ljsO����)d[ɕ-������PM!�����u�%���� j_�8� ������]�$�Y{u��V,X�ގa�Eh�EVw�Ag��-�}���؇7��L'f�I��M�P��CDb�ѝ��H�$����G���?�-������# ���r�xD����%������xd���q�1C�<O؞������?v�x�$!F���!)��lb�~S|a��UQng>JZ�r�y���x�����qq��U ?nD�u��X����3��p�?CԟoX�����VR��ݖ�F��c��y�l����ō��Z\����+n���>�Q�\8~B7-��2p�T�Y����o8��g�:c?R���
�3ld���R7�:��#�=L�N�)m^{���.(R��[��x.�6��jEr�����(�?cs���٘\�m�K�1�����I#Y��\[�.R/Z=4�<� X�h�R�\��q�
e�[��uNXvˍ�.�	�wp�⁳W�6m��T�n�gL�v��C΃��C�V��+~QuY:�sٶ4)ɥ3�-q;󪳒��Ebƥ�Д������D�k�R ��ŭ��
Z#��-�� 
z�`��z����/��B#�Mw�_�,*�q����9��=!w�u{OP-��}��j�1�˗@��kZƃ�5}�3?�א�H�?|X�ʝ�H�ڑL�*Y&|�
����
ϵ�&a˙�o\pL�zW=YF�9,aŦ�32�Zp�P�du44P�����Am�-f �qG��I�Ay@rV�Y��{��Gِ@)���Ka=�v��玝jI�e���-����V���l��,�
�K8�~�饋E��Lw_�Ha�&[E#�	Ȣ�?����g��ho�/�4��5����;�pǅ#�t/��	�=��ƞ`����1vt ����9�4eKk�̰��.�E��W�]/�@��T�S>7Y`��C�ָ���A���Q��[�j�=�pƣ$ֵ:i����|Yv����:�Ł���xt�<l���0L�g�G�7�+�$.P%�E3(��X�Rva��B��epM��?ķP#-*��4�C&��~��N�!���ɆOƜ���[3 Ǌ�$cP2cN;Fj�s ��<���� :�ҵ���5��7x 9�:��g�V����������]7���[�����?�F`����S,�P�5뇴B8Yqq�+�o���T  ^�R��Z	�Y��'3��5\��Ah������z��������[���z���CqA�]룚l:<���|�y�K�Ҳ�}sN������`��!��/�:�&����}�u�b�#N�Cd����&�D�XU���/xК��O����A^��Ǹ2��Nڛu�u�f1˘�2�y�r��g	�hy�=苟;c(���E^���➁��"�rCoF��y:�
�vic�����-1j�K9�
�]�I��,ɯmh?����J�߸�^��+�-���|>[*�<�0���?O39[����*����y���1�͒@ �M��vXK��~Z�h���wW���؝]P B�r�7�	����.�ܴI3����6"_a�J�`	�2�=ʦ#�����!  ��r�NF\]�m��G�z��r:grę��kg�ō�wM���k��^���e�� �0qz��oȗp�K����W�9�]}P� 86�$�G/y����.1�"@��S��c�O�pJՄ7�.j�`h�s7E{�%���)4U�s-�V�z}+M���gM�;�Klt_�>}"�L�����^��\���Cɤ0�U�?U H���GHhg�u�I�,����Z���5�f��/�5R_A��^L9�@}�;�ɞ���e�<]��[�6Td��~�U�3�R�l2%�}JegUqɸ�G�2�#**���E�	�p�w��;y�g���R��" `���х7}�d�)]o�j~�/5�2@��=���|��Q�R�ffNf���1Y��ϩqPh/3�Z;O!�|mPcR���%��S�`v6Q�u�ذJR.[6|죰@,�5�(z��I��y�~Z��n�>x#y���Z��%sA�b���]�'|�M7Tܬ��6��M6�tJI���-���;-xRu�4�T8].��oL�m	hb�mĦV�4�`B-n"j�	�������W��O{�㏐M&�}	�r(��We,d`�����'
�-�����a����s��TY�Zy_Z���VĤ�����7��W�B��J�v H�ؕMO�����G�(<Jn��6�@:�u���m��{?�df����V�ʯ7p<wU��*ǃ~�y~���
[-*�A�> ����ƙj�n��aUУ����e{%S�����%�̇CP���Z�?_��
0k��ܔ|:�;�Y�yy�ʐ��/rs(7Rz�S+koUQ�S4q��������"�4+_&)��h�*��o�Y�wW_Ɍi���@8��X��>��pٴ|X\Ş
�Ayqj��T̙y��%�F�.���h旳�<Q� �d�h�@�L��X��<#4x2*"i/�@���tz�컬�5���m}�0Qc�=s�ہr�B�-�E�5Man���g( �ivqН��F+��u�G�6��a:�! O��)��{Sx({��1-S�1%ɽ�yΖM����C<�'�Va�PB�wԹ�+�� {h��%	8��a'�V�K`�5�Rp	��]����#��q`;*�r0�$2�C@�%O��8~��k�j>g�0$��y��;�"�������"8��|P��$n�z^uO������A���DR!�3;�wͯ���^�>'&���w���oz�ߍ�Lܺ�/�D���M��é ��@>�m�ٹ�N�����OPq�:|�S�>QM�n��U�&ȏ��%��q�o:�C_�sS�GOz��kh�3	�!0m���>�s��EJ]:�I�O�ң�Qn�$x:G�������Tƪ��n7�M��K	t��r�M�S_��Ly��b��؄s�'�C?�7��h��e�K�ߒ��������(��c�5�.v���!�5���V#�-Ùrܳ�kL��7!��@׹���Ü�����d�b#8<���:�V���'i�ȵ�Z�Ս��5(�Ŭ������ZO#>��%E[�@Ar�
	&pa���j����|h�L�&��-WѬb� _�E<!/�~�ҙ`��� �i�� s_E�*��ů��uL1qJ��d�K��>�S�%�FB9@���Ϳj�&W��نb��N��p�-�5]n"�
	邸��8�`ǧR��o ���� �-Au�xeiR3�B���\Vb�P{��f���T��oi-����VM��t����@����s`q�.���%�n5��$ ������ޜ,<5��!���r3.�8J;�Iy�SC�Ԯ�����"�{m<�'ƌ��9|�'��zR҇5��>�������>&�p�;�RR�f)Ԭ��x-!�T�p�����vV��%��պ]lX������zz"�����xCo���T��2V�#Lm��0����4=�V�i�#C7��3�{XL�u�m�&k��E!r/�1�����v�����n�R��ʆ�n�L��z�YդRxT��%�W�q�V�٥��Cj��	�)�b�v���eF���Rj��\���bB��賚�ܤ�,+Ri-�J��`��h�� ��� �HΏ��#�H]+gu�;9�QL��5�þ���H��šUÄ�u�?F�I�w`_N2�*�KE.S!+ƚ��t� UT�ny%]_�LNW(Ehd��J$l��=��寯�tp��F}#�`0
�3�_MH&���I2�����kqe��}��;aa �e�?9	B��/�����w��'S�t��h�f>�͘]w���r͒38:65g�o���١�J"��8�fu���U� j�.�4g$C�#Oڴ�m#�S�\y�uu���4��V_�0��S�U�����N~s֞����T`H���D~�TE��w17���2�r������ڷ�ƶ~��p����Uc�ķF����8�8�tdÝ��m�Ȗ84b���a�m6B��1���V: _��V�IL�;q	f��>H)���>��F�?�Þ7��l�c܉Ė��S���b�0���N1��B�e�o$
��r�L�S�����KC�������!A�u��%22�=v���U�8�F�`{R��L*�I���ts��И��w�#��bYW�f�	̃A���ߨ���u�-�L�`n��?*N���f�;����{�`�i���c��u�M��LU;!�hL��l*$�	����8q��"IG��Kx��*��d�8��M�e��'������Z��Gd�\�B�=��$rL�M�������Z�3�j��8{(t������vg������q�W
LF��؞̼��{�?ա�ԛ���5��:�F��1�i.�ﱖ�����ْ)4A���`��/E��{�u���s1Ѓ�����=E$Ni�z�垡�z�i����3ech��L�K�y�lr�5Y�Y �j�,{hT�pr�� E���b^���Q4�d!t�&��`��C��ͩ�mI�<�+��o��<8�
A���SDQ��^Ѽ�v�s����KE�&ts��V�)�b1�z�Ir<��u�2�p�n�8i�'%s@�������j�6��B�����-^�E}�s�+	��PR��	��K����7C�����$� �������&L0��^-=n<�'/9l;�<Q�l%��2%!�ݒ�3�p��mR�,U�g��KRϲ��;���.�;	�>�#h�U�H�[�mNrʰ�q��k��\�������:NA6�-�N��z��Ю.[�Y=��Rk#��O2ՆI1�Z���2Itƍv�ĵs��I)�S�؝�OY��Sr��zi���f"/�OP�Al�Λ��>�)]�rb<;���x�*zO;��j�!n�.��M���$}������[l�3Ũ���_��.�JQ$�?���L�y�h��I�X��աƂ}����5W#�e�s��G�QJ�|�2kx�9u�\74�b����e��!�ȱ�;;"���
�1��j��!�n^�:�P����u� 3N{U> �@
�:$�>��	���ցg�;CW���<ʖe]��(76큿�o���ܨ��%��E}��6�E�����%,�!���{)1x��c�7��E&s�n:�ô��Bo] �	�[�\V����#�r�:1万I��M�4x���-~i��V>�O��-���g�{%e�!o {`
���߷0�u�C�.u�	���	�8ۅ��/�x{3�ڮW��ә�x3��s���&|�t����p�T~�T4��t5T����'ԚI���q��k2ȵ���*5�n/�����h�X��Hّ��t��޳���D�6P�01�3�ylY��.m6�z"�
��J�I�\-�Brx��-��t�M��R]
3��K�����贤�fXp>4	��,)�5C����4�U�� ��7�+c#n�3���X�V����D���ַ*
A�w���_�o�GC�*�����c�+��[B�ڙ����@
%�N��B�X7o�/��!	��c��#��g,��[�F�G�����g�1L������ԦQG�(����myY��b{i�����|�j�?�����O�Z�j�=v[i��Y��M�〬�
5ƽ	�	hP��\�P���Mv�|�/j@���&Yr6?�T��f�Ӂ��r�r�zV#�✪���$��rI� �Y4�{�D�]A ��a����d��C+���-��`,g�� ��0����&]�V�%�I`&"h��*�⓺��f�����G!m�<�rW�W��;��^��[1�����V�f
�lM1�Ug��
p���R54���m�39��W�?Mn�<Q�
�%&αg�P���X�U8t :��Y�hh<4�	��|otw�a!��3'�������������]�_)ĠaO�N�=�uR�~tNbS@�9L��H����i�8���_��|�(�	ipoW<����"ԢO_+Mj��-
����y.�ف�߱�U����S+E�~Z�#g \�N}��P���Jk
 Z��i�re8�+r���db�t���fs~0�J����#�\����	��_���	>D���T:Z������ɩe��Մf$-���@����-#��e �!���
u������� +^�j�-hܿ	穚��{�~f�1 |Za9��B]`�M�+l`�"�?k�H�[5z�gnc�/�L��q*1!YR�fӌ	J�i�udف]�L-T�ϑ<�K'�de���ҟ�gs!����	���]�4$��֞Rbe���+ao�.�nR�񗡲�7��)=%N�cQ"%�_��~��Ut\�D��WCǊ�.�.l��/�{����R\4��o�RW�wR�(f+���>�l�<�m'l��ɿf���n��9."�h�>TVA�I!����<�ksj��bO!y�+����^m�xl�O>���
�H9jK$H	n*�<�Ʉ6I$�{�RX	�\��*q֕��G�ELH��sBf"��m^�/��vz�إێJ
W�w�EnGE���{�Hz2�O\��N佗����7���i��J5�Q�����Tõ^#�P�r���gf�O4#ez�4�bF���?Q���ٞ�۱ӴC��#!G�j�p��%� )
^0�f�=kq���V$k	��~�F��.�/�]���*/�ݽ��}eH�֘Um�Y� ��5�֘2dd��IǊ��sR7�UA��V��3�%���^L�2��Jh��9����F
�����Y����Q|0X.5�:�]Dj����6�����6̅���%�hv�
�Y���u_=��6�	�
�S�弸�dӿ��8��ءWM�T����}��N��.��a(�Y8$n��wf�=�{�����~t*�s�^����A�!��)+	�r;P����oMv_�.y^�J2�o��]G�ro�?�gn�C���TF����xa��'��C����z� -caB�����J)��m���Z�~�7C}�hgҩ I´E��S��R�vEo���j�m�j6뛠��}�\�,�v	�L��-�ŉg�=�Ŏ.��<�M�Ow��rH�&956Ċ��fCu�1�s�V�Њ#�c�]�`>E��i���B�4\f�����	>�A��>������Ν�C~L��B_��XP��C�ӣ�#	��rV�#���5CU�,�/�� R����Zu,��ޮ8oMW4~
;Q)0����{z�u���#��Xn�@��c�P��Y�!�R���q����o���m�d���+�U;SW��w�곳�������~`��ş{����<�D�t���/�i��v��<�t�},��֝'O�g�6r���v��5����fR�U~_XV�/y�\"�܊G�a ���1-���PI�����wk�g���/mD�C?���~ �~U���W�_��ss�Qf$x���e�F��&��Ke�X{�Ȏ�E��O����j�cd�����Уv5�aVMn����k��a��1���N��|ݠ�0� �k$�eXG��?�s� ���O�.�[a�l��U�E�����s{��#�T�Ӳ�s/��M"�q�o�KT�u={��C0tӫ!$7$��4�����O����L�m�o}�������~
1�6���5DD����Dm�p��-�cwˋ�z��xd
�.�Ŷ��	P�!�0���)�"��=X!��m1��_<��w�
��fFS4�M�E&�2��/�{$ٕGG�l��e���=��R�(&���ujdՔڰ��_
l��JAxC��4ЗJ���3����=�o��!F�5S���ΚYi�	�%��vC<��k��k �8�|�+���s����X�baelG>B�u�M���(��W�L��N;��B�S��8���K*\��[4wx��͛�֍��M0���\8����0z��UᘆTr�Aiw��dU`�@�V_vC�7�z��t���O�Ǔ�� R�����ZtB^e��̉fT�M�`�&"Z�-���9��n�Y�'/IMU����}��	(Jl nnI�h��Z^t�f����;�#r|B�Xi���ٽ�B��e�W$6��=��&8���9U�c�����^�tN�8�x�^��")2f��e����"Ҧ_�4D9�,3F7j�y�XL����wT�e��Vb+]ņv2���4駏}�~��@-+��qi968�e[Fqi��Y�R�������Er˝$d��m2\P+$%�׊�2�xy�h�4������b�|yQ�q�IQ�qs�ó���O�^��UDm��ǽ��Xc��������1ԩ+�@���'���o��H���L�{�i���b]�5���eut4Y_�ҩ�[#�Wh��D%�7���8���y'��h"U8flt��1ACڷ7�[K"ߔ�ڴ���+L;J�b���7��v��a�fx0��rFG\A���{���%	��+&����#��5��'�>=� ��������!7��L��������cv���A���r�I�u�\�M���<q��+)���V���_2�֓[Zu$Z ��Ԕ�z�n8scA��P��Q����v�������e	uG9j�̾l��1!˗e�
d�؂	����~1���f����a+<)q�׺}<DK���9p�<�v��2,B:�2�4��3�ݽ�t4F�՚<s�M���i����X2j{0�C ~m�ٍ}?�Dk|����R�Ve��n�K�8�Y���
��a�����_E��A%Ⱀ�Vw�Y֏f|�ŝ�!��a���GE�9,6,E�Pݷ��<w�&��[#�4�pj������dnZ~M=��ɺ���R.�M=i/����U29�� �b3g:{޴eRWq�W���mIl�=5iB���:���B��#��"SOҐ��zG
׮�ϟVںC��3��2Z�������Գ{,s�ˈ�@��h������娊7'{l����w���Oķྻ��ǬM�s?c������Z��
_���D�QBr��	�65�)���N���6z�6�j����?)�涤�3�I]'���6��>Hf�`����������>�ֹ����qp�?d����ig5��l��{��E³`h]��WO���?���uoI1K^D��=�%B�S>x�4l+�SRe�4y��B�X��eRE�j���(�}�<��k~�s`�q.�2�TkA�'��it�����%H�����$�:� �$�vxElJ�0<��c��zX�{���U���!�ף9�v>��O�ֲ�6I+���j:0�����a�۪ >�9���8Ӷ(#�V��"�z���"#���m.�QY-��3�x������%��I�/�jn���GBHn E|�]/�^���Rm�j6���`ӊ18�`sn%���0am%���:s>�zhۯ5���� ���p����z�ݝ$� �*e;��(�@]A�kl�^9�DRARW#�KJ�́{�eU ��V3�_�~C�(d&j|S�:�D����۳'t��T��$j���Z�J���.oruk�1����� �P=�q��{�R6AP��{䛖:F�c9�~���^�[��<����C�9=���ڬH~M�R���v����r����*�j��=�D� �㇨Ř��X�NC3ͅ��)k��G� �"��1�07���߇�N�7�my�u�Ū��D9=V���VS�¾���q{�G��O0�帮2��/ԕ��������}��]��<:�?f��)��a<k�!sd��y�.)"��jA�$�+��V/%Yc�J�B:C	���&;��I���w�Jv� ���/m�z�c]hSq=Z��	��0�[#=0����|�G��a]2b�$���4�����]�Ү�d�F���[���>������VK��禩L	����шߦ��c�ޮ���a�.'l��ߖ]6��(g|2W67�z@�^�/�.!�)��M搅�8��ɔ�p����NB��oZ@M���c�~�����;G�#������}�����1{��c<��P�Ǧ��*�+ZA�N'x|��O78���q���Ł!ڀB>h���DH8�o��&p��ϼ}5���J�Lp�,� ��������^Rˉ�>a���^0�hxk
� �VŦ��O��=��O��O��2�I��.��*�ɒ��Ƴ����9�@be#l�����N�i���yz��tp��|PV�u�fR<�4�#�w�?���Ai�q���C��B�ODX�'h�S�2�*fzW���ŕi~��Ɔ]fB~��+�i����d&3r#qT�J��v�@��G-�WW����9�-�ae�߳{Jg���v�� 4��:�:�^Cfw�S�eCY�th�:��G�l}�����$��ڛz*�/J�9�t�a�:����f�T�ب�p_𴡏�'NRY�=K)�"@G�ӗ�eºg|��H=D8s��K��D�t[��'ìH>�^�[Y�1k�r֦Ө��-.��;g��W���� �I�N�Aϥ�r[�Q]+����9����s�1�^b���X�i�3�N�:�ݰ�d]�2E|2ҷ(@��"G��f;�&pp�wC�[�TA�:O�LpG�����$F�߷�>	�>�z�v�E��Uc�ĝ:|l8z&3B��{��q��v��vs��1�؊%.ڬӓ7�_���~�0P��uF�<���i(�t0�H����f����-u��y$��b��vs�b۔���1�m,v�&�}��p��D$��������Ra��4��ڝ�p�<����t��y"��z5�h�?X�q^��/��b:�
g�{��T���d6��)�d�R�Jʻ��<��7
0�~
���e	9GYÜ�k�o��?)�b8>Ęg�l����k�4����,�ŠF��{2 ��ue�@�L�fl��w5��I�R%[�Z������Цc=��php���E= ��a�H� ����(�c��0x#��רv:6���^ʎ�b)f�)�����!�6�8�!�`��Qw�6�LAJ$7"�	R{(�,�Y������}�;��ܳ̀}Ä�����u#�6*c����a��MG߶C6R���^Q&�ۉ+6�TG柗%��C�d�Y��BUzR���ȶ�R�b1��En=� {���W�G-0��;��@G��ß��3.�Ů��1�šK/Xo�~��g�����N������BG
���}#18^��J`tx5cqV93��7xL���mK+w�G��r�+O4ζ��ϲ�����×�0#�62�)��0��]���Mѹ�'�O��
~�$#����Z�O٫A�I�bI7?��r�</-�8�c��׬���3y�V�X��H����M��Ұ�BƮY��PΕ��p ]�K��Z���HV��oEA����*�~ԽM�nCw6		�Eg_�����\��&|���D0	�zFk���0��D�d�A�A[$���h�B?�qTL��\@�\(.q(>9(щ��. ���w����55�Q�Kh���|j�:F���Bl<D��P���j8�]��Ep]��k�o� �,IS�����6n8(A6�)׿q��d%mO�Y�%��R��$��S�$/�,ef��Ɍ��.�4�=9�~��7���Ap�����O�Y39@�7�:,AἅV���TyǋL���:�7sz���?QG�O�tX)�sQ_o\��d�?�M!����2q�6��r5Ac��K�`	z�.�ou5SAg�j���r���k�-�v�%|(�ʟ�Ko���.$q��!j�򙅸7��9� Y�N\��:m���5����y�轖��,d�-�iO�@.��� �M�G������c��/�z4�U�D��	疳��҄�7��]Ғ��T�l2=)c<���2ܫ����6��T�|kZ����,XdgR<I("��H��<;�4���'�Ұrd���VM��Q]Rb��q�Q�_q-W�Z���w�w��<|��?��0 :j��v:�o��N���@?t>���A��}�S)Y?�ߔ����=���׻3�!JM�-�7�ԑ7�1.����9�&��>���}Q�L��bUW4�ɒ��3���Z��I��2�*JSߑ��g���8:~���UV���4O�U�_ٝ��z�B���w4L�x�E�Ȑ+�W����s�΂\8|��eꯠ�.�~��C�XN�j	�;c���l�;}�D��<�*V��0��"$;�;�R����W�Z��?wի�x��l��t��"�Ԛ�^ `T�����{�ͥ��(i��p��M ;��Ang�H��&k��E�Iب\��'���mi߃�ț�y�`��R�'�6_��<�E�&�p%EKn熓��F;���<�Z�
QX%0�=/)���}$��W�&rSmA�8z�F��2��:e����@7�U蜤Q
�T�~#I�Zdǌ0]H���K&ȼT��"�-�d�jF^l�����+�o\,$�[/�G5���VF�����c}JQK�pc�����P�ģ�)be�#OL��/$=��Q��>��"���������H �,8�H1��"�pD9����8�O��(xϛ*�Ȯ
WL,�XT�v��&h�Ɇ���G��H�(�r�4z��1g��-/xFx���j�Z�!t�첗J�p!+�c����5{hnµ&2�n�4��VMu��t�a�g£_t`v�>Z�]���í��悲]�7�f�ϧkf4d�L<5����L
��Ӝ|���X"h>$uݔ-��9)�눻��@y֯mֶ!~����-!ݵd���� ��BR%�ZO�C��dQ�*���n��F"�	B���;{�m���),��G����NPV�V���C2�gM@1=�Hχ*��]���u��2�p �n�4OM[�������wr �L�
kFī�EgcY��`������X�#��7d!3�dR�î��K�J�+_�
ir�}�dׅp'���P��͠/�
EYb�=2���[!Q�Z)O�&�^�m�*�
�_��9�ۉ�a�]n�}'��2_(�2��r��b���Rƣ��w����kBڼ�^�-�E>�A�6�~�L�8+3���_*{f�v�vXr���87#Ht
�;��FkkC�红o)(�)����3��o�����S|psO����!�t�;��ʽwE�s��O���pD�愰o%x��(b�%��h����Z/pk�@C�Y��1O���=�ڥp��Fn��ixF�p��|��T��3�<=wv�d�h��sK�V>���_s�[`�L� ���bP,n�ԭ���%����2�k��2�`ǣ��}Ѱ/a�8&�0j���r��g%��s-�0�йF�3���DI��7�V��z46��/ȹ���´�P�[���ț��W��u��8�+ �F(j�Y���S�8���Y3a��	 �W5�������ݚi�����߭uu�aɃߟ�>����Ut�l��Z�r��,1��/&R|�ڔ9v�^%��c��۴ʻt�/
�z[��>g�D����@�<�s��)�}�j)��,�Y�V$#B��c��mvqy���TZ��GW{��i>�`�`�t��u���t��H�S
�$��Ҝ�^#�9D�理����H�`���^~�"�2�o=�˰���B��0I︔x�4�S{��R���E��L��,Z��r�~���6��QO'���:Nnk�|�-/��O�5tU��M���q+�^,2����/p;�ηi�m& �A�U����m�kw�)`��ܷ{ ����� 	� )Ft�X�Bh������%���!F�k���@���چ�V���#��������G���K�?N�x�K�0YD�f����Ac ��h��C����<@�@��O�S�7K��h�<��T��5B�]��E�ͣ����0S@Y��{���g����R�/iH�Q���a��k�lw�>��:0��S��)��/m���&�-`���;�3k�h�"���ID�m��/p^��R�����jU�5���Uqf6���I��i?;t����Y��o?�we�L] Dڋ�!>� [7 �r�sB�ط�K3���+�ax�&ܴƛ e�C��G�Ɲ��!'t.B� �(��9�+�uHz�*��ˍC� �O�7�7=�D�Q��,�G������j!
{&ش&V=kGYɌ4S�Cb0G�fgq.a�.?.7U6�W��+`�Q�l/�n6��qnƝ:g#�ƴ'Kc���L���AܢV��S���!��6�yM��ZPa@���� &61c�ߢ����r�5�'��?+G��¾�8~��چ�6��S�������B<ϔ��+5Z.��S�ɫ=�Y�~N�_Z7\�VF����tI�����NÞۻ�/��f@C�-�}��|Ȣ��%7g��6��d�ӻ]��H2��^N9�=9Qy��j���V-r�x��ʔ���8��,���4:�n�t1rm���By�&��W�K\{�,�kP��lV��[��ܬ�Z�!YZT�����cI@�q�4;���s�3g�P1�(k��g�?E��3Dy���[{y�#���V�a�e;���KE�;q`{]��̡�� P�s��ާ���0��u\�ف2u�8k#�1��9��:����%x;^e�Wxc/�;����K{h�� y�1��)�R���uXľ�+��N����M�j
rL�����-�հdkPJ��#ip>��Jn}	�js�9˷�fe�(1�4aij�GV� �:]-�_��sb>��������t#3y,Y��p�o:|�p�otoc��Y	�qy�9^���HXY��:Y9�e��2<�!P��%.�%��iS�FX6����8�x��p>l�^R'jb8m~�^$B������]�X����tWX��p[��7=��w3ܤ��>�7s�M�~I�`h�?�y�����9�RZ��-w�А�^��V/G����k�|�D�dA��@|� K*��'�����UM����l5}�o��$���ŋ���t�tY8W�״�r҃�#q������0����-�V�=�ɧ��:�R��U{���zN��e"����a�h@Ĳ��X����(�YLf���~^g�Ӳ����M�L��ɷL�?YT�Y-BR�X��	K��Xy0A��C5C�є87QW�z��Q���cBc�gc-�d���/�sF3���O�F>�	?�A'����O2�I@���HjG,7��;k����0����=�C�Y����k����N�*����z�Ų�
���x�Ll�*�9��,�Q��&6������㞡�Y*:�D���f�_f�0鎕���}Џ/����x eֶK-!\��N3�
� ��t(���o�׍�]��65ӆ���m�`�GY����/JP�2s�д.�-�v,~�4��Y�T�޷��YX�`�`X�D��0� �ϵZ���a�Q]��A�m'$�,���}6 ���]�';x>���F� [P�J�k��V̘��g9�X$'�`�4�hS�YY�7ufA)�R��t3�P�����"��؆���e>�2�qdH��O1���^7l�~��M���g=�k|�N��0	�D�����hZ�LZn��`���#�2��� Xƈ��Q�J� �	���5�̚�i3��!���A�{��u���z6w��b�:3�d��T�l�G�%�J���i�Z��x���EL��b5����l�}����KX����Pm�+<�u �ar�e{>��&������F䈴�O`���C��V:4�u����G7{�y�E� G�{��nG�M��3��I	�Ů�+������<c��
��>lȌ��ҚZ��,��lRW)����h_�H2�z���Pͩ�\�?� �,�W�C��'���S#���k�](7���������o:��z#����_uUPl�ߠ;�QFj���=	�e�4'�ӡJ,XP�zj��m:.uv?g+�Ttu�{ۤB�77q����~�7��b2eٲWb�Jla��DG%�֕	{y�Bg���|<U,��.�ԏS��I1���L���=��Hɪ�fC�C����6z�������
��6<���,pBC�,�	9rgr��U3v��0��>76C�(g�7�;iq�!;���B*B�1s����-n�ֳk��-�*ϩ@����55�Ud�"�w��H�?��sa
���@�_z��<j��Nuô��1)�	�=�=�[��l0YC-[2�l�\��	,�X�߈;i�:�bm��q�:���_%ҏGn������%��<X�����0&I��vcs�W������9Y��i�_N����S��V.¹@HԪw��q3�De@�ie�:;�YZ�B�x.�]���ѢZԕe?� �4���V}�C�u���Iuo}��V#�5�5��^����W�Z��xg1�0��R��';�;^lڰ�L����q�Py��%�j|sf[�><-��r���2}��[��"�_�qi�ҮN� \�A[��AV�|�2ˌ��{n���mqJ����f�E� (o��yi�q]��Ȧ#@ �oV%�j.^_��|b��2��T�v/hf��4}h��F$�߽ٙ@Ա���}�N��"w2^\#�ap�]��ġI�<5�&KU 4V�;LH��롳e��uz`��}���Z��i����q�O$�c�/�[oTؐ�ד���]�gJ	�I�8�
����̭��ፓy��K��%�͆#ãx�]�.rZ��5��@�?=���5�?;N�-؍T��*�
�g{T����T�#� y��?!���'�^�
!t���*��X+Y��L^s$䙷������YN4��B��B��H�!�<�g��~���ƬL)�/�Vp�ӝ�k�^8�w.dlNr3a�h�>�˽{T��W���-=V�y���D_F�A��S�I.����m�BNh9�>nu<ˏ6,��$x�y	�D��� ?xQYo���������hZ�Z�eF\����k�����h����M�ʮ�~ 8< 3E�!+����WNY7���E������Ȇ��-�~���JR�SC��gZy��ql�������{��a�)N�gq�}F��*j�����Ztkb�s�v���+Jy�TJ��L�p���7��^B�%�3֨Yg'^0��gy�c6i�]}�Q�79��4p�n�G�Ղ��FM���q�I(_{��2�3�<20�}O<�����E�ّ�UKĻ@Y�5ly�����
#��k����w1�=K��E+�������s�;�/�@1�J6W4�O+V��U��S-��^����ʑ�5�0�^�8�!�EM2k\��v�����B�V�$��Yt}avf�믭*�7�H
�2?5'���w���v4of��^�X`���SM�L��JKY�|�^��X���m��b�+ϡ������T�����I&Z������Q������(�N82wm�򋢮Ra�IH���ͼAxm�+�~O���?�:'z]v�U�4Ф�f*cp�J9e~�ֈ*V�(�܅�T�����3��֏]���qV�k��ޝ+ݏ}���B�O �gS�v�*eg�AU��X���uG꒤�l--�����0�U�~wל��KCTD7�T �.h�ҚO��n�Z�	�|m�?��WҠ��,P�ژ�a�4�3<	��<\��שY��΂b��ӊ�
K)od��o��@��;p�k���8Ъ�G-Q�/�zq�� S�����i8?ö:�w�O@yD<N��	�=D�O��ꄻ��t�r�<���Bi��𵿻�~���Z���H���:�7T�M��N~Ќr^��� ʛ�:h	�y����ؒ ցC�&�3��梵e7�JZ����є}�}��$I-�dhO���J:�.o4�(�d���K��4���-�0m������+�/��&vt��`�`iM�V@�ס�����hʈC�A��7Y�{�֖�(��ӕG3�_!I8#�Q��67��Ůi(��T�ko�>J��W�?���L������&Ԕzf�>#���E�p�3�|G�ˆ�C�*HT6�H�4-:$W$��\�����t���P��,Ps�QW��A��ɩ�@��U����l�2���4RDӻE��G5��,�%�x�Y�X���I�jV���=�R���7����=R�D+���"n�H��C�v��*mV&�=��舊~M���b$$�l4K%4�D��NF�-E��b����'�uؿ2R�����*N	*��5��c��sk���nL{�!,.%q�C� �ʋG�;�g�5%��2f�|��&X/n��}��o���q�Q����у�cax���@��.V''��� _�#�B:B�Rô&�Mnd�s��&��+^�K�aJkRy·�:&���d�*����a��R���}{��!;K��� �SzlT�?(��<=cfΆ�;����}lr�z�;�B�xU�
5����!a��b���m���ΰ�/I��,}$xS�����tb���|��r��]�~��[��wA�!t�_G=�J��8�,�A�c	-�9=���4�p��D�_�N��O���z��ɼwܵc���K\,����Pȧ+�px�W��8y�I�0 7���ҙ��qPU�L����u��!�A
J�̞��[�K4����'gZ��í񀳛r��c̤Ki��z�F?F�W��i���3net�=b�A�3xx�ߙɗ�A��E�F��
|������S��hh��_�0K�,٨����y����%7�v���6�OA_7ˉ�B� %����H���4C�Z�{�d]�b��32�-2�L���!~7M��w?ڊ�Hѡ�a�A����]��Z��9�sMI��
xt�\c������#� �R�L��HԦw���E�碦��zI�Ap �ӯd�C��O��I��4g%�[N�r�I ws�6ɠU� I����)��dFcPE*B��77���P�Կt	 @�F�D(�~�]�O�~=�������Sn��׭�*����>D�" ZM�)�e-��L�le�����_����8�~�!�_�Z��K���Z�*=�1ʠ�Z���=.�4*��yY�e�o�#�`�������]_'JZ�*��ת%�7S=Y�_L�Q˝z��׌��_>����4��2,�ߤ��I�mij�QUC�����zĺTt;��*���8Hb
���s��/g���O��H��r[��X{�A#�9Ȁ��8nX��:F2b*���l���K�"E�x�n6��L�S=-	 K�����q��y�Ԃty�A�v�ꬬO.e��E�(�UB����`�I��M#���8��TgD�!����>T�`r�؍p�S;�.��#��e<�:n�@V���x���`fGz�ae��B���h�,
tr	)����$TC�]��)�1C>8j�J�5{�%?���!�	L���T�jwVj��&��UԧOs�KE!���� ��4
 V�ʌ$'s>��l�-��b���w�qMrn��]c�d؜;��8uf�TP1�i?ZH��V��w��Fڼ���
u��uЛP���������6�AW�D�K�24[D�+W�y�ZL�^jX]�9�O=��D.x�W>��#k����Th|��d��f��'}�(N��*@�� �T�����c@J>g������sb	ހ`�#�m�B���S��_�x2ť�8-���ScH��܈�~j�Z �M���t"������i���C/������P��']��`+�^�4�`2���l�K�r�p>��d �oX)�lӸK���[�b�T�/?g����,��#�[5P��F��)���A:����i��֏.�Tu/�.w��f$|ߨu�|�ٲ�a$��M<'N���;F�ll>�����P=��&��8��FR"�Ԁ~+���W�F�XЫ�Ƀ"/[Ո��>�:�!KeҶ��:��L����.���sr�-���՝,��M:�O�;zȠ|���X��S'��I�{�}~�k��:�"L��U+=��H �D2\�g�j�fH%����E��W/� ��u�Y��M�sMq�d����������'9H���C��2�UZ�A�%yp���s��1[�����c��t)~���W܄"�m3=}�KS4�j�*�u6��o��.��0�MǓi�����b�IHt��i��17p	,���?Î(��t�������Rt{�r�,����h{ق�A��W*UR�?rM�e{����;���ޙ� |��� ��<<@U M
b\�J�d���J��i�hث#�ԯ"��S�{�Z67��Ǡ��\Q��\�z�4���]�q�uz�a�r6�ẓ�o�=$Eo��ˈ�/GX6�JJJ�.k�;Tg�K�cJ�1��*�����B6�T��#��7���ڨ��fvy�.pIX.k����+���@�^�)�;\T��&������k�M��8���F���2�jd\M�tf�W徹?�˜j�!��_I�� �� ��ZEZ �I����#H��/�ڴ��f-.��`}9v0TS��^���z��RwY�b_\���,BK�HB����� R@��	��!� ��K_�B1Fr��Z�T�,�{c�Z���+��=�J��q@�J�'6
���@=�0�P[+{pxW"̫v�Rw, �<�>�-v��"lPy�J��'��.ұN	��7�^!�a$j�61#|3��)]�!2&�UH ��D����,<��q��)��{��>�y(ې�m�_���R�8{��t}`��^*��G�O�Tv��Ŗ��W�N ���R5&�M5~����L�V���p��H x���1!�7�
��95��}S�O��(��x "}Pau3�|� �;q��|~�B�<r���K�j��n�M��+K����M���������_x��L�����#;�5��0pu4�$��`FC����\}�#�(1<�+��g\�X��������z@�W����$��(*\̷��L	��_��L!� Pt���/T���[��]���w}�t�@#mjoΤ�=��\d�(�މvu����V�}ES} �Bv�����y��ІK���|��1�J�9THBE����woL�X�zO��.Y���g� �N��tI' �xw좱��Hs7�yG�f�~2���JX�=J^�(���|�b�*	eGQ1���b����BO
��O��C;������2���"_������d�Q�X��Ru����֟x��~��y:�LhM�������6�w���H^rs$�~}�^�\�9�D��~���
rp%��I �i�y�� ii)_��bq}�L�Be��9��(.(5��J��&�J?g�}���@�M��i��JW��I�%� �;S�ፏGDKZZ?L\�x�,x6�k�Y�	:T�l�1	�a�C=��&k���.LXg[Dg6�'��U�r�F��v��\b!1�]��S/���hi� N�0����|�{�p/����2�E4<��,�xS˰3��0�Tގ�7�����m��qG�@�����<�d�H�D�Y�㼸���IF-�� �o������w�1Fp�2��[����B*kH�?��ӎhQ�l��	���e���Q�%Bg(0�	�
4���`�0�
���'��3~+�F?�A�*´�����%v�w��0�-X�d��eyG4���M�Ɖk#*=pc2=T�6a��~W5�yQts�o����I�F�����"V��?�?��ef�����9�1n�uY���jH2pa@�c��x�����D��yθ��տ�F�.�F�_9�k���f�	��[$������S�ozX���72�}�5���J�f�#a0�3|��mC5��)u�ƝբqN�Z��#�����ޫ�5��2��G�a�v-�lzVq7T���a$2�;�a�#Lh�"���3b2����j�N@���R5~^f{q�`�,�>!�f�{1�%�����e��x  Hu���;�Ɣ&����i1��*�/ᰙ�sH�a�Z�����q�m1�Z��N�~�L}ʷ�	5�����>`[4ً����wh�&���~�o6��B�����(1�}<;��@���*�K�:��Yz(�R �퐟�cJ�6��q=�̲u�<ߺ%�f��}�/�J��fA���g3|����= ڶ4��}
[% �G�G`�7.�W������F����(uLפ�5_����uD�l�y?��d�k`A�Fq#uYu�+�bp�L����mN�����������b9H�pZ$g�w�P�+cn����=P����0� ��xA*�[�+��6�����M�� ���6Ld��;E�Ɇ=���#c�Ph-�w���n�� �&4i��XGT o�+� ��B�^��N}'f�p�$/���IK���e�ӗ�I��9�߲A6��x�m��$3.����d���_�;������uR�?(�<_��B�nmd*ص��Jk����C�N�ϱ6�@<�$I���j�=��&�U[|��]�Z5>�%���n?�Ua�$��F�M�1=��PE���\�|A�|�t�O��xm'�l<�YlV�pIe^�g�e��AJ� ����]�.�%�z��"�@��*B�G��5�[��dɎxH�.?Yx��}*~�h!�;a-J�ey�k{�u���1�-"�'��w[U&��aH�8_%�LlT[��2�V�MhN|k�h����Vr�
�m(M���8�;�0z�&dA��d��n�5o�n?E���B��-K��)�X�w����}�e)�o`t��?._R��������4ԅ��o����N��n��pM�^��8���a�]hEr� �0`��}��h������}�=q'#{r� :w�4P��/�l��4���W�n��G.	�r�bB�*J��,��Ii�8heA�<�ٱ��3�4�[
Z��6[��}h����[Ƶ�)�r��bꛡ�A�� n����=h2$���+�B\M�I�����wh�w��W��]��#F��gH$�{�`��NTX����ke�ݎ�ڂ�ҷ}�%'�'4�W��t����7Y���?ڄ��1���Onɘ<Ղ/9�c$�{֫Q��G?�g3K����DU�Y�x�`�
���{g4&����q��X�^�N&4�{�,q5{M�J�C�}����Zi���S�弄������׏�ıɸ�����2�x1~�2�q`����2�b��}��塚������D���KF8��Pm�Iȵ��Q��x'H$�VԒ�X*nE,���XO��8���[���W*���8D�he�1�oR���ȵC�k�4]Q�/�ɭ��h3H�(>qy��h����v����`�+��Kh풓/�G��h�,�.��|�X����z�1ggd{���\ H;+��c�ԇ�/2 8��ɂk�����O�K)�k���^4��>�$��Q��Q��&�F�H��3�������Q��p�!��	�{��X�-�f��1T0|�*nA|{⛉>�<�s���� (���,_.!�W�@+fn,}����X�,�qt7EW�'�3����h����3�]�����=n �ʪ9�w��|}���o�G� 6�}�"r;$��������D��&h\�f3,Moq��:j�ͫ��FRh�Q,���9�]I� k�H�{�S�x.0�]�`	����~��~Xso:���iș*V��<y`6��N�i���E�f.�������5��i�G�\�GP=j�&0s�����E��Y��h�v�~�>ѷjB���t�.举��y|$�yD	�+��o�D�S��?H�������7���)e��h$$a��D�B�w&x������z���v�%�m�%�a��X��?��AW71ɸ=TbM����X xUϻ���a0�s��Y)j��tM�B��1?��M�$9(�#cdr��4Q�{]pUJ�-r6���z��u���Ƥ,�"�<z�л�%���
��?�[���BLh8����/\9)�,�U4��k@>���yB�oq��ɍ��%p�^7�Z%��������hyk[q����t~�t|cb���b��.:����&�پ4�i	��#'c�/�"�|U+��i��>h�;�;?���`�e[r�cz�Z\+���N���*I&l�ȱ"�;��{wA%�l9��!V�Z�x��,��O���6�ItTY��l���@J��� �W�ֽr��FC�r�8'JD�6�6�[��2����k2%G�edG>���~�2Z��%��B椳��
����8Կ���?�ߗ|[>�U��AږTh	J5��7���%tl�SGD������Đk	!�3.n�,k)�(��� ˇ���U+$��R�9x�ڭ��_[՞�.{�Ӑ���Heou��ߦ�����V�W�;t�0qu�)�R����U!�y)?��m�R��O�A�C@���n�J31e�&74%�8�3�Zg������ɻ������������;�wt��~
�d]!~>]H� :�_4�|?Z�N��z�G{&c4P���$@,/&��<i,/�s��������Z��gs���Mr�נ1�K�RK&��t��q���@%�8���f	�N�#�5O�{6������e�(}�:��(�6r+GA_��,�5O�I��jCr�E�$!0��shq�6���t�x{EÚ���XC&�q2��*I:�� r���qy�^'���^L�T�Ѻ��bwu�)��r�!���1<�s�� ����Z�s�ɬ �U��8@�+�;���C� 
G��o���KQ�0��"�D	������P|aom
���jJ�ǅ�v�ޙ&T�%C��hvݷ�#����|�|*�Hg֏�J�������g(c��7����[Az�o�+~ΰS���:CXwŔ���E���<��#�B˖wX��+�/x~r�l��mq��#y����G��UY����uQE���ӋtN[⼿#).S���B
k0t�KzDhڥ��ER�H3�~&i/�{x�?.omh(65U�*��d�(������T�|f�cǟ��Mq�-ME�\V<J����e����3w�m�K �~��w+�����Y��,���%�e
�?�4^��;p]L��[æ���:G/9_@o���1Քv�℆?SП� �+tظy��f�ŖVt���e��\�� N�����C�Սd�K�f&�ñl'���09�?��]K�ڮ.%,��{�E��8�䈘5��[D���x�Үq�JU6H�Lr "?��ƋӮdN��+�04��z�n���c8�V���H��qdw��F��Gn��'VN;U��?څ����}y��������sм��ތ,:�9L`0J�~�l���3h��n�S�i_�������S�2̽h!�-CЪS��]����X�K'w�HN�(��Jl�<�k���e�3*������}��<���Y�!���"I�z4��LC�o4q�BL���Dod<[�v�#��;(6�<�V�w���o/���N�4�nZ݁
�<�!%z����b�iI�ms�Y`��u�%`XSy3-�-���xʐ��w�>̉"�>�$21�΅�Ǿfӕ��Z��{�:9�j3dϡ��k�ͬ����(�5��t�t�����5����'	���A("T6�Ԋ�LS�x�W�J�lZpϥ�	�J�G�Hk�)�f�P	�G���9橞0U5e��	fZ��/%�@���x���$��������g|6����^�!���騺o٧kx�^K�<���y����@Q��qb�t��'���[��y��*��>�֥ȏ�5�� J�/B��J2���x�ʀ����G<���#Y�ݦ� ��vx��~��B���� ��/FhH�'l���mcC��U=ƺ��sDo����FMX�����-@���t�<�`������b<�q�"4������F�*\��v�'�t��n��tWAqC,_C�Y����߱�e�4�nX�k�r�3�ֽU^Z?JA,x��k8n�����h�U�G�ׯM⪬���$�KG"�þ����~x��˓�Յ�nΈcb��W�ǄH�^o��q�9�2ۋT�y���`���'Mֱ���-7{�	��g��3��E�S����h��1}�b5���[����x,�~�l2o����vi���U��
:�M���0ϓ�E�M��)J����xP��s|⟴�M���=";���PLnU��Q��vλZ�ku)#��Q���|���
�qt����!u�o�?��n�s�E<� �V%�^)�Yjs��'͆v�V�ڹq��(����E�K>r�� R�Q�4�?��y?Gp0�z�AV�7_�N�_e��gˬ�gC��綊ؚa-srCLo{m���J�a�\Qq�ʰ�� �d�-��Y�㕽=��q���,�N���k�ux�~j,nr�z	
p��5!qk���6�l�Lw�~���>�n�����ȷ݈��D�5y'n`��DC�U%KqjZ���q3|;?�w߱�c�@]4������Y�d��ip��o�ϙ�A�]#�\;�&_Q����1J3gi��H���%�]��5�|g�,��:~���Äp|O�y��J�Xw�^����ȟ��2� /2vOxTL�q���6���a�Ԋz��17�gl����{p��I�_ �A(��K��ș���G�9�>�Z8;Ui�!�RU2����hC�o�>u���]�E��``K�eh04!^�M -r��b�f��d�����f�G?*t��2�$��c+���?��\����E߾����!����]y��?��Cf��
�f ڥ���$f������!������Z��7T�(Ѻ*�/�7ݡ���"q��hY���81DWxk���Ϧ���Q�Tw��P��2��g-���m��o�3�}��Q=40ǒI��;��>t�4��$������� t��SNꖣQ��-���F�X������r�A��HO��� �q��:V�=5�??*�D�2 �R�����l�p�p|9A�E\Ț{�y�w8o�w�9�`����^w>iQ$���!���\:�f���-Dh�i�l0��9b�iZg�1On����:������`�4܉���f���!���z�R��u���9�s`�������4��X�x\xyr���= H�*4"~/0b���|�a���@��N%�c�R�8ԥ�dbuxb�P�Q��C�7�zNl�1���D��Щ�q����6Hv���#F� Ի�dh��΃�/0b+�t�:�p�¼���]u���RE�� ȥ��*�~`.#�l�+�2�{Ӎ��X-����f�
y3���'��	�Ł�+�Kp��.������'%rU��IX+��<?�DpH.a�q�ra���Nl�{3p��ƕ���a�T�K����<.���2�g���\�hB-�����9��"�YV�AG�҉4F�Z�R�Z�&ܪV�H��'IQmEN��/]Ȏz Y�{�T��7'p{O5��N�Fgeuv��^�����j����Rl�����%�{+f�h�-TǢ���->L�bXTfO&s��[���0�,v����c��]���}���!�̠���~@{/��	���\Ɣq)I����/��Θݸ��Nt�H�/y����)1�-�b@��asԩ,�h�}Q�װ�9:g�6%6�A콢�ɩ���K�%�`Fi��&��M�yZ�9���wƢ��+Uo��GH@��ChHA��I��6�߮I7��
_3��Sg�9�h7��\���H�Z@9W+ �*D�����*� ������x���+"���%�V�7I����c���BN�T�ϫ�x�rР���ԋY��G��8�g�1a뚜s&_�2�:��&�`��5��r9̈́�^X��0�I_�
>�\u��Sŝ�b�X��n�\�0 5��z@�7�Ei�[�o��Yf~pY��S2ւ��s-or������ш�i��*��q2@I-�]��:�A�0T8<��ߣ�S����w�V��%���* �� 2���u^���C��Ȗ�j����N���O����܈?�.��=q���5��]����)9��%�b�
�J��W�D˫��U��gmYzc i��@�>�C��m=�
-��~����$�э.q�l�w_��w/�"=�q����:Yh�p�*��:�0vk�������\�R��W__�}��M�N}iӾ	`�R�4�K�w�[a�EZ���KZ>;-���2`)	QnG��0=*-���Tq>�hu4 3��-�̪d����'s�{_�z~)*��)���J�>���s���'i��gZ�u66�v� I�$�&��m��t=\%a�L/D��_��}�I(�}��I�0�N<��t�;˒,�-)!�_�pXny7+��{�`;<#�N%5��4�b�s�����^3ک�n'�
9a�ܳ�b�zOD�!�7�jH���C�JP�`(��������y��� �<$�G���%otb����ӽ�5u�kԑ�H/ܺ|���18�ޡ�RQ���6)w�n<��k;���Ù}۾Q����ytuHI���"����L���k��1���Xل�ʉ�P֚a��'4,��W0;)�������u�ެ�x`ӣ���EWz���Ň4^�K��}v���	��˪j�r��j�l�R�S��rK9L��j]��J`�$��=��S�^$P��-�ȦR]���������P���A�{�ћ*
J{o6�C+
�K���t��D"�������f�}����r�G25�/p`��P(�����Ttp�x$$�i�\#Aq,m��K�\G��E	bA�G;c�;��;��@P�y�G���xFS���-���+n��O)9��_��:w��-nK-�o�3p�u��jDb���`l��J�_�q�F|]XY0\u��4�4,�Y#9F/Zǵ��E|��iP���.�T+R��T��h��mL���FȔY-�A�"u�o�B��X�K���>[��EÊ��/��c�s�銹M�x Hh����,L��İEC�֒���НjgE��r*n��x���Ax	N��X=P@=���9�V��}|N�P�rm0@��4��*�)k�X�;_P����$�:���T���r�&�֐:�\�X$]A�vks+����k��6��}y���1�j�^�.�A��5/�����c��J]�+���<��熠�0��'a͇�}R�j�3_�N��d�Tw�p����ZǇ�@i��Y�c��
��z��啂��}@|�8*�� `S^s����X��'���ߐ%����s�t�T����\|�0F\�צ�^ж��W3�D)AM;�G����(��q�/�T���}3���P���pp��ӥvPx����c~�`u��Ұg� �����3��2�Ez�8�GA �&��N����:~�P��ě��ZC��}����UȈ�ƢLEX� �u+{�������A�VOa8�]ެЍ�_](J��*z$)[~Rm:�4��NI�C>�l�N�s��M�/�5X���f`+���v�B	�o�d"���8wS7�K�3���&N�3������lf�v?G�du�|��GN�����$�Z5��Q��A�5��j(�^̭/�z��ѫ���f��U��((��D$"�����1�l�� nP�D%�k/vPQ���l��}ğ��J���	�X�WZx�2.م�E��{��3��*k��܅��x:{*	�@� ���#1D)B�>��rhIN�a��?*�|��