��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t���0�*z޻�1�M��}��j���@���v���I��L5��ϵ��i=H� �b��.�$���I�83���fA(P�˯��%$�^J��S�xe�b���k�6�©�JD�f�/�aS��4ڔ �DK��9�ս2@C�.{����D$�Y�&&��+�xYn��_+���N"�����H�o��L��)�Қ�Ώ��|���:{�Qx�"��J�F��o���[����וTe�;�ɛ�t�����^���,�e��Y� /�F����o�m����q1ge��g��5A��('u:��> �go��~�^�U�#�[fx�F�+� *�׼������<ƶ�A�JEkg{"�2l�������:�`i_QK�Ki���Ji�\��p��/�!�E�Rj������@'^1�1���.�KF�C�^UM��_m�D���|����������Au:�#�}��!��Ó+>rx��B���$�E�����B�v��^7��	m,	1�D�[�K\���e�e�/���(V�,��)�:�J�\�y���6.�V�Vs�;��A#�2}rF}2�#��c	� ���s�ੁc��Y���v��Z�/���)=}A�8�4K�"��@#�0�桿�Xs��@��tZ�f�+�F)M�N	9�.02��<n��e0:��t���ʴ��KإL���e��'DOw�t�M�&�<_b��nx(�0r�&͍�DԻƺ��6}�j_�Uj�G8/�8q��:5V��*��C�=3���VWS��_�g%Eׯ�0�	�<,j����&�N�z��Y�w�����75&��$�`K�Z<��-�Յ�XJ�	����q�";�ٝٲ��l�	��&U�Vb��p	��,\h?&ۨDġջ�v.=��b/��ۤ��!YP�����v�+4��Vx��Sm���[<!�˃ ���`���(
�-'h
�p>F��k�v�G%d����IO�O,IҤ}&:*.���}�)&��F��R��J����[xz����؎���S�d)fEM�Nl�`M�KhD{V���8Q���C1hQ��-���d~^�[=ܹ�j���ȉ�I��gϏ�I"�wK:�\W{����r4�W+�r0�7" �x\���홹�7Bt�x����gp~�Y=�1����!�i�}'l���������6/�/�����	_���P��lk�h�C�n�����!C�^�����E~v��T,%'��a'��]�Z	4"g��B׬-�}u%�h<?��2UҲ�-+�)��Ҏ	�"�46�m�?� �K����	��M�ͥ	n0�W[��Ku�/^	��3��v��`���JZx�.�s�R��Fjb�}kP�?-� 6B�2��U�w�{����F��
(���&�X���<2�e�p5�Eջ��dgz.�Et���Q�?�� ���HZ���;�ɂ]�k�.�Q�3;BSLN�֙�<{I9�OXs�2�B[��O+x�ڔ�c[���K�0�GO�RX����n3���ڷ��?����U��v���j����lR/1�{�W�>^­J&`9�e���%',�|K�����l#����T�i��� �Ps��㐓�:s�75̺mY=O�K��R�&~����T��d��s�F<���'�˸�[��+,��c&��\��Vp}5���9��0yaW��!�3�lR�8X��r�·b�F&J�+�x�h\e,�L���{������䙐Z&W"k[r�D
��E�ܼ��&d������нW�ϱ��Ǎ����4�A�ͧY�Y�/W0���D���k&��%��KZ\)Xc��2o���Y��x��&����X��S�b�0#S75�/p~�? �7�My
GOKQ��5�T�����5����#��_��ӎ%��n�U͚�e?�`��WT�D��7@�('�!�k	�o��nQUt�V��o�?��6�D�����KE<TcS�8���x:_+��C�?
�"n��+ɴd�z9bcT<��1w���p�dhnpJ�>#j��sI�Ҿ�D�2|%6�z�9Fd����gա����v�py�S�o[�<S7�b�֞� �X������˥x_-���1R��w��T6�<�,�;x|��lI�T�s:�#^�E��\x�n��B�`|؍f{,�VoI����dL���#�P8��S2����	}brn��L���f�[���'Hn��!�To����ְ��GV �>�,:�'aҀ���wS�hgҴ�FQ��QO��[ �T�7��Q� �+4v� w�>�eS���<.�%� šG��)M��T17���� �Zv�h�:\���^���rc�Sq��~��?z��m��N������B����[ja��r���j[��������N9��%��!���fU:g�����h���Ċ�l�H��"+�z$Y�0��`�ܺ�����{c,E��s�5�)���[���{:���n�d"�/��>�V	n#�klgK��w*T�E���)�����Q��-������A�NuM�t�7���	�X��y�\��: ��IÔ ��-���i2X*z5��(��ڎn|<gT~ӽ��N9<�Q��"⣪�.�އЪ��ӭ� j�8zPh;�#'u�ǳ!��É�E[P�Cӳ����#�WR�w{Xa���.�%����(sR�yE<Ÿ�py��;��吇��"�'�wi_��T:��ٶ��Pq7�'��b������-,�)盗�) ����$��o�TV!��G��������aZ�d�~BO3��]H^wb��&�\	�	F�㮗�+��I�ci��Q%�R�$�|	��c�P�;�l#�1��/��f���k�Ԡ�*��>"B�ghr"�⽸q�����
 �p�p�斈T��x�zf�8���⤨�F	G���:nH.M}�;E��#	�]�Rj!�S[����n���(m��8��m~P5��N�y�aGl&(��f��VӚ�3*��^�n.)r�Uq�)�LaY�n����1�=�]1.�^h����miH����>��<���7��)d%K�q����SK�����0?�ٛ�\K�W��P�q��S��^g�d�LL6=�>���l���3�1L�D2��Fud|���1�&�k����t8(�	�y.�w�5�A����"9�U~��=�:�����#2S#z
Ԁ`�/�"���k������EuE���eV99ਹ��837ʡP��0�+������0$	jH��� ��y>�Y�\��5� A1�5g�Ei�� ��]�L*7�f9�V� ��!��_ȟ1$>��vǸD�^+tl�H�e���$�����s0s�Ok�O"�EKZ������G�Z�B{|�|�Xi���]R��Wͤ*/��[�-ÜK;�����72vy �l�3>}Q�O�+�����b
�����D�<��o;��3�j�mK��$^J�+��K���͒;K��L�3�}y�c:���U �.&��+L�a��*02����)����̟}_45K$i�cG���`GI�n���W)�SO��.���	�Z{�Y_8N��~J��6�B���GJB��@���<聻k�g�`��W ��o���K�}`R;�$g��w�L#v5�Z���:Վ�v�w��H����K�
�k@�x�BJ��rNM0���f�^�j� �� P���j1d�`S��1�qxFi)����$����ĵ�)�Xy��vy/��*����������|�ЕWη��rDM�
�ϧDt��)��GS�Pi�3ކ�d��|�E허ȫ���z�,X�31�B*�W{NVh&o0�W��6�@�0j���J� �I	>���d9"lh6����"��&f���H��<-�>����� ��G��p�?�����U����jƍ�d6���֊x .}�_ׄ�r_�kM{�jb�{]����[�1S�m�3EKv��9p��3�5�[�A�)Ճ_���(z�ni��>�<ɑ�m�A� &B�|%"C�87�<�	|YXV{�<��9̾O���l*]��ԣ��/k(y�a.")JY�(56+�_)���"r#'}Q��p�f��m�p�CW<s"�ӦMe�y��!���x֫��VCb��z�@��>�r�C��*!�x���81��fl�Wؔ�4K����tPD�Z4��%<����LX�� ����"�-/��) ��|��K&���.�L�E;X}8��	�,��m���"�{"���P�7If�����OgI*y�֏��s��*���q2�P$Ա���~��m(5jzð�n�%N�!j4	�&3$k�7?��E�/�t�|���	�+���F�"_��Ã��}ص���we�uyhb^S�P	RQ�O��b�`mu�����< ���>a�^�p=�ެ���0&�A���B2��=��:���>�E0���ͫOӜ��CǞ�1jr2�����ϓ��ʅ^l�W�Y�Lyqk�3����܎�KH�+.��8%(�fg�[�&n���ug3�Δ׋����?�k�t5ݣnt�3�}޹�������F�]QI��X~�# j��P�x��$�B=�*�x`�d�T�,G���\�Ke��]���8U?�Y��X�\�L�ؖE�	0Y�u�7F��/P�4���g����&�-��"A�g>���i�s"ɳ|Fj�*��|dR�:\�{�<�v� BJ[��-'�*�:��&�Eλ��1!cY�Pi���8��1�
,;U9�:Eq����$}�5���6�X�I�x�#�Re�R4��G<��T|������e9�-�9 5J#X�/u�Y*C��c�Wa���'�c@�,R�x���m��\y���Jy��A�	���b�7]�(vXy	���p���h��=��]ES5wL�յ�c�~#S�N�(xr�g"[�#�\�,\�i��6&��lk�O��`�N9�j ��~.2L�?d.���ȯ�:Y�>K�	�l={[r�T�l���%��X%�k�dq�[����I���T�י��2�σ�������� sCSp�� d��g�g �[����-Kˇ!�[��~g�Fa�F�(��B^�K��l؎����I�Ҕr<J���\S��<��5ށ�.Z*+�!$M�G~�]�)J��u�5�a�x���d��btv�����5����.Zj9�����q�d��\w���o�͎����#���{�4�Y�sr�����`�[��Wd���JN޽�$`&{��(�Ϡ,�hZ�����3(�l����K�\�W�}������� �s�0	G�ZD�OM)���Vxp��'
z0��r����XBeE�����0Քu�_�"?N�P�K��fG�x�,'�5�Ob�ٚ.7�짚�/�9Ч��o�{r<DA|K�Q��^o���k-�X���e��4�f�P'(lCv�$���/��K������$��FI�p}|Z���fd�Iج��^ւ.�0١���SO��O
���.�/������J俘EÀKDA���<��K��ƒl_�v;�ي�>��m|���z|>��nql�*7�|�Ntm��פJJ��]�u�� �nt?i����J�2˻�* ~TS11���㛱�A�%=��nA�J�Z^��=�L��A�L���Gc��C�3��y����}N��Y�%�
Ye0�V�X�6I��2�/H�`A�Z�`V�t2��A�ee¤>�kc��C���s�� O�H0�C��%�u;e��TJv:��+�()��_���،Zf��s��g8A�ǻ�ϭ��m�j����iA���LOZ90�)���l��9-��Z��z�q�ƻ��ʷ�v��;TS��(DT��p�f=��%dw�.���.���]~�0K��<�g'��f���R�S4��Rg2h��3���7w{P��I�����w����M�׬��RlFLn�����@y�A�M�B���~hĴ��LH��/W�
�3����:��ã{pq����}1J* T�&v�Qa�%��(a�	���Q�T��$�R��z �0
�W�PW9��;�X|���"�+zqZy��)��t����*���������D��h�RKx�5]�t�Y���4Bj�*u��UQ����+^�
pc:�Aɾ�G.ꫲqe�WA^S�os'�6U��������R={�߲��f���l����t�F.�c��B��94���]����}�W�U��~lA���%�h[��r$B�?�?7�T㪧�8}B";wI���+�4�7L,)��I���Ն�L֕���5'����A{��E�%_)���i�@d�A^p-S�A;F�G�,ߜ�̾=���ݯA3��K�T8|�^��p��E��j=���c+�~������hNN�yiZ��Dv��ss���p��/�
@�'IJ>�'�y��(�z3ؓ�MG��?6;�<C9[�8�ӽ.�Z�v5��OM�Ӭo����i�;�)�K΂"���Xo��(�q��y���9.(�d]� �<'�t7��?�=���:��뭚%�����!���kx�a<A-Q;f0��{R�pnL��3�
V��Sd<�� 3;�y帍�u�-��*�m�{�`&�D���}�v~(��?=\jA��D��)3�-ua6�x�#���#��������!�GCM� �1<>R��Q ���e@*wD���:(�����{������~O�t����b��J�Q��;ݡ+�w=-�o;�>�tE�_��I�J��R��/�9�e;���=\ǽ��P�N�Y��v}J�����)�i�Ç�ȸ��"�j�&�����1�V��ϰ?U�}q�%@�fD�!	HZ�O	FsWS� �Ӛ���]��Z�D��S���F�6�7�لp(�c��F>����ݻ먏�V��L�_��T/,�(��
����Wt�˰z*8k.�F;4sw��"��!�?h`��ڟ��\�xr����׵��Y�!�/b� !�1Z� ��&)������d��^`�����0�N�"�N��>,�t��~Yik����&��/�\Y����y��@�E+�Z̰�J�:��1�Q���X>���{�ԡ�:E��/Ο��2��F����2���bʧ���o�~ɲM�8�od�{�g��{�띵�/��������L:;�+ "В�d�2g'"�j�@v2�z+��Mzb#�q���}4H��,��m�$F���|pB�;}h�q_<D������U����D� �G�Ԑ&S�nn�7�;C�9�`P���'z��8;7b?�7�-w����/"UT�nM�ٴ���^�tˮ-�����.Z Q��A��!��H�Rr�Ĉc�v/�2!=��ܝ:�Z�
�����j��2�$|���jws]�;�C�N2A�ǉr�NȓeiX���³;�gʵ���/����H3X&��&�p?���^�:r��^9��s4;�c����消��ZDTյ�&ˋ��;I �ed����O���=08��^1�)~�����B+,1��a�F���^䈙�_��1H�m����|X�����a`���p�pk����+�5K���
���� �,^��1�]�y)=�oq�R�g�;pw�R�c5��/2G�͠->6��_�d���u���LB/hm��<���KL$��>���\�������v���Iz<�e�tIrH������Q>��E��Ձ,h���Q"��|�(RQ�Z�3a���U6H��
*��u�A�j����/ELrm��M����tq��_Su'�m�圻}5�
Ǉ��+�R�Ť3Wd3C=j	��k�(UF���DMX�8�LaS�T���؝/,�j����>#F�m5P�X6�/��*l�w���Xw*w�A��Ǿޜ}��[�O��U�su/x� ��0@5p䉉P�T�%<=ɹ�0H3,�05���u}A��6�k�J�6II%#�����^�r�{4\_s�@1��likbe�������Y��'`/:�r��L�rU�U#��SPp���	@oH �_�c��$l�f�A��=|�� �S�`��jno�1�lJ�3��[�ޠ ��I�AW�`�; �$����%�p'{F� �����[��[z�֑��A}���+�2�{��䖬eM7��ע�%���3<Q7����Fmx�zˇ>���9�[P�>��I���'�&�q'xx}S'4َiK�]��f9ـ�B�3"��EħL����R���Oʕ�h\�/�����ix��SV�]]{.
������T������i���F{U����X��SsK�\cH�	�U@e\6籇�1Y9�����Ƚ��b����8��NgWQn��	P�|�=��ʭ���	������;1�0��	�$w0�r(�``������i�A�H;��Ɣ[��I�9�>��Fb{�V+�^;��D�]jzZ�����CE�'�*�c�6=��
{>'���ê'AL��CK��QYi�!d�׏�[J�~s�]�;(��%�r7��$M �HTg���A�������-��șnD�6�j�����=џl�gCen8U?�\���}��D�	~�EC�,9�yt#�s����J�e偁�P�v�34Q�����wEM�_�h��j���N~V׷�$.u���9��x��!��wmk*��׬%- �{)��o�[J벿�(ج�ZS�*$ I1�>,)�1�`tPC�Q�n��י�l)W[}u��/旋�'a9-R6�y��z��ASVi`(s��LO�L�M�ZnF�sHx"&�h�@�ח�:�� �j���5 ��k��l���$BTr�VN঑b����:x��������|[`�/�1%����/��BQ%�xzW4��7�4 ��ꋞ����_��7�X$�d�ԦpG_�5���)^�]��d�qj	a�Sf/�X�%�rɻ���ǧ��F&J{�T�ׅ%��e>��ik�<!��� ��������j��;X�*Gժ���5��^�[�"��\����r�e�����.��2���J;�_�A��K����D?�bs&��k����f����qC�ݞ2���SQ�Kp�� �	Z����8ǝ�zL=�bU`6��Ha���߉��}�F�u9\��XMH�B�A��Tl7��]!W��+��}��O9|�>d�8n2&�א�.�z} K�A��BdPUkf���]P̻!~�zG1Ǘ����';֡�!5����=�"|Mz*����]F�ޙw�����i��.a�a�y����i<�x|�}-���������Y_�|,��V�J ��
8�
ƒ��
6؃p�l̲��抲���u�%,�ߐ�n}!K{⹉��+�4�V�D���G�d�2������
���Z�����íl%�)�)��pm}jF�ǣ�u��P������M��w�-�����.5��b��T~��wP9���\tA�.X��u^������=�5�̈�&|5�&G�j�/��ϴn��To�a>��i�Ccn��'1琘$d��;U޾�b#���'@�4�v��@�^c@����k���`O�S���Z.�3�=h~�Ӽ�i��{�(v 8|�u�� �3�.�ڦ.�X��
�S&t��V���	��$pO޿%�w��<�o��#i@��,1j�(�]��[�a��!�n�](e[s�݂�v&�	\�&Og�9P`���vF3竀��!w8:5�ݸ�w����5�� �⏫HH�6�R�e��J���v�_�1`�x�'=�HjjR^��h<@�*�9�V/�*=4s�]�V7n���q�VkM���$���[��2<!�A>��h�����%���.3��܏����]Y�@M�~߶�Я���������\��a����wV�����h�)z�g����X�BF��~7=D�j'��6�;2�ҥ���UxLH}/�6kzmBX �^�*3u��{�_X��8��bׇ�%��v�fsM� S��Ȍ{z-<j(Mn�׵0��u�|�B��䳫)���'�X�@btm�L����^t�<�fk�� ���0�H"�Dp�Pf����ȎZ]�8���?���b�c���?9fQ5i��iJ�\m�����}U�k�U�How�׏*ٲ}x�L
�^�V�CZ�5/-��]��ve��Ĳ	JC�Σ&�I�*������"��~��_���~U�wj�;f��Hsť�2�}�u=�	�bi�P�A""�x�rё��D�E���ג/[�ʓ��n�A��w}4�῏��kA�,���s�+��`�N��!U�|[�v���}.e}�W�i�J4��6��h��18~��\�rc�1���>�?�A����LӕYNԤ�����Z�i�}� �zQԽ�����'t�9 �a�pW Ŗ��-_��^cF��o4�����<k�b�V��Wu9��$��{86��Q�{ˏ!1+c������ɚ)/[��~�e��~�&F�O[�[���1MY�q��-[%Z߉
�)pPV�)��V�.Q)���Fz(�\R�z�}�-�J>�����Y�&?�I��ؖoa��ɝ�p�I:��'���>v��5�;��qT2q3(�.u�c��>��u�p�I*�v�����SWiX8�4۲N��0�g8��
���� +�k(`di��5f�0��j������N��`.P���<�Q_�v�b���Uw�J)NMAxY�*��*Խ�K����jF����v��K��/��(;��I�ZOx���dKi�qxa||m�n�Z�zI`�m�Cjzp"Y�^��Y�O�?�A�<b�#h��W g^�M��u�g�$�afH�z:0k��B��ȸ���Lo��˾�m����gzY-��סT���l=T�]�pCqn6��p���6�n��Jt��P���4*��}�Ccr ����,0y���T����M�@N ��r$Β%�vd�� Q��7�;w��C�8�M���S2�s�O�^��X�h��b�ǒ��C�;L�%?3�T��U�^:�'.?:����U��m� zq�TV'�2�11޻&$x+�m��W{�~�s��?�Aγ�W�4�d�I���Z4���� hP���?Ր�U�F��	���.�����5QPV��.���-���g)Q�((=H6G�]�~�It�j��*��X4fx&��Y%u��V���pl3?��y|G�������Hv�
u���� Q���C���B�d|��m[�D�0�L�'���S�K�\w1JS������T�?��Ao,m �	0d3l��|��u#�'���Q�g�ߔ�BUĝ�X���흲����?�2�6�|��q���Ð(�4���a!���Gw�� iӜ�Z���k�&&�v��I�����^�2�c�/�M�6 �܊��ͩ}s��cjI�Փ����ƴ�n��4�{15�6j	���LH7]p��
D5�:�ё�QDK9Qv��&p: �HG��`���&H��`�\Y;a��&?�0�A
�4K+���j�Kl{O�W����zD�"A�J���u<d̑���k�݊Y�K�g��-�	�n�
o.��b-3rC�[q�Fq���u<v}���(t��m�'��R2z���}>Y��ѬQ����%�����8���t�`.�;d�-�	�S�A1��� ^��pX���"*���Ȟ�����q�O��=]�T�j^;L�Ǫ���V`�;����ˀ�o"��2+�JmvïwE��'�n��xM7^!�],p��d�^bn��6��h������"	E�D�~n�bx�'��?�W:��ک���3h�m3�����NN�2o7��
1jm2^[r211�Q�_���X�x��B_�H
�x� z)q!c�$�����|����q �	Hz��B���z�}�~�*��,k�u]��UL�\�Pĝ6ї�o�O�<�5�����-&�{���� y�+�ۃ�]��0p;�7��C�wQQ��y>�{�v	SqN���P.B[�b�88O��6�\�V����ʴ����(Sj���d���dfO�o��Hfrp�m�rs�k ]a��Ӱ�{R�]"2�O������3���VfrT�"8�*�'���b�8U�'�*q�d�;��J䆋��T���.���rj���H��PO�%(���)
�#��z.\w���$�(M����>~=2�h��c��7.�S�� �^A�:�x��W�c�I�3�$T�v߃��-�Qd8M�:?A�^h���wc��i�=���u0 �'�|��j���0,7U�\���#��wdu(��B��'�ݍ�X�u[ci�荲�I��r��$O���O�������,W}8)ƪ�݉����k�$q�������im�q&U�Z?��Q��1B��3��T�	�������U�D��j�Æ��+FO˪=����b�oM7^i$7������P�y�Ƈ'������ށ,|"�<�9�j�`���g��(4�"AAAtь�E��z�~4k�H��ԶL)1�H�v�1��5��v%�QyO]6�{ ӵ_���I�0��!��#��v�<�<�[��N�A�>ˤD</�������[�]Bt�T�$�=Я�u�v�u>�tc�bw�?͎#��D�xj�'��Ve����F����)��2*�҇��X�sA�J���k�
�	�;�ϭǥ+��:�-�����k<�Z�']�L���_�������MnK2Ij��K����H`��ۮ֣E��Uaό^K�V����b���n�1.:�I'�h{��Ei����J+M�
Tcc�;|̚G̗!Y��}8�G�����s*� k��2ҽ5�@��O3c���yB�T5�1������ �ʅ��Rp���Ů6w��Q6�02_�'
��y��X���Zb�)�*��y����rZ���/1�p����>��F�8��f�9�R�Tl��3nNvA` o&�A4�n�e���D��҄���z5�Yi)���/M@��z�%�?�C�ـ�-f��Ã7EH�j����+�i�B�"�|�>_�
s�v�����lY�CJ�ia�C<�S��]��\���%꾽��spCȜ����kz��p�EάC�)yk���vP%	V䈞I���G3��n�ađ��Xܮ���(��6������wh�S�N��*�=,q-�='�l����B��U�*<�A}(�Т�%Q�[7��O�X�_��Ua���iҒy5]�A�R��3*�1�B�ɞD�x}��iR�H-���t@�M�Ќ���4�>�k{?#&��IឆOb.�̧�̩�ɛ�||�e^������[M��0ݙ���BC�9��f��[Ԗ{{<)?o�����uOZs��Q�Q�o^>Y�
�bV��ϼ|v����C�>�wSv��.FG�.�4�Fz�_����ڨ2�W�؇�0$�ީ���sd��ʆ��gix��Ŀ�m�L�m��Eѡ�>�c�r��/�-
A�A���dœ�r�a���m���,�VW�;S�w�e�>zrs�ߑ^��b9�5��U̒���l���*-.VU-��Ƹ�/���.��k�ȏ�~
o�<�'����5`��<7�K(Y�W�H�oM�A��V#���<�W<�tU����sQ,���p� za��`)���X"}�ޤ��N��j�8������Pl�,�-T;P�}���gi�&�&pL*�b4��. D�N�m�+������K���!4���O�q��+��d���k�I�jt�d�u�>�]�uC�]+�稩�����0'�;l� 64+]w�Ι�/	����_3����A�������l�T�v��|�C��!�/�U��__�@�9�j!!�4B��|�0��r�/�6��q��?��׌�lq�Y�CS/K���G�p��=�-!�tS]�w!Ϫw�u��f�|̨ �,��)�۫�������+Q�j�����&�hL(6~��N�O�t�����ߑ��j�2��N�+V	��w��8���B�cX\�7�7�`&�Q6����e6���-�(������!���$l򢆆�u�3/Yz\���Ɯ��(�mp��~z79O���>��N��&
��>�y�qga�����0nk�C��rn���'�	��vVN�rbh��R���C��U	����93��w��g'��`�Ŧ�0��[_�H~]�_8hq�]X^ׇ���K�]o�a��7��!,f���Q�芾�P�_ ��>V��S����Tn�߄����S��������eL��W�z������9�J!����@��;���M簾���g���Bj�υ�U��F��yn5!�r�{�HM$���|�w�����n�9����$��q�H���C�ޞz����{�N6Ay)�(�֠������
(���^H������-��(9A����?0���~� ��Hp��H�@��7Q�6lR�8��W�%��S���z�s��kߪ7��%�g��҇"���q����~�<�6��{XR[e�C��c���^��:�Ƭy9�9�Xg����'��R���q�N��8|J8�^��u���K(z��!%2�#��+ݛknk��$ &0"�`���8�yt�=�<T�M��uĥm��
�Yg������9l�a2�^|7ߚd������tRTӛ8��R*6�fȢ��O�Gi�J���Rf�N�!鑑� �$����Z<�v���b4��^#�E_�r��!X���|a�X��o��y�KG�18ƄV��g N/�E�8��-x\b��ĥ���bu��q�#�c���:����q��b���:w��Qe���v��L��QP^iߍܱmi8�x{�V�X]�@Q���fI�Mb��V��G~��t�ǁ��xc���*�р�;N0�]�	��w�_�B�/+1hq�K;�嚄v��pe�`��]�{;�����'�K0K����-g��h��f�5Ӓ��n�iJ3;O�c�X�^�xL|3y>��z.��Ѣ��r�"�Q2�8&�g�EՒ8��g�����w���@�J������hޮ\���_/�����08u8}	��C�_�t�4h�
���й�p���	z:�rj�&�k+��q���y�o{��k�9n�r���v�,1Xò��o�U�o�c}�$����/I
��Ц�?�X;g6N4���D;v�5�b�ӓO��{�L���Z�^Q�����E���j,���!���E=���#�	�}"o�HƮe���Լ�9f�/�
)�4c[�J2L���34�Y�i�f1��6�`�IO��	���N��ʄ��{X`��f�%��@U���N=d n��W���jn��Y�X0^χ��*�S�U��,����+�~���ijx*�eiK���( ^���l�9�-R��{����I)��l�0@�t�C����m�{���(��BD��J(��.q}_M��C3�<=��(
�������Y�a)d/�m��~m�Qo�*H�Q"�t
��h��ΗȉB���637��-�%�y���Z�	��h!~>���$C���È��Q���ߓ@5��}b���g�<�k���V�w'���ﵫ���T�:���uo�v?���Һ�����ОԊ����xW�(��׍	�t=�fd��:n\3���t����$�!C�@	a��he�"	���ah0T-l7���IY���A��]萈���󷇷w�m��}��=�*1D��(�be��0�H��r�I�Z/� ��L~�I�]M���Z�'�<+`��M>ƹ�9d�.�S��֛�Q�96G��3�y:��+�`�ؗ>���J��~�s���s*��qy&��>ܢ���D�J�� �`���E�zf��9��3=�B��������-fmV9}�2������^�t��������Hqh��B�[�^G���)|���V���%$�Q��6�|�v�hI��YUyָb��p���W�V�n���^<㢽�w.�.8�y��`����%��L����l���n�փaYg¢"̚!�+��u_���A���������,-���ivN�~a8�����x�K(U=�ٓ��T4$�+`&�Ք�je��nM=-f�7x���<o�i���d�b�F��A�=,��/��Y)��w�CgR���s�j��~ZEj��4@%Pw��7$��l�	8N`pq�9Bto��ڥ�,�(G�����w�Z��Gz���@UJ�c��NH=��IW��L(U�X�m����\D%����K~�x0o�!�8^�dvbݍ�jrm����]�� wEV�g@��QoRh�v���UL��o3)fB���e���~A�|䍶�e ��2��7'��I�l����-e��(��mN����o-.h<	[0L����U�Ø�e�
���uW���}��8�SI,�j�.=�8�l7�b�5� G-Z��z�"j��"}:Uք�(��6�RB��}0e���iAp��o�� �s��b�o��!+�����7��\
�t��#`�,5��� "��� 1����&,	}���������ۍо�>�o��l�@k�����Ȑ�ኃ����*	�/�ԓ�I���"���,�ã3c��HZO��������u�Na'_��0S.`'��Ū4��;��
%(g�31�n�{3��5`���Ru���Z�d������f�E��3(${v?F��>�rG@੆Ώ����7����G������M�OLY��r^!�OEK2�ي�F���0-���ry;]"�,�iU�h'���(�I����+h!i�V>����b�	%ߩUul%0[�:�%M���AfQ������x!w�}�j����������j�c:�L���D�(�oE����%|E�����>�<ǚ���׆�?��p��������u��|�O�����C������F�=Ɨb\W�?}��8�R��d���VI��ܐ=x�{�U]�R;_&emX��-[%d�}+O�3sb-���s/�S^t���8�iuqZpEbX.����w��ʹ��[��$�?mʁ]�N�ӽmhSGQ=���J�?�֪Wm'����e���[�!�Sǭ�of�:_�`A�b���i�k]Rƨ�q~%.�bPKkì�j������xU��t���"0��Wd��緜!ٕG�VR:��D?d5O�hө�L�O��Ȼχ� >�&�7�`���H]m��{�����b���w���%�
MM��V��B�ߓ�ޚ���C��2e<���*�A����ԋ�K��xK�K�K@�5p�^���\0D�#��G�O����ph9a��1�ץ�#�1��; :)"��w�l������1�����Phz�nl1�ۋ�F�>qy-��R�'�4"�2$ͶǢ� ���� �fl��#��c�@�Yod�-� ,���{��By���a+�| bo�/t�Bʯ��i�@Xn����O�k�`��'Lǜ�B��u�v����S�h�����'�;��B�e�� ��e0���o���}����t:�` ��3��}>����:7-��|m�BЂ�}�fg��jڄ�m�P�b��zt���񳢢��5�Ǎ���M�톄�R���ٻKï �����̄�������ac;�0��bk͞
�F�1���7|׼U��b'�'v�Q��E9�9sy�BH��.����|?�7�L%ij��8�E�Ϥ�y,�1q�Bt�c�=��p{l����	h5��+>봥Q*N��^Ҹ�dQ�QDk�] �1G�h'
�D�նJw�}�8A}�^�(~�8��m���9��,�[ɼۄ4���V���?��.�h��l,(qo ���![3����̰9F��;��)��_�^n�^6>?,��:��}[}�ɞ��e{����Lp�)�.�L��2�w5=ȏ�ث*���\������������n�q�3VA���V�g+��YP��L��)�,��S���}�b�Hk�{��5� ��ҁ�`�+?d�#bN�����_m���� Ir��ZIbK��[JE�cWʳ9s�f��\;�����%���m���!  ����%�lLE�/Zo Z.d''��:�9��X� �S���q�o�:ޗ)��W&8J���Tw�������r�6�p]_���sר�3שz�>���k������0+��W��|���iLQ��po�����xˡbG�H9ɟv�u+k�nh�*�8)3D��/#��ƭ��oˢ
�}׽\ŭ�'mɰ҆�)w,t��X��)���ސ�	:[���Q����p6x6�>1W������]���L���S� �D�E��T�AEģ��l���m�O����ćU�7A�����Z��FY5l@ͦk�V�#ax��D�)��hcli��T�wH�v3�@V�Y�k��--�o�Sx����%u0��66���Ƿ=\3��r-.֡�Zf��E8R;��H�d�Ӯ0�y�!����M���PU��8����<z�QQ�|7M�د�^��C�n���y��[�`� g���qK��%���B��&N�,#؇o>��P>�b��h̳Lw]�-�]b�Q�#F�x�7�Ԇ���c��6����"3�م$�q�N]J�����8�N��~�^K�yv�t�g���KC#iC�3�y���|�~�T#s��1xds%��vͮ4�DI�y�f~�k��Տ��3�uS��p�4C���n���,���C"V�;py���gU��~;��J��1-}��ru	�Fs��TA��r�'�x:���Z��EN�7�t�Zג#�� :�rf߸��"i]���i��.3"[�vv��k����ZPbH<�����Hn�^sŞ��v3��"~�NbW�W���fY�ʟ*�[&5�*��]�MC� L_�m��2V�簙L���}>���&C��brk����c*kڃ��^6�|8g�E7�8 -ڮ��*û9�c��y�W(�@�1:�����QE��M�i$��"�U)��v%��G��b5&��6~�1��.�4ö�{}!��88���e	�[p2�W'�"�v?�Jq"Q.�ٚ|?��V� ,��S��ڈ��p��[q�7G�I��x6V�^�DGB������L���6���Y_��@`��S��I!W��Ǫ܆I�x��儦p!�S��q��a�����B �Yk��S���ZJ��@����K��p�.{�	K�(�
;�S9�	� �*6�;��+H�_<�r]��;<;���-�n�i�{MX���w)��o�&�nϓ�zP��u� �G���ꤔ������kq���4W����i�_[��-,]��hb�w�:�����qH۲�7�1�����WSO��O�%��V�?%�Z�,�-��._G����E:O��/x/E�Z��WI�Mg���L�:a�n�\$�����<��^�L�p�L$g�k9��=��1�������!�#�-/q��0�V����[O�(y��)�UIu��^ʦ9�ߺ�쟋����=�;�������MU�ެ���ASi��ÿ��.��av���8�����cw�{�2�Wi��/�X�ݺh�[�y�F?�<x��85V��-�c:)�}����o���$Z���CCa$��^�\h]�Ė�| �a��!�%#vF6*���$��C��%�s��9������L~-]�Zo����x.InU���s�X�����7Q�9�N�e�;��{��ڌ�YK]��pqJ>�fu��T+��_����S���'T}���� �<�4 n�����1��S��!�d3��L1H����,�{�����
$�7��E�8��T��B=��{�����I{��z�G�A8�� g�#v��^�j��Y=� �~�kcY�����
}`�i�7�~=
�VH������R�+���%�Xo�gt���
q
�����?��T�?(�C*���/�Mi4�Q򬶠p�N�D%�>7	�k���hd�|��
�yQO�����@�H�%���/lp��nZ���
#�!D�.���O����/���ś9�~�ˀ�+އw�i�0ue)e�Y�g0�����!�e��gm죾�j�ͻA4s)��c�����{���3�v�����p�y7-�����.EW���Mǭ��,B#�wٔ���Ѷv5:��=�%n탭�z84)�� �~�g�>r,ޚ.yg��Y��ϧY/�S=�݊�%�@�96�8�8hۊ��+&�n�k�C$������f5�2���;�7fҰr��!mϞ^Ϫ���ژu�k#��z��H	��8�	2�}i���)��中�7�@��d���>��݌�*�����0���Zw�����sN��?[g�?�f_��!��o������wÞ�D�����1g%a�;>Pі`�����I�2a�������3k��D����2>y�}yp"&�y���W�aܷ��ަ7A��y�w�XP��)7o[a���j��X��w��N��a!����%�=�FI��Ϝ葲&�mh�X"����j�����Ut�E�Xɳ�����s/�������~�{�N���S	N�KB�[]ŵq�U�@?����+!Kڐ�<}�$����D�1����@���K�*cj�T�7<����n���@�Si���L�R���B䣺V6]�55�t��l��9�z��Ŷ��z#���,�;�TRּ�����۬t�km�if��H�)$õ���� o"T�S�o^=8�~���hӍ�irHBx:�\|���\���h���E�.���a��,�` ��C�pP�+��w�\��VT��\IJ��h����ݽAzJI�qN��V�\^�:5K�k:�`�Z>��4\���׳Dd���f��R6�{~>�Y��q��G�����AN���k$"�\�xm��툷��Bn�j�p��˼�.5�����ň6��~5h�~W�K"��ZԆt���s�6K�ꐠ��d�{�e�禩��a��3�Fa��R6��9�n�,>��^{��K޲�:��������T5�U���u��Z�8���sUe8>&�d;+���P��*t��2]�GuX'X����UhӘ��c[��W�ק���Ѯ��4PaM�K���i�� ���uW%���a��4�w��r�q��'(�L�I��a�vЇ�亷�4�ig��޸ċ��m�7+���5Ť�p�����2�m&�5WC��e�g�5�_�����ÿcH�#�
�Ż�!��.�,��S�6��{U�慤<�ц�?F����������+G}i���#9�M+���������^�_�]+�?�HwE�'1 D@%UR�)�r�x� �=؝��[������H$�U�ڟ>"�xq�$��*$��f�z�⡜��݈#o�"����q�T�ޯ�������a��@F�\:t����2��Nipz��U����v�	��L�"�.:����uc̒Thpy�O�t9։��E�e����0|x^VL�1� )�˓j��ܰ�5�¯��1�	U�˼���Rb%~��"׶R��6����F����ݲm��
�����i����M/����d&y/nk����n�0r~l�f0����-Y��~�'k���~*����������O@��x���y�`	�?"��8�u���r�؅>cu�+�r����������"_�\�ބ��&��r�m��!�.��k���v��o�P�A����ǖ��q�n�n�J�
,��bG�O�=W�V4���y�KݣA���QOL�I�Jf�0�����\�-{6���%����,���eS����O0�������(�7�b������e=�3�M
>��#�B'��y<��6������6��Sh��f�6����NL%h���b�OB����ȵ6�T\�F��ܳ��/�S�}���R�E�7�a�߃8��Hz�4��� ��z�N���c��]x��l�q:y"�����F�姝Ucw���,�����"�jdm��G<O�,����EDɎ�!�m"W�;1i[��-[P�i�0E�lA�vɇ �"��L1]~�p�
O '�\���2z���Ζ�lv�r�˫@^\_Mreh}���F�Wn��ߗ��?��<?wB�ki��_�kMJLtz�݇'#�ڶ���)=6|���j�y�p�4�M����P����&�|�댳�<���5�2���hѩ���ol^E�e��O����]�Lb6E��Ĺ5*���U�~n�oo	�A� ��l�/��m)�:�\��)Ei�X.��hG��
�P���6�9��kYނ��{C*C_��_�e�LP��ڰ�>�5�6f��=H?�	i`�ڭJBa^�0��]v��J�-�s������f���-R�*[/<<4*O���.Ń�0B˾���3��6E��8��'�e�m��5����%��&g����������OH�$N
'�<��$�����i�� �� UWS�ĦV�up��zѤ.���?�t��6wwW
�_6��'����sN��ʜ���VNZy��	Jn�/�??�8�]
�r�M�epμ�Y������1G���H�GiV�rG$���`P�S/��Q�/L^a�o�����nԀ��y���7�<���7_�+/�$��uy�(iA��zX�c׻�v�y���N�����~5��=�6]1}q�%��F��x��(a!���Ͱ�!W�A]��!�q�ULK��+�