��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��e�A�����������*�65`ϧha]|�fcJ3���#c����:��*d,!�u=�����>���k9F���D�ܻL�l;��z5+*�$?Zq����t^_y����ml���{#��L��"_�ѷ������L=
�&�8E\41������_�}�Re~�_�!��ȶ�5��AzE AK�%I��XT2�t2���#[h��i@�
ò�yF"^��D�6���,����5�I��\%$ł(����W<�!n�x0h�� �ۢ@|�g.��č�fbI���y4Ǭ�~�De��>A�J�+$H����ηַ&z&vJ����%���o/����k��|�Qe:�z���1����Z��4����T zG���݊@�A�}��N�}~ȵ�=�m
H��G��OU�+B�p��yH�'�k>?����, �ۮ:�)ϋ2[�}XN�@w%�l�K+�N��=ܑ�7ں$��m��/X�*����U� Gjx)*�f=��2���n�BpF(�G�@�{��W�q�o)��c ���QEx���QH��p�x��g$5�D:چ�Tc��;❓χm���'�a�3���HK!Q&�,�������{+Ճ�Y��?��sm����H9����ɠ
I�����c&�U�_�:��e�� �A��G=�o=�ZIK''Z�j<4���m5����	���X��'8Mf�uXV���3��[G���tl�3��C�ʼ�q�Wd�kCϨ�T��,���G�T�b�-��؅��LH���fTI��	n�v��IG�Ul�	䄘�I����VU/��6B�����@�֭�)}X�*��0v�^�Yho�l�θ����
~~�k2�Œ��*"���|KpD��;2Fw�$f HFK�2bX]�d�X��5�T�>1lco��K@�^C��*r^_��g��]������+p��߻.h\Myr���8۬�����kWfeq�F�J�G��h�P.�iV�k�"̱(
���0�Ai:j�ʦ��+�Qx��j����*�kض_8+2�{�V*�`Oa޾�W��\���_�qp�ф�w,ŭ	���bĽO��aH�P�3�{��rU}�5?�)��Ҹ'��Z�]�u���b���Y5�?ڷj�X�fkVܓ�'�jݩ�Mv�'�� R1-�����l-|s���f���lvbE�?�}(|���.��ʥ�>�'����&�.�L#u�
3l)����� -�C&�j��vF��nB?�, ��;��@NR���,6�%Ŧ��N����:W�G�ǈ�8�և����A�랕vɚ	�P�G����O���%��i��>t.oi�Si�;����So�{��%�Gq*p���Ov.��"6��
NM���k-Z�	H\�)
��{�v�$��$� �ʧ���H�律�:��-�"9%�����}�
����5Y�( R/�	��a�L��a��%��Ԓ	j�n�fnh�6��aO�-����BoTX��9ڴ�sP�ͤKq���k��^�4��� ��� E� �������|���iN��b�4%��E��Cq�C��h���fs�3=٧��i�R��v�A]k�v��4e���B��^o<Yg:e6��A��O�=��8w7rYZy�Kh��n��GB/�`m��l/T�ə����އP�MpƩ.��-��LfFQ����hs�!W�$��W﹀v�Р�fl6i�'0��\�3��a�{j�ZW���`fV0�-	������#��l�h�������n;��1���G��ΰ�KQ��ύ%TI���W��<�?��Dx��n�1�x��;�������g�G���ꗟ�[��hn��&F0���)T���������&«E���"߰N(O��[q�JP��N}Ӽ[���&b�caHj2�|^��ch�S9}FMdG)�a�-n�ѿ�O�m��X�,?�4�isw�㍯V}���B�w8�~HT����U%%��Wk�LT�b���v����v�nf)b�GW�2(s�]�NF;�Z͙�w���q�KҤ�$��:`�"J�l�����c�m����_bg��+x�꧛�R�����󅍎ڳ����j?ƜEg%[�4�͌��Cǵ�&�Q�$�q!���p�e���T�KU�P6���,u2�˥*�i��(`QXG���
@v�n��ͅ�R�.r(b��a�����=�^�	\aY�Ct�J��^�i�&�Jn�{��la1�I?�Í�ϊp�#+	�[�_af|$1�������b��HP�P���^=[���"�Z�:�3�f|Ë��$)����n�W��g"G�l@:�(�% �]�&ނ��e�`�l�P	������u�͈�	�Ҷ��WzyyA�Q�y���b�]wJk~�r�Y�� ��}�$���ϣ� ����.��*˭�]� �e��ZL���T[��[4z6q�)ț�&��2�S�_%��Q�/�6�`9�}�z��W�,�� L���ֈ�xC���xJSf ��_���
��$*�4�>]�#�<!qq�vÝ���b�p��.Jp���yzV�^��K�~�����O7ܣɥD�5I�k��hc� t��E� s�����D�Lf��!�B��S:�;݃a�+mL'�{T�4r����|glЭ�?��͈_�k��R;i���:c�O�x�Y�M=3�U��'�2��c�j�^��O�rg��S�Վ	I��j�CWa�.�z�gR�����t�9�"�ZH|&XJ�s=߀�@�6�`��m^j@��΀�Iݸv�.�D��(P%̇ �J{��MMӕ�[�7h>]�)ݩ}*T���� r�@��$�Y?�t��/�͈Rb [FQ�k!�VZQ�@K��x�oȭ�J�E�{<H ҒfC޺�y�j3����($��Ry��Z��P��������q�Gv�4��^��`��r�9�7t�6��4<��U�h�����o!]� �̢��=	D�/_v�~��I��y����T�e�"d����0���,&�o�ص��C���}_Ġ��?��H�&���e,�޴�Buu�.mĀ�f�m���� �@!�A<�@��m'�F���l flQ=��>�Q��j�F��̞.���Z���Z�lǍ�`,�\��R�z�9���Qš�{��$���]�M΅�S���,��t���F�nԺ/����F^�Z�޾��o~�9��-����j���[i+B��
,HL��\��&���j~����ȟ��%S!7!��u��{t�|�J���韇�	i���x	1
�\p�H��s)���ϛ)CE�V�'��ū$��#�2۹kI���*y��g�gD��LTR��c|�-��}�؄zg����8���v}�5���5��}��}��E ����x}!�ʯI۹e�j�g��:r�ǺW���k�R���f�<�l����P"a��������ſ �)�?s��eEY��x1ך�k�	�1Ia�9Ζ��y��H�W�Z �M�~�W�$��x�]�H�~d?�A��6�h�Rj�I�j����@�l*O�O�s��~�G߸�s�ե�c>���;��KK����!���3��m�����^�˭��:���
�j?+�&��-�,6�l�݌C�')�eP\�@̂�О>� ��ޣ�v|G�)��K-	�yHg��O�Z,�[ԙ~{�G:p!o�-���$�I�NĠ	�un��+�5��c$	�Wy[�*�@pƔ�zy�$������}<3I��+��;�8o5mXl:�����[�p�&�����gɜ{�蛱�F0Z+�bn&�+SV����fx��W]��dFVx�1������z��b9�
�Ex��zg��h.��	��yM>�\X���h;C��3R7+���R?��u���V�o��N*��I/'�@$=��O@F/�`�Idho��o7�����i�$��m��l����e���fv�.��A�`�ݵ�ۡ6�Sh6�6��!�X�f���s
�p�36g�ĩ�.��$�[�LA�&(���a.�6i�A�<�C�K��@o������N�_ :��K��( _�w*`M�\�t���R��.�ɐf�yp�w�4Ĥ����Y���*���[7�=.��E���
������*�T|8�<������QX/UB�#޾1��꟣� Sh��?�G�X^����bA!����l�1���=�Wvg"�q�s:�X*�6��e��\£WNY"��7(:L����g�46^kB�[},��̔4Z#� ����:4;.�i�G[y�zߙ����UÉu�iD�lY���*��8�O⹙�76�th�dq%J�������r}N�F+�\��&�|ǆ�-�q��O��_$�V~���ۗ�J����n���M��-�77�NT�һ�r6��y?L�g����P1ki �>p��D�������DE�b�
>ʵ]����Go�C��з�l4�1gD�[���@�W{N�z��I��[[v���G�k��=Z��1u���q���:υ��k�h�N����K�CX$t�4t�c,Γ�����6T+�/�_�ܝ����1��ǵ�m	U�f3Uܼ�1�lyC5a9uL���hc6x9��q��D�ԅ�Uo�kN�8�����^og�Px�-���Ƴ>��p\� �w܂�g�a'�׻�ҟ��얦,�C�#�9{�{,z�w�5���#�@J8�E��S #,A�)����^�zS�����)�s���2�/��w-5-Ы�_�܄�E�W�ך:j�3�~�PJ�Z>�QY�����>g��Z=�H��q��E������ē9�κ�  �Z2
8` �*�:U�bq�祊�%$`�:���K�Hq�ccM�G��o�DRv�l�?8K�>�m���/��E�I�_W\$D�B+�>37;�)3$[9�&<[ 9ڢ=#a����B������r���+Ɓ�XV@�Ф�9'�׾Q.���=�[��=��'�T��̓ �|B"iJ��U�@	���Ѫ�5O��x���K�[=W�0>Nږ�!h�;æE~k����F{F�-XKZS�Nx2�TԌۻ%���㺭%ي��T��i��*�ͽ�hS�k�¶&b���+��s	��VyG�~%��	����gU\����E-B��D���M�)�)m�ݿۿ���):�l`�����|����剭�.y�������.g��frK�R@S