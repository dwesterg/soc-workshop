��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t��m�O'���z�p�Q���;�P�ӱ�����[�kA��h��{���f�]n�W��E�E�5J*+|��\0�f�?|��v�,�<�j��ls&�u�A������}�n�/�$���f0�܁\H .J�.d�L�뙭𺪛G85���ۿ�<>�셤�D=l�@'hkJd���<�kݽW��?딘���ǯ�Ps�5:���Y��k����ik9�z�tr4�	��9���\��Q7�5L �M5�M�]�H���.K�$�A�#h�X�p�n	���5&M�Ѻ����ؑE�S��:�u��	��#\���͇틖�i� }�n�B![M��o�!�6����Y���e���W�����7�v�g!�io����IGݗ�k�$Ī߾ ��>��K����:��J:��eK�(�esW��N�Z�j��f�I!d���䪋�S[���O�-�'���Z�yv��p5_�8&�"�.?҉��aZ�{���@JU^'��B�m����J���*�&�u!�r2��v�ӳ�ɮțVp�� ��T���
@ֹ�����/��ۑ^	��l��;>�x�B!n.+4�]�A���v��W��F pN�n�Kk`��d<���"8�wvh��i������z�n�h@;*F���:ui��c�MW���C��Ǚ���	�����8�H��53�XC�z���$q�
�?.76���E����4M��A�3��F˽�6��~7�v56�Ex�0e:�M�˟T$�
�k� WV���5�k�L�jjI?^W�?���J��ť��g~:ǘ�>�)���b%D�`��	@���-��s����d)���P�g�ϱő�S��.���9����J�rD0�	G�!�0�ܬ���	{G��,���\?�5��z�6�X?�>��j��8�Re�.�2��̬����Q�����]������U�_�)�SJ���|SIO�!ַ�2̦]�9�K?�n���f��l@�	�3�}�A4�DƔ����?V9�I�/O݆��k�of+S���_m����[��M�M=��o�����Z5��e��V�l�\S��ƁI~������֙��\�>{�(2��Ɉ2�?]#倴1t�sB��՛N�;D9��X�y�K�o��X��F:f���qQ}�n�J�ɲ����`� [��Z���7k�?"��̓�RI?��;5 f�<6,��p�N�:zR�xQPP�`L��cr�y��Q�+���&�����@IBa%�4~�?�r�-f��f�z6ٯ���^IwfD{��.�;��ɏ�?�K�9x��v^�&��ܬ
�lDTlR�}�l��}�w�D ���7`C�sw��<�� �!�����賶y/B&6�Kg��Y����o�vj�o�cǰI�E^;�!�8��{*��=�g.���F��e�稗���>�)�/܋���{_��+~G��0�n[n�c��iI5|����ǉ3+�ʉ� ��KB�X� ��e[X/��I|�D�A�Qز���]��B݈I��̧�.�K���4���NL��CF��P�2����Y	�k|�]~���=�j,}�n����O�Gz�e�$0�O�y�n��M-Q�\`�-�ߏ� o�.�1ɸj�����p�#q����`��a~�O��g�,�����̥�ϣ���)��tºp7�k5��{2�*��M:_���y_ l�����I�9j��'tU�H����~l(�	a�iB�#^ʠ���֓�Yp����E�,z����<�Ocu��쥀��>
|�����`��	���!U!l�W!�gc�Ri�a��wY�����zkH�rFB�d�+�yǒ�y�ܧ= �����gg^NW�1X�!V������o}�|={!�w�(p�Tf�6ǟP����r��g��m����Μ�@=���1�(�^_�9�X�L��E2�t�hkɦ��ɒ󑍮v�o���	U���J��C�?˝a�p%�$�m�e��;�1}����M�����5��@�Y�޼�3����Qq���¯����T�,/D	aw��K�@�㹦���#�a�T�<?����l:��*p܀�
��]��'R̸$SsZ�������2�{�
 ]�2d[��v�<'��i+��q5�V������E�7D�K�/��T@�r�N���������Luo�)&���(�k�Ѯ�/��T�;�M=B�c��/�,����f��'�W�:5�7&���c4�KG��}�6�G�]�F��#�-�����@��q,�Z0�=��~�1ed9�Mo�1�4age%1��|��1��T���E�)��x��{�� �ޚ�G^涥��F>���S��}��׾J\?�4U���G2�-:`�l/���5q-�[�����Ol�lݝԦ�2��w�B�_f�e;_���Y,vs�
�|N���1�F|�p~�?�L`�wԧ�����N%�f��C�G��o��zs?MeO�:d
��O�f≔w������N��R�;�<B�����8���*,1��������c�X��c��T���| ��L�|UW"���&��w�y,LG�CW�F�u�"�)�G*aA�h��6�CZ2�vj�T�旿A�9�M2�d�'hg�/Y����NN�g6�Jt�c������ޑ�1yQ��g7�+�U|:�����������ú��)h� �C`�����b��RS^V���r�Ȇ�!¹̺�h�h�o�(�#[�-�дn�0��³?቏��d��Bۑ&:j�SG�ݻ���I&���2�J���Ks7Y&��I?GO��n��(N�a@�[���
���:|�q���乵7O:"St$���c�SYٽ�U5�9�'��W����=�^")evJ�r�)��;���D&�-�R��l1�t2a��'�QC�����qT�sv��^)16��*4|"��A���(�3��~�)�C������X��Φ�Eht>��l͟�,�s���ӫ�"c��x�U�nVm
+��F3<��F�?�|����^��!R_�A �a��ǵl�W��,�B2���[��Oԗ���t��?��4��\˴S�J��s��Y�c������u:�k�9�0�#:��-J�BÄ>�;�!�T�Z!��������f�PQz�!;rۘ"ʇ�����7���^=��ҹ2� ��K7���	/�Y��0����/Br}�o���k-�����?7Cg[�6D�Lgꎖ~�I�b�J�d��q.Y��h�S���s�ܲ�,u�I.�I;꒢�IOm�3��#�]�M����"&�eW<�v��!����JI��K�x��Ǥ���v[R�򻀠��E��eĨ�־��mή��� y	m��?P����,��sh~!�_������*��9tq�������;_w� �X%��>��,��':�m����>(2��ĳ�V*�[I�w���GB8�C��O��7PѦ̋.�4��?��=��v3�ǒQ�$��d��U�jL6K��[��H�����w��!��,$��sp$�8>7�_}��1c@�����J�J���K�қ��� ���M�yHT{ �����ȧu�ظ�:v���֭�����3�(nF����zh����Obς�x�j���D�T��W2�B\��J���>��_�p�Hl��Z�~�W�aF4a�|�U"�G�����ٝ�)�t���P�jH~~��z���c܆s|yp�&8{�8�������D]f��1�Xz�4�ǿ7ն~���γxlz1��lv�n/zUK?ӈ8��x�7�Ɉ��ux�md���ȷx���n�N���dP%��zd̚qc ��_��j�W�yX���?�?����\�@v�P�-�O��a|�5_p�%����=��[_���	K�P�;��j~=���y��@�l6�jC���߆��+v�+��>R]�u����ۉ z�U���j�~N�WF{5�W-��Hm`�i$��y�����e���~ոs����z���7_�y�ˇP�Vz�,fܨ����
Cub�d]2����������J��t���EP:2!'A�x9G&A�"����I�3�q�_0\�\�d��-�^6nA�����.�Q�C����MzA���i��L_��c_|pz]7���>�Z=9�!֏��}{�	|�~&׷ kR,<��j�魍V�>9F�|1O֦�uuB�$th��r�@���o*<�&Zh^�}����
�Z������saç�8�έ
9���qp�L����[M�kW�7��M�����BTL�D?
`À�2���sQ��
�����#�i����%�X=��o�]U����#��h2�N��Q$�f����|�����5��-$�9�{�:��C��,����6�3�О]+��:����k���if����.E�NǗ�a%�[�H�l8���?v�A���y�������ci�
S��(l�k7�)9���,����6�/~A���� �r���S���J�[4==L�L��j�� l�2�F�w�"�M"�����:t�;�kM9MF�ZuȞju��rM�!��/��36E�z�Y�J򾩋�C���>�`�7����e�HO��������a������{̭�� ��zs�7��ۦ�iq���k)K;}���KM�w��{@�	��F�a'fy�)�	����0���P�J&��܂1��ڴ7b�w�����÷фL�.��]YJ"�O�:�e�">�&V6�9�x�M�������so���=����z޸?�[�rT���tWg�1��&H�T	�&[�A�u�oi�.ތ���A�Z���DؒM	q&#��`�j)���v�W�����at��eY�wm�T	<�\�L�ۏ$B��24�ψ��k����AQ���rY�1���Ƿ�߲�A6\��ִAD ��״�{��j�
�hUS��6I�c���+���k�4u#s?-A���-`���E'z�;�^G>����nϪ�bU�����N���ch�?�)�� C_��m�轠.Sk�r�L��fjޭx��e��V�>�E�>�N�O/s1���n���y�]�O�Y~	S����Ia�QZ�7�|�f}�z���g�O��1��+�A�UEʨ/r&E��)����^+(�B�\�`y�L��p��%�(M�/�U��e$�Q=��/���)��
w���z�Z��M�S:>�%��@��4�C����O�i�ᐴ��~�t��V�W�v�)#/�IM륹 �3-�Ș�tM�����'E���}����-�jA�"e�qyɗ�!2g�1�72�����Sç_�W��Y��+4�4�+0:�v~`'ML�\%��;ꋬn�)��#k��B���O�bq=�ȹ��󟚯<T��u���`̎���	���zp�ҲH�טVr�(��"t�ݔ�����vt�����+�����#X���g�n�4<<�7*d
�'`2f6�a�R�Q�x�vH�k�l���.�e� ����U����`����ٵ���Q�]�?"��K�����!����p,v�?ة�u�/#D"��8��*;��W��olH�����i����,bx�'Rv�X�,C�ϫE6E�KDO ~�;�w�}�+>���v��]de�&�B�l*�z���)�N&���:Ѱ�<D�$��:v�)�0��>vS������{e洝�懤i�e�j������ �@��DDB�"��L���2�tgَ]yzN�w���YR�&)��=�b�-a�A^-�Ç�:���/C�?�!�*KR��s�� p3p���8t /:� %>�T��4}����S�-:ȄH$bC�����AO�F�⛽m�=�a�^�H�_V��m�U���J{�͙�=�1�ݦ�juwu+�%nX�T��LE@�5�d���XφzY�&�J�o휈p�ޟX�]	�-s���"|��i�����?Q� ����-�WL��j�h��fǧ=��S���!�����uɋ8/����cS�O����U��昫���}}$���"6꿬�xy����t���BZ�v�r��Z���w%�`�#��������h�	$�\z��.��)%�
��O��b�Ykی��llZ#�ܗ��^�YY�
�Ki�N��,�1��u� �3�����0�>��A�N�􂭂�y���3؝��=��=���ĳ���e�w���3<�3t�骣͎?�-��y�U�7����Ky KY�������������[�4��6�	[pm�q����\���,�h߶���g�/�I�#U�!�)z�pE�Շ���s��ݧ�7��փ{q���\C�� �&r-I�;���kR�`��sN�d�֓f�$b�K5a^����_P�n�fW�1"V����#�ۆW OZ�u�Z*l�H0wҐb����K䍳�'������vL�-����N�ހ���_Q�n<���S:�W�<c]]ت��&"�\m�%���E�Y�����	�l���o�ʽ�Lw� B�'O\���4��h�	NL.
{�5��Z���f�y8�3։D�˾6��P�\�0Ϥs�T����C��ϭ�y8t�b�m/��<�8�H�_�~WF�i����-�ڼ4H�p-�}<�=m����.��d@���!����PD���v+�CL>��S���]:�?M��i�N؈�Æ��I>Q\�%a$�M��\Թb��r�pf촼.G���\$�ڹ��xv���H�tωٔf+W��H����f��-߭h/alԶT�1ÿ��m?ťХp�P��oe��N?� f$��P���>���TE��#Y�:yJ�k���1�I͙qT0��(疢NfI���)�y�Z)�C|��:�C|?�X}vJ
�������{q�Zړ�T�=IQ �)`��S���,֩�bדY�P�n�Er	�����#��h�4��+���sq�$C�2��1�B�C��R�
+�A��B�����&�w廓��(�-���D�GRH�fe��݄`\1�k�AGmC�������9�x9�5�*�z�#��ײV~:^�W���U��vd�?��&(��S[�ms���;�D�@�Ux�Z�Dh��;;Eڼ&�m��~��\iS�x�o~XH�?6H�þ����%����T�'�lk�a�j1�Q����hO��XϦ�}��o?�w6,��/I�$��]e4O$���B=��c���H�xAR?�S��[^��Y�<�~;��9�3�$	�Ҟ���:�0~���Ǻ�y�9�����^&��P�G�ښީ��ѯ$n������ٶ�zw��l�tp��L�E_jTp�� ���[��b� \�����W�_�p`�*��_q��B�Qy� 9zנ���
� ����>L��~�\��2h��?��U�����-��)!�*�Hw��1<�����θ��c��=���/�����7B�s$�~�8�:�����"x�������]�:�I��H)�����'䛢�繜����\&�L�ڃޏ��g��ȍ#�ӑ��.�L���*ՠ+�N��6MU���0�=(_���/Ƭ ��X��:*Ǭ�c��+���t��L&��^(g�U��I���pͿt����8�$P��^DwY$]2W��1�ح�G��=#�_��GZo}	�N��Z��X��,	e#|�V��fh�nF��ܭ{�����>+�����Tnp�|Nt�a��/eC�ŏ�:�������`(�؇�MǥY��3K�gٍGX��R�Q5�Q�(5��|c<v�}�0��DZ�����Β��{�X��Ȧb���K}�w���p��f�1(�'�NH����f�>���y�.�CK�}����*�0%"���q�%��z�>^9��4m6���n��Nsm�)*�!#��1�Q͓���ϩ���G���#���/������ 3�G��o�>X6\[��E�~������-�>T�{�<���X�~be�u�4>~��8$���3�xt�ڟ:K1�pz>���PP�`��ҔC���<��3Uj��S���)��"a�#���O�B�Q�qo��*i�5��҃��d�� �tr��K!�"j�ҭ��9�������7�����ce�Z��f�v����"�9/~�r{sJs.����H�Eū0�!&P��|��7�����R�����#���SO*)�r�V�8k��:\�Ǉ�� s�iD�wϱ����|Z���"=h�}�(�CэF���)�J��;��n��E�����������H��JJr��, �r�J�=�SC�"�i֜y��+qm�T4Ćn%�pEr���ח�-�V����K��E�ux�;u��9���� 7;ҥ�.A���-a��<���q��PC�	͞��N�[\e���өq=��)@p�=r�C��v��l�=��?˨	}_enA�����4�'�XJ��9g[�c�K�,���7qf�HDS��"���m�~ށȼ�J]Ҵ���(l4�Ō��6������;/w�=��KɮÒwQ��c+Wdy�86{��P�&�����w�`���AӃ��X͙r����청���P�csl�HM������MeH����D�8a9�pI�}��WEY�P��ze���������X��%���_\��7�ڔ�Q��u���]�~�%  L7�X�C�w;���� T�7�7U|�2���zE>؝�n���\[;I~p�Ø$E'Ɨ�f���hޏ�(j�0MCyV;�jzx�i�C�n���[{5TE�)\���f��������KE$��Ak�����n. ���z*A����WJ���$"�p�+QRYXl �k��٪���R�������Ǐ���F�;����JC�#�@��(�tz��i�dJ���y����s�:�;���$BM^����u�9ˢ��1-�P<o\�M��2T�s<�#��7�c� ڎ��M��1z�I��o`a�C����r�_���c�ܩ���W����TN��t.��

�9��J�/�D�����|��SgNz?U�&H�p� ֪k���q� ӛ��4=PiU��s�e�F*�:y�Qu*	�_���X2�����Wk)AJƭ�O�#�����ǩ�
cjVX:�.��y�jGCG�lz����l{7����5���3�x�*��/�H��">胠�H���W�NR-���1è���u�1�<�L���S��hu���t��=8�5��P�~y��P1�̪C1�h��t��ęN��?���O�E�B�H9��+³�ak�bX�]�U�N���q��O�Kz/5��N�S�g;�7K���e:���1LE��#/��@�n(����_hs�?'�	z=u$�r�"Xq�����R>U��)���W	�Z��'Yi"�:�O�ȃ{�*�H!�v���?8vB�aA�0��X����Ge���x70���c[�E������q!!w'�z����{��N�C8�S����c�gT��iQ`��a��bJ��N}nS�u��M��.=�e����-T�^Q�f�B�H4'�0b�	Hv��I_쀇Wݧ��r���Z��"�ob5i�s|@*P�oG|2��~C?���x�wļ�Z����(����D�.��֣�Sg��/��cz;Wj,n��YN�Ă����>Ҽ��G~n�{f[�����WI��$oQ�,�4ӽ3g�(
�eJ�$k=	����z�����}N�,"�50Yp���^�2�Gs̔��7ye����6��<������h~�_�2$me!�����>�D��&��I����%����N�	%��Z�V������~��x�d�ۑV׉�f_x�+ ���D��jL�^�7>��o�����2b���V���6���e0��ZѼ�\L�ԃ�&yp�⦪�L4o�N1T�qJ~=����ߣ/Kro�70N3�ڰ�O���G6�P��H*��`�C6|���s�DY������<5�X�J@�����6�Օ���7�{�O������ :gj�����%/,�N��IdM�bg��5��`?'ܠ�%�ـ���F��R}����)j5�t�6��� �ب��=����A��C�@q5b��5K�sW7�q<j��T{�80r��n?���y&}'�����e�w��6�x�/���_),P��01s��Qt��*��i�zQ��w���l&���^b<�D���t�1�ߺ�c6��!�O#���u���R+\�B�x�5cĕֽ�;��U|qK׮�f��F��?�ݯ�|��,�+�Oޮ��YH������tU��C��=]9�ƕP�Ɍq���"�����*i��NQ�^��	�N��+_'�=�7T����T���E�/%@)�/\Z[��AA8����&ͪ�G�k}�]�c��H�c�>�=���{�8�D�:*����N��;W�A��Q�fZ�a��#�b�4�9y�{�]�����󒍭��ĝ	`+��=z(�P�e�:Lഢ������@Xd8��k$�r�M(�Lk>}��%�����C�b��M���MA|���i?�CL΋T��ȓᕌ1�|�ap��)��6�K�0�M�Uł#\jKo�����`�]aE.�7"@����΅��+��c:k��lg�7b�>�S�uh	�B�GW���'L��C���`��_"��Ȃ�m�����ښ̽�Bdx�&L�Gv;�Iq��AwZ�5/���tX��T����	~��j�孡Y�1���o�~���y)G�×q�D{,o�9S"o%f�K��¶����gD��	�սB�(�i\�O�j�Z@r�׋��n�݃h�=;������nj�-j{L�O�	?�!�%�i��t�+�4�es1�c�$l�C��Xx̎��R�ڛ��c���*)��A�|gE����i�<M^���\��{ ��?U�1j�)D0^%��aH�D�q�J� ;�?�;���-A
���?��w����FY�XfT;�<�����5���" �h�=l���}������	 �1��SK���6�������#9��/(�Wty�VJr����9�F� U�}#�ĉoq�Uz(/{�PP l�A?�_-���zLKdco/��0$1����n{�n�?�w�[.�s��n�_��8�n�@G������Dch}�7+�o��%��t���B��h��L-R�'��K�Ĩ�*CcAZ�w���E��d�E0����Ww��^����Ձ��$��b�<�Ê@E����Q+���XT-��w�vӈX|ZgǤ�o_kfjF��K�!��׼6U��ڰ"6�Pt�d���*����1wF�Ur_P߈k��H�ˎ�&������͊b�@�u𥎀��g��/��ㅜ�������z������ۜ=�� �S__k�]�K�$G��z@%�*�x܅��L*�;�.8��p�cf�fq�C��x�l�{P6d��L���:�c�S�)��J`�J�fz]�{�n���Y��z*��y�d�O㻵?�c�:U��П����v�ȹZ�P�
��_6��71`����=�8�+����\DG�����D��7�u���9�Σ&'-y#���[�mۯ�x3�k���c=�3����K.H�v�M�{|L�Cr�:ߒ8Vv4�(mN�#�2�1o���
���~�a�b��"H�Vٗ��a���(k.N=�0+C����A&�gkN��!��&%@J~%�%&u�4'�"���r@l���"X)Lt�����{�HG��fT������c`�I�`pC��V��t͊6�L�d�Ab�#��@�1\��ڒoq�6��?Z�c��4���S�)�H����C��"��/�}@{	�tFNR"����?l���t��遵�(��nO��\�^��>�ϵ-������G�SU˙M������
�}�:7�� v�~�p	zm�ih��4�QM�����ʻ��q���뭘�bf��1�Hg����;�
m�Y�_�E��el"���ʧ0�
���1���Ce�׉l-�ETf��u9B�8K�>�G�+�H�,��b������co8���]���J�J��39b�;tƗ�LݵXBOl<N�p��yW�"+���3Ɉ�4���Z�_��*f��P�K�d����ˌ��_܅�|+�CB���X���ûc��hHͥ���!F���z�ɤh}!cl�4�ь@ِ*}����(�z�����"���'|��u�},~b�S#�Qu��v)7�r�䝜���Hn��O{�/�(��ߙ|5w~`��q&��2�L��I���w�Bq<Q��<�J�ep�2����Sp�ʟ��'�CXm�meH����TH����Ό?�l���\M����C�P
�q��dʜݒt*/K�%��C/I;E<�}z���ຣ1���v�s|J�
�{�(UcH�9��`�y�`�I�w�?�t!{�ʑ� �V�
>}Q��F4����y�0g#dA��`��2m)m�t��kDND��K,�e`G^�?���#�)�����T}��+N5���XJi���+K�]y3��̰҈Uͭ6�+%���� ��W>���d=z?Y��W9���*z�	��"$�ڼ�	z����U����Y�歧���c���ty��17�HWP��l����,����B��mew�1��t��z8�ɹ��<�)�q�:�s�]m����!*�����~��P�<�0J�	 ��c�uI�����ഈ)hZ�C������b����-e��ڍi�,)��~xK��'��9E�3�l���c��U�g���@s1��e�z�7�gO�G�ԓIDd���-XrbE��E T���}���@U �.��ٴf�#1�<3�gr�:��̛ �y�������=�~�a�|\IW�̈�N����7eA�"Ϊ�^Ц4"���Hŉ�Ҭ�-�� X)1|.�
6�0i6Q_c�#qܝ+{:��Z�»�Ӎ�7${m�Eǅ���ߍ� yt�n)c��.RrI^H�$���"�^�s2�@z�͜�uc��o�/�R�J�?�f�gMO͖D��#�᎝���]����D� (�tZ,��N�do�N�\ov��{s�x�\�:�~�D�·h>���S��c�$���Nb]�f�^�X��d�-mξ���S��t^����/;f@���XZp��Ւ�I6i�����1y�sBYPZ�����c�����'�l�[V؏]E8T>���[EA3�
4�-�M@It"i����es	{1dڟ������ud�JG"nhw(�q�[ǻ�K�;��'��a�I-��
M��I��j|��D�"�+#_��j�#����쀶d��E��;�"r��������̰�b͹,RF��X^=�f�(csW��k�Kzq�ߨ�r��;�K"�i�t���i6V�5/�d'�^"�E�{���!Ld��_��3vv�ɞ*���gۃ�9�P�} ��"F���a��.c�r�n%d���*���V�R��̵�#u�Z��^}�H~�?�Y=�qJ��6�]�X%|[ L�#�FaFfm���n)F9�>�ː��� PA�o�eտ8�+6����M��#\�ţ[84?7R#�!4�1�B���3`��{ܭs#��WW��a�"����~���h� ,gqr
ȠP�}�E�����8���e#nN��d@��;��[Ef{��.�0��j�>�!.w�/�[J���3&׊�#2�:lj�mh8����lr�ҳ�;W�Ʈ�����^MD̎4q��P	��>�f�H�'�	�?�A9�"�!�ҝ�B�5�wל�<�����-�\i�&�H/����k�L_v[�dK��TA���&���@ݽ�Dr���*˝G���(.��m��]z���v�B��R�D����:;�F<��R�	�A���4(X^�h�v]�I=N�ѰqF6��8Pݽ±d��MQy�O�<8V��J��< �LW^�<b8����������7�A�W��'�%��X 2^�;Jȡ�'*���h�:�\b"®�RDO����:����	5Iq�B?c\��w��N1Gtc&[`޷f� ���՛P�κ��͕����~Z���AZy��WX�9̓���?���'�K�ف����6녪_Y��Ż��#a�,!i�8�]�#=����ߖ�>�[ d�U{�L/�g=�-1�E�O��/���n�/��Q\*t�z���o��V���� �:�wML�sE���?�j�2ŏ�m����8�A�R�;{q#���l�n�a�Ν>�6�Vj�X����)1���]��,����
.xњ*#�9?Qj�Q*��]l:6lX�Ȣ%���g��X��MX1�'#
Bs��w߷��^�!���q�=���ӂ�ֈ�`XD�'������@�CI���⃃-6��>�� ��6sR���A��q�Ҕ�hs�"`�T������R��)�޵��y�x}�j�Z���O�+ĉ�&���B��u��YUV;Gv���\:V��ꀭ�yC>9}���r�;Av,���n)�����`�ь����>i��#[�ܨ:����zL��=��9�]Vu�"H]M�F�ɬ>�-Zq�A�-�6'X*6��:���B��� �E#�b�����O�EYo�}�'����` &�!g�i�I�*�G�Sk�A�rg*v��'O[�������JKcE�Մ�4 y�-o����zG���a����X<�ޚߧ�ۯhPV&s]d��s*oR<��8��c��`d�Nz7Q�b��>Fux@%�PL����e��v�m���KL��P�`w�Z�𠡟�"m�V�Y�%������E�7��Z�F\���ѩ-"�2�Q�Buh����W{Z-�K�����"RE�a�\��+[.S��e}��p��7p���h��F;���㫵u�rC����z�K��|�7�`3l�I�Bb[T���X2��p�(��\����F�c��@��~�Ѭ�@mz�NX;��.���9ՙ��r�d��-|�$���g�J=�Q'^�V�^@����u=��sa���iۙ�?z���̏PF�� ����6s/�G�;�L��2�xA�˵}P0���l��v�hI;�F�z�J�|t_�����$�\��p�T�z�_���p�A���8Ц��l�8�+��&�ee��Tj����!�ZQc��X�2G�
��Dɨ���y����1�V$��^�
��8/V�d��}R`T�G�.k��`x�y2l�pN����֫�z�z�;�Uc�GpP9n���6[u]�K�o�.��Y�{U�|�e|�vi��͚�<��^��M$>��B�Ԟ���=�1X4��F�PR�~�Ɣ�~�xdIˈ��~��}��Ư�1�wB���ޅ:�����4�ۺb����\���M��x
X�[�`=j_CN,-;�< S;��mH]^�G�J*"�"��.��J��3�Ϣ����|ݻ�'C�U�Y�μ���M���^"]p/vn9���Y:��h�;���GE�x7�neDB�u�&B��)��ॅ�0���*����)�J�b�WB��)t�˕S  ]T=6^��a�\����P�����F!/��۔���HX��"�rJ��B�7_����9Tx]}�s�y�t��A�qۥ�5�>a��3�B���\���!2c������g�˕��� �a��2qHH}R��q�g�՟�IGs����t9w��Z����9j^��ݽ�h���g��O�2����d���𡷤��
����̒�?|K�[��ő�(Z��D��<����63S"� O�\�i$x��ך�1�{21�͓:�r��@��WJ�-<�a2=[�O���m:���V�Q�i��S��Pu,	Q�<Q�ī�$�{J+v�a�+��悷%z�B �K��ʓhl�r����<hy������?�}�QǷ�����|_��ڿ��}ƗWf�QaXKںW��`��ax��:��:Ew>�G>���˓�ρY�2&�O�=��D��o*�bׁ����&�^�&|��#���J,�%0���/�l؅����'f������%��t_���UK��Z�|tV	4���hQ3Þ�d�4��W��0��A�����T�ĪK�X�%�M�(:Ø�h�<5'FQ끺�4���c���o���`�W��ܖ���nn��]�1���d�.+���X�E�D�LS7���76ϴ��#��`r���+р#��6���DZ؈L\\#�����b2�$��H+;�:g-&4��R�2	�D�x� y�rM��\�x�G���wQ��G;���w�\���?�8��K�YD��q�c�1�ˈ3g(@E�?�e{o�z�;4�Ӳ{}��X!TŜC@�rrD}�4��ʈf�@�z#�]�4�48����v��bW���j�������*2��ωA�:[�B|~ �Å@~&�h�H�	)A��������^u����)��O��Z$A9LD'�	m���e";s�N���7�~�I�X� !�T�Q��f��H�A��'5%l
�!�?Ȏ��ѣc��z��]�<����a��5P�X~q{�'�����_tz�1�w�m����Rp�s{��	��6��K��7�K;�D��Oᾆ6�%O��7�J2rJ��S��P/$�$[]-.� ��Σ�l�����zE��b ��6M�ޒI�BB?O��@J��韘igi�{VEu��m�0��!)A��P���I�Q�xc�D\:`Ȓ�Bkz�$Ӛ�Ml~A� ��>�"@�g�vŞ�'�����
M
a'(
��;$Y�^�d����]�1�b�)S��|���K����G�nD�)��~�ex�p�3Z!>_��פC^6DP�K41)S������j����۝ 'g�iտ;4f,�kt�U�T����9�K؟�Ե��S2���Y�If�9I��L.�E����3v�m$-��ko/�-3�C�ZL�w�RrX�	��z��AC|��#�U߰�"�RD� �{p�Hؖ
u&��A��.�d���&sC�"�=��M��6.��?��m�X| ���j����&�Ί18t�T-sK^�P�.�(��q���Ȓ/����P`�FtJ$1A_��םCI�E�����'��È��ǋ�f���$OU�0gU���>�K��=X��ֿ��Z�K���<��}Hv)|E���
ؘE ����Q���FT�0a)6Қ�������u��r�������ݻ��d����>y�k0�/&;���J<ğ�Lji!��~Oۮ��$~3�
���: ᦉ� �4w��{4a��j��
�+����]�+_��@��P���ˌIH�'�2�/pl�n8���0�k��!��[�SaV����U0����QC�)�����c_�Ɛ��Q�,�7/�v����ѳ�����}�o�a�m�5�h~)�:��7U~�Tt��.|� ��Rp��ض���s�� �S�9_��]o#yj6���	L;íI����$XlCx���nT�tOa�A<�:h��j��T�[�bP`���Mp��خ;�atM�z�):�w�4���������@���H<�A�Sw�A��R-��| ᖡo�T�A��N+K0�u� ����`妧)�n||R�^/�!v��^-�;��0�s0�Zϫ]�����^�h*;��x0�z�$�E�z�K�C����� ��hSs�^6�O��뎬�\~7A�,Es_% @��}ڽ����+Ğ[�:���k�*�H ?>Q[2��NUQ��M���f�K����WZ�jX�dD�P^l��;YO!j�5�C(�\\�&���o��(Ă,Ǽ�ԁ
�g���Y�~��/T�Qϟw�*A�>�'&�#�kfB/h������~�V����l�t��b"3�S	�
���UHs��	n������(��4�	���"I�������[~bll�9l��^B��h�d1yj�:�K6*�(�P�NJ��Q.�k>S�o�\�*=U�,I�k�ɵ��A��N��/�����U����4f�H(��q��ߍ�ĕE}.�^�����1��~��:͕��0Y�֤Cl���l5	�p�Q�6�5���r�9!��I�Z�\�b8�#ָ����ټ�k?�S?���UN��?�U15ZI6�(�Q�0Ĺ�[�ܙ:�"�ˠ=��#t{�Bٲ�؊l�m9�
�ԯߌ���Ϳ��6���"^Qdl��0;�P�Z)6�:��e��J�~��u7�T�+X\�c�KZ6g,Z�Oy����;t�݆�%��ϋ���gq4�:rc�����ů(c�aw�yEEit��x2HE+��Z�Qd�S�(���Vf��M �lCq�A>l�JW����ao�uO���נ��f�-~r}�)`.]z)��g��6<r��R��%$�a7TpXl��>�I������ġJ7p�j��t��/�t�7�>���pq��J����,%��l�Ѿ�Z�f�'�Ŀx�ٙ�M��<�Bq��p2�ظ�#�K��صb�޵�����D[�ʚz��l�rW)���q�(5h^tEU%VG���!�,x�n���"H����e]	�A=<�K��=�4P��@�A��,�۷�i�o�ʳ3((}�\�'K�ˬ�H,��W<��;�۷�:ټK�+�T�M�6��[
e��/��% �?'l�3�������j����w�O�ײq	���ܣ��~d�뾭��י�D����L��?5΃2 MU|�Y�a&X�����g�A�2�Û��զM �&�7�����k�����tNuϭ|i��S�L;9��J��i
���1܇�3���p��ijK��CuS{L_][��}W� ��#[J�� �hay���le (�H^��޻�0�g�����M����,�şH77�crr8�
ةR�����f/���7��ޢ���d�A��BƷ�_(>��>�d:���� V���
:����*&|�������������,��w6�o��{ �i=�?ˠ�ƪ�������GW½��)�6�H���,�lJ҄D��O���!�;��"P��pX׭#��W�f����X9%����ǳ��Y�X;��K�0~V���MTA�:��9�SF����ksdN7OZ��ې��t�A��
�;(����ݼ���2īh	�?�H%�&�
UY#�`:�����y��h�K�r�=\x���~��>^��GX#$�2}E��_&0��������Q�e��=?��/ѫ�<�ؖ�Y�~��&ٸ
G�tu�}�+t�ʽI�F�3�a`�(1��46�� #��� 4�m�P�J*�� ��V�����8������IF[9G����Q�>U,۬%w���Ȃ����^�Z�10L�Gc���6x'ֻiC���ڪD��[&~P/�u-a�D2?z}iF�F�-�q�e��˒܀[!^��%D���w)8���لuV �k�I��3��UaXIn���1߭s�}L�5*�h�zX3X썿/���|eMPf��N���8�3]�Ċa�s�+�.� �)Y$�j����6�:@˼�yWk,�����rL5��"g�:��N9�l��B�3̡_�$z��� o�GOu����(�h��z�]�3-v�GcȪ�} �Sc���`n�l�Ě�Ȱq��5���Ad�Cs�6Ƞ5��x��; 0���[˸�	���X^}�+v���p�*��}��%�MQ����*Hy�T��҇ܶ0;�*����wP֮ptp�^*;s{�ui"o<D�g�O��q��!�>�]K�D���	v2�	��X�hѐS�٭��Q?]bS���!���b]w��"�ï��H
�
�;N]11F�F�j�&�e}�8<d����(��8N�N��V���p7��|?�*:�8^Ԑ��.���3��1�v<��O�ך4�Ɵ�U؂>9!t7�
��W^[b޵\�������wm#�[�V��[��ӏb���L,`=CR�C����KobT2���4���hONe?�hdP]��K�o 4u�g�s���@	 �f̺�
h�mu��X��6O����KΎi1�?�i��ؼy�kXz\�1	D���D�l`sT5��N����߁�'QA�,?�.`78#��?�)�e�bO~��JY!��\��S��[]1�P���ǡ�(ι��'F�Bt"��k��츶�x }Tƞ{˔Q�v)���Ǧ��%�]����W�g��uwm���	hU\�h���S���s{ߨO������طM_8=��8�����^�_��ݦ��tµb��JN\�D��R �|�"��?���v��9��-��K~����Vwq�\��`�z2z��NL�f�� ��P��E�N���ۊ)
9万Q1&����xg�@��*�=�Sd��yu�@B7	��J�`�2/g�daW^��f�eY�O�[9��4���pbi��gn R�Zhب��ǃ��2Q\f��m_hg�N���4�5�˺�l�kz����(]'��fTހ$��.<2-��_]~�`x�.�����)���F4��ŔpW�P��_�_l�;�^Sm�:��&Iۿ���Z��R{�����x,l��}&̡�&e�tn�³i�_"e��T@_���&7v�UYwP�ț+��Օ�o�%����q;6Ou�������Pd����qveW	woI�:�Ѧ��L;q�}�[���fyi�󁌤��N��)Z���b�4�3�ӡ�6�b{��7W>��CD�{ IR�����r� ���
"S�e	�>�f���Ӳ��k���J~��u�i	���ua1|�;�i��m�(g����>v��$�C(�������o���38�&�@�j1�&^�`$���$�d�ƌDx�8�}�՚i��X�p�8ՠ�CH�/T4��R!`S�Ug�U���'+M�x�f�M�fw��uݬ`��#4L�p��ڃo�֧$���]>�(
����-땃�зn�+� K�qUM�ۀ�q+������*Ex�cY�"k�����P��k�	��7צ�zV�9��Y>4n��Dv'l�%7b�3�����ɀ�GM�Cy쾗1�:�}��֝>��4�3}gΘp�GA�[�7
��j�G*� 9ȫ���	؋$���\]qhX:y��WDe+��	-�Tv��ݱ�~�	�	���yz�����H� ��ȶ�\&TĆ]���A��;��q�+��3��&;g���b%�a�}�0M��ܭ>p���HK�M��D��� q�������A�L�iq�O�=��Nܴ0�)�}&'
�c֦U�!��Ӱ��?�l��H�s*vSPΏl�۠_/ϲ)������9��gu�p�2�X�-ǰ=��m�8!z*y���&S�M��	R�����#o����Cd�0��,����(�8/����s���d~E���y�&&a�f���Jz���eK�;�Q�w\OU�3�%#�4��sDZ���Y�u��'<햇��e	J6�YZ\�7N^���?��M�Ȱ�qg1��28}mK�m\U��IM0ƅ�7�K(��Q�ʯ��:P\�W�ቕ�RlnW"x1�������)ϻm�n�Tuzn�31������ 4��
�Ƹ�h+�P�+�������iyd����۳iI���G鉈ꃿ�5���,E-�(GJ6pP��Y; ��4�h$���Y�~@��l���jBop`������ ��SD(	�9����R��r��c�:vx%�+&��y5��h�ʙ��*vFE�:1�'�x�����B���&7�)�@܄#�d�<���dH�.`f�ǁe�'��)&�⁫���8����?*�˰��%�g���j���c��mc�B�࿻������D6X7�-��7?���?@�����+��d-�ZX|���-i���j�捓�F�g�<�,�%-,�q�\7�4F�9�Ӄ�b�������9������~UƉ�����\�3^3�;�,)X#4p�/~�Xʧo��OޱĬ��Pt���4���K\)�~^�lX�.4��f��1\bY�\sPl_�hM�>�oE���e�G�cn���d�/-��������˫U���J	]��s:��T�hHu�]��u�v�{m�8Ȁ��&T�;�U� �P�`T\f��rG��U���	bg�N ��c�b/���S�sѽ��:��{����k��E{B)�;���k}:#�D�K3Kʉ���Z.:g�%;��f�6�� ��.��dB�q8-����?G<�1��r>��1O�/�<F:��~�1Ly��/�N�f��Ge}�2�X�N ��o�N������(k����T#�@��$�ݓ���9���h�E6rG��hA0��qg	u���:x�#��*�uYhGLO��&�^q�[H�4�\Y3�NWIC�W�y(�&ϴ$���[��j���xX؎!��@I\��_L��z�~�I�sd�)�Y�^��>J��Ol��ڈٽn��D���"~�Ӣ	<>3y!����`y�W [��ѽ��m��3�j�ەQDG������g�����������~t�\���f5������U��B��v��C,8
�?�A�a��d��ݒw��ev!� �����J[FN��3؛���N�z�S�,�s����^"��|9ޚ~�P;�|=�P�|���=�$SXj-5��O�;#>0��l�t^'v��:~4�~"�vP�����&3!U�e=��G8�H��P���U�-�}�b��K�;i��sIJ�x[0���jd4W��>���S�Bn���;N5q�S���Wʉ`�I�ab�����ts�h�?d���0�/��7��q�СJ�o?Ѷ2KS+���*6��F�ƦtQ�	�6��k�.� �&����߇)����0��ւ�ش�fD��Qt?���{���S��?���Ο�m@�)$H�b��j���D�Ъ�h�G��X��^�	n�&��3�Q�b�ZVBGVA�C���Q��)ah�}�nŶĽ�F3S�,(h�핚����S��t�>�H �P�K~��J�ۏ(.ŵ����{���1?�T�-)JhHq?�:���h��!��έ7\���7D<�����<��f�>!Β�Y.��.�PN��1k�5�!5괓{����.MoO�]^ɗ���T��[J�Z�;��<��������od��Bժ$�f���4Mۥ� (�-m;���n
気1�W񟮂n3��B#��Iu�V�$i.
������Cg�)�Yl2f���=�F;R4��D�2[�i�_\`�Uj��*v�2��k*�����#�3Wj��i3�|Z��=���m6�^
���L6��x(�{PvQKu��K��8;x�5��D���;��l�^G9����hs��׵�+4b� =@c>ɌX62_K\�4Й#�Xl�k�������Ǌ�:&]��Ѝ܋kD5�\8+�F8�d�0���=����;����nf*7+`�H�o|_�O��Ӟ>��dwI��*�Z!�%��QO�h�BD�&p3�-��&����Q�?�f-)���/ë+��y��q��)�e��r^T �kH�u��V����1�%c�u���C6�Qȭa�~Ӟ[�Ĳ{���X��@Y,�Ġ��e��շ�lW>��LoO�X�\������sPz�	3�UTаZH��O�Y�jo�Y1MK����6����}��pk�`L|�eǆb���8T�=A��%E72�8�iF#����^9�4	HM�$���s=���y���,g�gq��>�s��Jɖ�5x7#��Ycy��[[�l�@���9�O 	#pQ�;;�a׌��Iۇ�ǔ������j��>�Y��mφ���������lC�7Ɇ��&@�,n.b�[>kS"ֆV��xL$66$����?�71s�g�g���D/R�Y�)��x�(���b����H�xJ��ձ$����FbX�r�������t�B�1��+J���gu�Bj�;띪8����ݟ��B��u#5�ȣL�]t�FEr`�q��O0z���5
~��Uu���G���xNzR� ���0��ǩ��,��җ��>Ğ+9��L��eH���HW���G}"�/Y��FL� �Hi��$���M����D	��V�b�&K��UC���
�)���E��*�d�MZDk�ԅ�*�n'�y���q����1_S�RO�}��?�C��iހNU��BY2���L*V�Y?����xǔ�ǃ�u������������ck��mh�Y�\����u\��{y�j�W©%�U���N�H�Ē�A�X����j�m��w>���@2w��]΃WPc�li*2���钡��UG���9�*Ѷ���3�G��h��{	��F����	W���
G�9�.-f7jޖ_��~AEV���3���y�N�)���'�\*�E�OӲ����b<�aȄ��h���Ҽ�k�����ӄ}Nfoq&�s?�l��另k;r����}���R����QTn��y� z���
��N����JH��<�>�]�wUL��m��Q�Η�J�l;��f�J0x˴��������p#��Y��E�va#ga^��A�B�`�-���z�1�����$<���ȋXZ9�E�#�Y����_�b���5�8�7noE��Ly�bc����������
�O��Avy����\��1��?�n�&F3�z4r�C�@w1���$OEs��k$�c�&�g��l�;o�C
�^�iɟ��CGe�4^͜�W��/,3t�q�<�����^3ٛ����R��BM&-��l�b�f�a�&�VY�M��-�Nh���/���?�����!�����cI �ZNcAz�.�oʂ�ձ�f�#؅���R����L�з�
?m��Р��(X1�˛@v�}p"SeWt¹j�k�H�3�N>�e��	�~?"�ַ�TY�m��'�f7���n�#d%����<t%Z�U������/0���8��}g�Ϙ]�20��`�f�IS��U��Ko�=�bM�}���Xy��,{��0�������
��Ĵ��P�� c��:#ϓ�X1tW��K��W�1 (���L\�m��'�uVy�g���T?ἇ?��	�-�t�K�c��P*��Ո����J�9j�w��KI�S|!0��o=IwM{h��فM� �ܪ�|���g�嵺�JX�xrt4H�sn��{���tY���#n{�`�3�ʍ��AM�ՒG.�%�9��ٵ!��$�����Y�A�Z���t	�����*N޷�/�.�C'���-C�z���ئ����C������ČJ�(���u�V�
�i�0����#�3O�|�(;g ���AaJK������؄K2@��0=mT^B��^�ĳ��,�W�iF�|��6g���m?��������>����G�����4?TƁY�IJ���V����m]p�À��q��<�sY
wW�HG�1�&c��\Yt�r�rƩ�#Q����n�7ӿ�!���>���!�y>�Z>���f��!/�lc[OJ�<�쟵�'V<o@��{9�R��PR���l1Vl�y*ف+���&�����`��F����3 &�H�V
���D�%�G �1�;�:����֐䬰g+���g��<�쓦?<�� * 6�*���>$����8z��!'1��S�e|���}�la���Ⱥ��V�x5Ρ6��`X����>��U�'x+Y�g�tù׏�s�R����sjr�Ąe��2�t^��e�P���7�X�oK7�����My;S�t���,n�Ι�k-C�_�1�#��������~X����c�B����t��G/YWwIc����w�n*!�c�~M�&X�=*���rF��3N7,�G�i+c\���a]E2�:k�T�P��~�0�-�N���ጩ `L�d�a�K��.��Dh}i��DL���V�G@�H"9�U��u���h�a����^�)�IwǨqJ` @��wl��(ˠ`M�_�:چR + ���.�(~e����7�?s�'/��>� 깦F���ث]pq,��ϊ�f�@�4��������6��?���;b@ Ԫm�y��{���x$��T�H�� ���5���V\�Nvkz~������
�w�P貘dT��$5�w��|;M��s�=����[j����B[71�dO|��~��)�����暹�+�!��LU�0}�_�	�2=��~���j�/3+dFF,3�dmT�E�	|:�L��(+y"�_�`8��vU�iG���t�<�U��&s�D���o�1��~��=������������v|�hT���_�؟����*È^�F^�?k?���aɶ�;+`��g$l��yv��&S�[AX�s���O#�r9�Q(��X9����0�<;B��n�h$h��ky~��Ӳ������r��ĩk��U����a6���5 l ��[��^p̾�=@����RG�u)�zl��8�v��tap6]�;Q��Q$�+zp�V@���������[v�'�"� 	y�9���h�_`!h���� ���Y�3�����=s�*�P�B�7�qvKdK#"[�QUOvgsY��������@�P\��Yލ0�}	���a��l�'�� �6.b%�<����%pq>Q_���{��hƬ�gRx��<��53��b�F���f^�db�hQC:��O1�'�p�� �|`]�?�y�:�P�f����
��ٞhjo�e@�\���P{Ŏ�m۩*�L7N����O���VP,$��~��]�s̗�#Q��08p*#�656�jl�)�,��OT���J�v����@)II��u��߾��,o�<}�@��6ܫWg�|�hv�+��dm���!/�߀����;��GU�d������f��b����ߋ���+/����۟Ƨo�!��]YG�?l�wk�yƬ2�����0"]����M�*Y��L�Zf�~�Hw}Q r0���R`��!Y@�4�0�7]"~�-`6[>�cT���7��H��t�Ӊ�!RB7=�g`o�S��È@
������O������|�C�[��Au}��07����[J�2�?��t$⌥��j�A�Z�����8 ��SM;��zLo�p�=�->��I�p�o�z�|Uȉۓ�rD���'i�Hx�fT�]�cl�y�����ɸ5H�"6)r� 0������4��Y/�
���kG'A-SIP.���jGT��3�x^�{D�P\��X�u�N�lr/}�г���[
]M؁���0��`���a��k�Ǌ�����@<�;�u�y4B^t�8c(w9�^���K!�^K��R�K���&E*�^D~4kE��UG�o�"�=C2Hm��bl�֕��ד<������4�u������[�y�wκl�)�,/Y���b��=���;��i��sR�Q/d�/�k����'Х,o>)�e� ��Mx$#QD�҂*%�;,N<��$����.o8%��0o�UxD�M�aԾ�4�(���-
p$z_^��ږ��;^Xw`=V�L��5gl�lR�Ph����d��cSk���Vh8��^d��2>6�H��^��R.�~w .R�ӗ���?��+7����Ql3��t\�S��n^��,I��Y�ߑ��NFGQ"�|�5�L�%�1T�3�ַ���>�<��1m��C��Ҵ�3��Ut�]u����X�A�W�r�c�U<�ўr���rl���2�Ӛ��?:� / ��Pz���dW4,��6�^Isk����jʔ�ؚ��l�;Z�?c7�f�-�W®\���,�<�yH�Ƞ��-��Vx�q>�v�SJ`"�貫���}F�8�o�(jN��V���]�~����ߖ;��� &�tb��m��N_�a%�2�����[ĥ��}�%�f�?�,�6��)�<*<�����e�6wi)���K�r�������nO���l�69������^�X�q~L�����r4b���d��O�so~�A]G�Nu�����e,���Ľ)�3�+�fd��Ikk6���K�V?�����[�q��2'���L�*���O����4]n��Z����v�%��"x̂l��6��9���?��q� �s�پ����F~�����3{�YrH��D�Y���2�T�^[3���Cu��k�1CF�s���aniߋ� #��hI:�
����!]�0J��a���@�I,&D"����c�~����4�|�j97�`�WhE�z�y9���	f�M��?a�6?����Z��ne�Z��n������+�9�
X$	��ՙ2�ޤ[���|W.�A=�y�^%��Z3�h��ނ�pe�`G��iw�Z�.0Yh�$3�P������.�Q�ƃnЇ�!<�����Q��wGt_�ZW|���Xl�1o $�~�;̡P|3��s��qh�>.(�D��~0	G�]�N�Or��Gv��B��j�g�.�C�NO!:6t�u~�b��JM����c�q��F��nK+���-�� �����Ѵ>L���W�nZ�'�L���ş[k!ũ�'%��</��.��St�K>��%)U�K.�.�%��>^e�V"�u��7��!(�Z������'nyM���/���z�/G�uδ��ѯx,&�$�d��Uo�@Ž����#���_~%`�?�L�8<��GW���Gm	_����\��"���[L{������0�|����$R��!����uɗ+�%�׸Da��q����f|����hF��Ж@�raS�ؼt���<��T��cvI�4d�7�vl
o���B~_�h1ԛ����a��.���6䁂hv�L녾W�~�c$?@f�݉�J�x�Sl��*U � ѳ�:e\P��
7h%�a�V"_�7z����`a�tИ�)�Τ��54�.0?n�@X�?Z���c����T�c�8�2�~�.�̓_��# ��Ϙn'�����q��H�TM,���B����&��P�;�3�D�U�P�s/sI��l|p4	5� Sk�e��_�~�)[�y?`��c�8X=U0�~����[��H���ǈu��шtּ�� Z��`�wSl$]j���>��S-}v�F@��|��y<��*��Xߧ<d��檷!��W�?��p�/x'���V1S�,�!5ߧZ�M��&�G�c���V�3�H�_�(~_3G'��I:�h�n�E�h�r�0JN�E&�ĵuw2C��LW�	1t�ܚ+tG��o����@�PB��O�g�^��ARN.Fs�!g����b���D�q<��ٰ�ki\������:(-����8�&�n���+!�8d2N�O�c��/-�hb"�a%-�܉����9�O��JP^ث�g+�9��0�g�2�ד��,���X6���b�s�Va��x���+�i�L��"���,��_�#c�RћP��	|,�L���?d�-�W��M0�H52�h�4�����k�N����B$t���y��N�@h��8�4t�$IG� ��hs��=B���&��p�"q�1Q�d����z�eGZ)��5����!����j��w'��P=Ӈ�=�thR��Yr�hS��M�|�Ɍ�<t�6�gw����\�Yp��.��V��ų�M��=G�k}X�b�'��^#�Y	�j@ă��T��RUf��@���}*���m���ɐ��^� '��o��	2ew����3.�j.{F���*���d&_W�,�hRnD��_v��4p�iG���n �l�/���z�%��4�����q���5�:h�pwU^�E��ǯ��[�"�>8G��v^C%r���9�&�B�%������Gv��E�:��������<�p��� ��(I*7�Ő��٩�)�&&��J��0�f%�r?� Sh7�W��;Fj:0��+,MͬaK?�w)aE����O��곓�f�\�gu��C��.;(#��$wBKm�i�#�b���u�^��Vb��x�������t!�1��X���V�T�[[;��ED3v�es�����.g��!��g~��[�ЀAG�/���؂D�)���Eu����(r���}�h��R�#��kZ��>���nr�[1S��$�9
1Y>�?7�^m�����S��1'A�|�1 q��������m�	ں)t�.���[$�7�sf��:>KW�mQ�E8 �;�^Bq&�z�а�h � դ��sHj�����o�HF�g2��いoCN���>���N���y���-�ȥ���$H��*�sKF`�����5�����l�Ѷ��!|@x��]qOz����.������
�&���Ʉ8���>��D0��O�NkW��PT��><`��l�+�\�kn�_�f�}���I�9�},z*	4X@�~*��2 4Z0�d���О�o����lY�m����c�a��X����9?;�zH_��x3�����c��޺�����^)K��N��]Bğ�:��R���tv�=�R2F�ʵlXr��1\?��ME�� �1���@)����e�����?�W��[/���^v_ˀX��/��G��.�)Ұ� �����f{�};8]��kJ��1lž�D��7��;��pͼ3$P�h[��J텚�W��H��vF�s�uu��1��n�?�) �5B�PA=V�b��9�(G�v��TLHKc૔����S�
T�l���U�������zx'cI�J�v�H����#nwDb����o
��e����5�CgA�1CEnا�[�M���<)iWt.����60�^t2uM��e#�>230\�( �絠��?2Q�/ޕ��'�v�8毼��`gE��y����$%��v��Z��p0��;�E��ز�?e���@�Y0P�ဣ�T��v�`Y�� )�qBQ_�ls{�6�N(�Q�� :�-I�U�FH� ��D+Aw ,������HH��2&�$��iF��6�S��w��\#h��(f+e_�-��̲���\��L�x]����Ճ�O3��\���,��n��9��_��HVݼ��0��	���Y�xɐ��m\�5\�޳�D+c`m���"����X>�Ϝ4}��������Kr9�i+5���OU[ņ�]:s���J>A��
�L�2P7�@bΎ��A�F����3�"�22bBlT6�U�P0���o�p����s(��u��N�f�.5>0.8�y����Ϧ�;���|Ѳp%�#j6�������c�O��ñֽT���� ��`��d��O��"�䵵J�<
g�fk�k�`����x	M�f�k*�j�'9 #�Pv��3�-+��e�M����Q�o�q��
Zʹ\�^�a!��R�`�3ΰe�{*[��Y����Ͱ2mzK㱣 ,1kl�R�s�=�6�	(՞��-D�)���ŲC�|wE�RRmK�=\�����K6�x�e��"��T�����r�`���-���89�MzG��s7�)�@��px����U`U6j
��\���˜��Üs�*]W�Pk�?� ��9��8�N�R�2�n��vs��16`.�6I{	-�;~�ڇH�M�/�	p�M�zxfM��o����;�*[|�X� �I�T���@����]��#��n�[,�j1�/������������o����C$
ƛ�zs��v�d�{�DشH7s�3Y�X�m�a���~�!�=�\Ī�gn�^?�����:��ktYt`t�u�e�md�az�����T�-Z�Չ���]S�Mղ��,���l��5�����~[�N;`-`�N ��a�\��ښ��� .r��N-���*�vg��W�A"�u�T̒M��*.��[��x�p�Ί��]�eu����ە�2P�������L�D�n%�cI�����	:̆x���u͘�@ ?&��5A]Ƀ�F�G%���������ŏ�����O��.�.�����ϒ}����
f������+ɻ�&`�AzY3����n<��'hF�6q�F��Q�%�HBS�gu�`��}c���I�ǖݣ�tYۺ&���gm���:M�놥�<E����"�+�+� e<��]dgQ%��j��z�r�~���E��8�~b��ujHuP&F�����t��gT�'�+��5�Ӭ��鷲W�)j��f�e��[șB��L���R�Z����2�*1����DQ��h�b�N�����/JV��Xy�1!�o�uw�
\��F�c}�L���uᢂ>�8�,��Kbr����u�h˶��<��m�A��钠�|�0�Q�#�Y]E[�y{��(�*�3��g1O��_����r���W^
E��q#�sp��&K\�O{��D�/Z�5�	����&jp�PƳ��T���ũ�t�z^ύ�j��n�zQG�ФZ��ô�T��� �B�
 Y���*EMe��-�0�.�Uh�����\K.��zۜ,���T�C�K$����HD];�٩H7�ëD�O��k+	myK��ٵЫ�g��Q�K���
p����c�MnJ�rÂ�S��z��z_?�4ݩ%�Ǆ�W6g��X�Rw��8J|�c�+vd+L'
�xІ�O�խ���
�\�:�<)i�uɈS�O)0~m
0�<�'���l!^���D��z�҉v�X��"��
)�*CHP�+��U��;�"�h�u�E���fzY����0��'߭��1�}Q����K�{X�;P��B��r�o��A8~3�x?�%��f.�����n�%�$����K>(��t<]B�gт��L�;R�2;%�?K.0�GBV�m���v��ks�\-���O�Yy�A��M�J��K!�U��ӭ�/�)�8��>S�M���O�m�� l"yz��
�S�r�h����_��$���
9@5D�\>>5�
��P�s����:�:?jB涠��������iTx-aK�Uʿja�� h�]��k4����am-D��R$����E��L. �Fqګ�Шk��I9�֥�ǹ�tJ�[�I�b��W�x7��Y�ї�==�p�P߹?���զ ��it�ȳ�ŝ�E �Z��r�i�P�Dx���w��˪����%D��}}£��ӻ�ʹ��s]��)�-�F߀qrf�#N��sŵ��4��=M�O���]��l�>B��,q���@L����-t���Ri reb�t���