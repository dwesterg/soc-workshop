��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�BdMjÍ���di�#�rT��Hn��k��gw9�~\�U��b��� �M�( �c��C1,�YY���5�`��&HA�W����/�Ԅ���u;�s�u_�{�G��%��^޲|^ew��0�:�u�;�ŽU��_�9I\��sYA0~����{����7_���}}o�܊�ǜ�L/�D�NK2<��FQ�3$�؀ᤡHٗ]�pn�MC�yT�]�R����@�D��rI68��X�x�����1������� )S++g4�+���p�-���S%2�1��L�b�{/����x�\��L��j����P�x����\K!��?1*�m�"�	��NfC!0`���M1��'����A|�]�2�U�q��YnhP�xN���r<*x��upt���W6]2�6�0	?T,���qX������[3�i�1	yY��2��k��� �8� �T�5���ݸw�:�Yc'�NIb�����d��U�;O�y%��e2�$jjS��/\O��w���#�@��}�E�z�q�hܥdu��T@�>4s��Y��A}3���H�����޴�c"V��X�g`R����>�?�
)��q�O�}�Rv>��3����U��i= O��Y�U5.֛��a��}8^��ܜM40䭆��}U�P*�1$S���aB;��ߩ<�j�E�S���a���^bVų��[͗%>*5���f�=�n 4{�~ D�/�ɛ�O ���%lJT���X��x�V��?�T�������;����3��p���.XL���X�,&)^��;�D�{N�j�@}�a�	�T�w~]��b*=ɨ��9���6�pr>���\�b�e����:j?������K���ܧ��o�d��%�X�|m���wECH��t����a���Z�^_v�g�����ukO��/:��V�F�4S��`���u23NL��sPS������x�n�]cX���]k����O�*�ؗ�;���t���{ϳH��G�$2K7ӛ���U�똻_B3
�*q�-���_'�؟D�[9�x��f��B�3&{��dk�۬R�gx�� P޵"z�����N�6f�����hQ{����x�A��E�[�ys����./�;��u��I���Y]�Όb�tP��I	���� CZ�z�f�Q�_
.W��U��+�Svf�Dϑ�q��y{>7F ��N�Wb��\�U �����$�S-�^#���xRJM���g��m�_�/����١Ă\Kw_�ٕ,�LU�Hs�Ѡ�c��Oy�1m��P{&>ڔ��A�#<JV�ځ9����QC������U2z5�_��}�'V���yv��PY���#	�n�TM�>���Y��|SU{-�ޓ�`4+|}q�]��\�HS�KMu/����և��aö15n곒�����t�����m�a��Rǡk�����7C�dmu��T/<�N���kB����L��pXwX	= 2�).KA�4D��)�����f�W^�|�NM׿Z��2z�5�v(�(6,tN�ݑ%V��3e���;�@�'�̛�vJ�ՙ/�>��.�2��9ǃi֑����Q��$"��|:���CB��X{��u�"QFG��W}��/�צU�_b�W��v�	��Au9TB�������z&	3x�V���!�u����X��/�8^k܅*LÉ�j�7R·!�/�KM8��.{��"! ��OTu(���<y)F��w{����W�avYV��Q�� k$�\�U��y�LZ���i���N�	��x���Q����U����'�l>��7���Jx�
Z�������U�G�4`���n!*H��2	��	J��s�QjW�:B���������x=�H�k˾��/9w&ɤ/�A�P��6���ps6��0�����B�T���Ïcņ�fb|�/�L�قjT���	�Jn�cv}Q
��<+i:����.�%J$��&G���Ù�)�U�N{�"�PFT4ra�����>[�?B��eD���nZT���T��|{t��k y�8��Kf���{������27gfP$T	���7�:9j,�ۃ$6K. �5T���\�T�5��B���E� �1��='�Ye��w��_F%hYZ�֪�+��������	���F���#��Omm����砽lw�R'ۊ����*�I>�m5�S��79	��p�dO}\c=3����H� �L��3%�3
d��c���.�#C�F���Ѻ.|�A{~���c]��[M0�vh�|�=M"Z��*��()��]��ɜ��f|r��J,�S9��'��$�ѹA�~m>Ș��k�b^�ڽ0����I����4�;u"����O<����{ۚi������J�݊ ��;`�x7�~����-ͥ[;<��?��C�(g! :�	���zE]�F1�����Q�?�𩱝�V�T���L��Z�w�zB��I�v�|��O��"i��}�_�������39��_z�R��ut�dKi)e��;m�ww;LkY��`��0Sj��)p�}
��> �~wS��DqR�T+��0�r{SɊ<��vGL |� ���#�/��J��p���)��>I:������،C�p��Ve�:��e�.j-Lb)����/3mi[S8�"iy�&^�Etv�I1��n��2U�h���>d�����5xh��be�j�ژ�X�d�����C��|����so0��8J'��ї��Ə�YS�"�ʺ�c/z��Uφϑ�GQdH��2��ĥ��z�������1D1	Q���_��\���t-�P\e7�Z)�m��S,�0�H�?|�y6���]8Jar)�<�_}0�x8w<L
��C�
��|;�y�G!JX�Y���1b�ۂ=��	�ç���J�ɕd ifA�c���1���9��"֚%R1���~~r	c`���㞃��D�|��E��񪶴*s�H�@3�a�����H��1:�Bf���!N�ҏA�I�A0ȫk���{�<�Tw� �6���E���Y3�Z�%ݾ�v�A��2�T��jL]��{`��ؖ��Of�Ÿw{��c�*��m^�X�1�Y�G:�e��KǷ�?ͫ��*t�C�%$�� ��M�c}G���3��+�<��	Zt��x�'�2j�6�p�k0H���-��q�%��+��_�V���-���bQG<��@��8��k@�*�]�Q��h/lA�',I�}��m#F�j&dޕ=�"&� @�̂o,��l��b+��~ut5�����;�m�0C#��	.����R]��=��Ϋ�!eb_�x)�����^�����e�ܞ~�-��9�J��'�W��U��~���!{ўՓ��:�N;E�v���C_r擾T��l	��f_���e�fs��H8� �v�"��iJ^��`U
���#����3\Ab�<�8o�Hg�>�"�Sk�Q	˳{9?��Y].".O���3,|������7N�+�-�x�E޴Z�g�VE]�dA���� υ��8F���@��Ȃ�>�㪰:d�/4���8eZ�[�S��j�~�O��}�b�@�Lq��d5	 ���2!˩����*S��Z�i�L"��`2N�w�+.0`?U�	C�J�D��ȳ���o�H��M�y�1���v��)E��/����,���?N�/ko~�ڳ~J�/He��Ǩ�g���f�W���S%v�?#�d���������X�5��7�Z;
z�IM�M���a%�μ{��NӇ?���xn���J��z�� ���3)��Sc�ӼU���qo���~RC�#�gǕ"�LN�J]�C���+zj���/�f��t�@�վ�9&V]�a���JH��dp�E�Um\��V��ZJ�D9�#*���_y-cD���5w��R� X.��ʾy���Z��/L���#W��G����-���l# �9��pT)F]�Rn(��<5����l�������<�|�O
3zF���qc��91|lY�թ��p�,�,�� M2��%1]���A�`sBP��}U�O�4;�	<Y�U�/���~��Y�q7�g�?��� %�_��c��T����q	䘴��-6��f�f�D��b�1	��S����p%�+(4��r�i�V���"�vq������y�~i�,�i@�����b�ְ٘�9hP"��L�"�#�qKk5��'q���n긩�]�P��S�Gm�g�Sw���FIO2|u�=�x�Mͤ+K���^ �YY�`�D��W0v񗍂�!?�4-��>�6;���xLN�8�Y����X@������x��}�ī���&;#�D��o-޽��\�F�y�S�"�3��Q��::�UW��f4�b��&�n�1�l��a����e8r6�޼��8��&e�3�S^j*ǫ�j�*4�p�)�jQ`�_����p�=�����~[+�|Y��l��U j8�g�8x4������ͣ��F�w:7���-�?���f��40���������]8��L�A�$z��x؇P���׶�@�F�1B��HB�*���d���pg"��=��)q[�EF�YԖn�|ܾDnܢ�l�Fc!!�6��dC!��v�j�?�M4�;�H�Lf-�]���8cA��C����_�~B��rF���/<F��@���ڂ*��ձ��>=1+Ȩ�������E]'��W�M%'�Z=]�����#�lWZ�0Zvm	Il�c�F�X�q�7X+mC�n��;��sGC�� �X�v���Ze0�i�%]	��/w$$�;�M�f꺽��*]}��}e8>���U�p"n���R����{6o��:3��6,�1\BW.[����������ςk"
����f�-�B�U�s�o�s6�/�O�QU���`��
�V
Q�Ngר������E�̠��e�n8/�t�d��6���%�kA��o��<�	9���)-��` "
Sx�=���9+���1��E�N�	DCӪk��g��ԇ~�u�%(o`N�Y�M9\�*�'' � &��8�}�p˱Tі��&É|�6.�k�<4c��&N�Oܱ��ϧ�p��3��A8�/��9E��vO.̏�9
��u���jH�d�$zE�ٵ��:Am	S�T&��wA�V�i�Pp�v�@�J>H��*A�2?b:���%���zP��� /����8��Y�<ww���&"����`���5����r�J�M����@�(kqa�4E��Tqn�mҳy!�n�p%���z	�@n��OP��k����Kw8�C��g'����/����/,�m<�����>�eAfM�~��E5�3��1#e�N�J#���U\���3�� |[s����$wjL8��r2w�$lD���Sق�-��	'm��ˬ#M�iJ"i��I��>��[�Hh��<j�U����x�oj����Y�!L��~���ϒ�C-���0����n��Ĺ����jD��- C�x�b�j��+���mg�bBۨw��8�st��$`��x)�����!�.�*:nAQ���k��Ma�Ō�rN� �w���7���l���>�2�k� �� ����Ʈ~G(����b�K�IiJ�4ڟl҇�Fkq��ʛ.Y�q�3�p�!~7]��D��v�1�It�&���Gl0H=�2���%}c:����;l5����[ah�>3�ߓ}���`d�D%Ǜ� U�f�a�h$̲� C�p��z�[~�+�&�`�*�&I��6�,�O�`��W�{R�q�Pe�* U���3O�'=���N��<I�n�K�c�V{hHW!�_�`��su(p�5��	M���q�r��<�W`���T�̄2���a˚=���[N�c*
uĞ�X	9��y�u�[4Oz������o�j��Xݗ��H�G3�]~k�����5�
�e�\�M4:bӊ5C8@֖��~T� �>�Nqz!ye����V�� �"��!��c�Ij�
�4z�W.�ު��ӫ��:�c}�o�"������������(���|�ЙKOS��U^Fb�;e%��O3#�#���x�F�4�{p
>�����m[6B_�	i�%&J�����EDn��A�I+�s�%�������}X�y6b�\��,qoaT9G�`�h�2Co#����>�]M���r�W<�s$p�Zd�K����=_
{S��nZ���,�jh�&#{��GҨ����c��vFQ'v�U�����\)�k����f��y2߸�l���d�X���ẫ3mi�~+X��J�ge?c�-l'ُ��*����D���g��|G�4�q����;�������t�&�$���Ld�G*�f:��4��>)�8x�����	��:(Zb�}�����
tP�L4݁�$r'�B6��S�v�Ll���_�ّF�A$w_-��Dt[�3��< ���jy���D+/tt|�/��2W8!���α�q*bO�y��9��Qo�m�!��PQN���L[*� P���L�z
h:O}��(gPʊ�duA�����,4u�s0M�`���j������Q4~z��CwEmro/���C0��cJ���vu/#o��b*䪁E/cTq`瓱3��;0����L�"�6!�PA���\Ӳ`'dH��wٖYm��S1*qӉ��=<�~�8���0�l��^�H���BG/��)�6=�T��T�i������� ��1ӗ}�I�[pK<��H.����(��!�C����V���F�D2�s�)3�k�nĲ�n���3�+ŀ|�N����n��]s���2�jS�@|dO��U����Ƨ�'	%`'�/TaI�`��PR,��ĞӒS����|�<�XO����/jf�6:�M�/��(F6�˅ٺ7�uΐ���u��*��}K �\ z.ۓ�����ʞ����3_a�j6���1)�-Dw���CBx�5��J���=H�	Tj�1��T�NZ<�J��߃^i=+�l�+�ҍ�`����*����Q�F��U��'!�&Of@�_�Au�2"
_���l�4z��-��?��-,-�в��W?H"�������p�in��	�S�u����)6�eS[��ܨs�������w��gK�Z7�~&��<�8��X��^x!k�BV�}��6>an�����q�Y-?���&�)�Q�j���&�%m�[/=|Ob�vJ�H��5νX3�S���f����c�-�Ȍ�)�w��^���Ҿ*_��;��.*����9]�ࡐ�x0E4z
���llG��bo��<�����-~\-\�}�4rw[.��Ľte�H���v�9AC���6�u�8`�l�C4�3~�(!�%=J��z��H�t^K�����}�v�+w�&�Zi0?J3,��B�U���&؄T˙�WI�"�zR`�jh�H��p�@��j�6�����b�����ʟ}W��zUk�!���k�`+_w�g�0�K��]�g���5&��=~ѤLt�n8�����`he6m6`�V ��ࢍ�� ;ѯ�6=�hч%e�.�&�
�z�(5�oЊy��Y�AY��v��Zi��EC����̓��� Ru۾U��x{��j�6�A6H1�=�B������f��+��y�Em����p�nP�}0�s��֘ �4�@"UtyxCVy$1�+4}̳����U�O��rB�|h����HV+�l��\{,> ��Sjr�5�REَ�����4(b���K�7,J �K�
����w�}r8zJ5#�x���4L��}��{���gJ��$��f98|���h��H�=�h��qk�������9'਷$G���O;�_�������?�M2,�N�����<�
:�%�ҵg�w�W7��r�pr�p,\�����d�����6N_5I�Ԝ;�S��t~= he�t�����B�C�da���J��cլ\q����4H�o^CW5���
�^_� �-x,��L�)�	����`ˈ(�Qʂ���� �j����Kn-�*t>��|N�!�H�A����L��M��rl���}�]O�/R�wn�zg��^+�s���=�MJ��Mo糦7U<�`?|\��Z������g��~%J�ܶ�����S5�r��Fj�^!4�r�`��]ͬJ���-̚����U1�����˖"͏��cgIZ�[:eM��i��]�-9H�o��.�v,����6���C�ǅ,%�D��0�{L����8�E@[(���F+ z퀙z��C��G�{èT�ĥ��"����!�M���u[`6C)�� u	��i�w��,�d�a3��c:�S6���+3V���Pz�N�G4���n���)�zҾ؊���]�f7��A��┤�#S��5u:����a�r5/�V2hK��(�K(8S2j�ɸҝ�{�/+��T���7������,0����e�f�� *t�kjx3�#ԡˁ��&ۆ��'��ؑ�oܞK_��*A�S�;�'��4�׸�w�*ЪG��W��K}�������Uzц�8�Yȗ���AȨ���~�@�4m���k� �N����hN5��}rk]}_al��ܢ��8��"��|�����=0��v��@�*Oa!��pC�G�8 �d3P}����x�R���٤;^u�KL�ې��x��cB�;����Ǥ��P�c�Bp���ˑ�p[�<8�Ā��N7�4� c�L������1���Pk~���0H�bU���ʪ��?;n;���y�
I_+�8R���@Y�l�2��=І.�.�;Y�ΑMV�&/R�����y�v��:��A�=��QN$��ۋe�I���=V�2�gV�	|5� �V�󶻂&��I��37F3�fbT�4�esm�ʺ��o�Ǵ���#Gj�7�a+lt�U�P���y���.�Yt=��Bn,H�j�l��5�H��dS��\���^���m/ ���N���2�{Q��ݎlFɷ	�h=�}�� mq��\���0��|o-��^#��d���qu� �)�*sM�d/?0ބ��Ucꨴ�m�՚���n�J�jf���˸xD����h�P�;��{�V�חr�F��&�%=^��ɪY:�D1eJ��L��"���y"Ɵ�K�D�yݘ;�="���`O4�}e�b���ؑ��?�	4��:�b�z�L�L_�qD��"Z`�F�^�xt��@(1���+����o��ܐz(9�̼�'��[�Q�� d���][oN�08Q���PR3�s��[��Jzb�lX�y� ���N�'(m9�߽���l[
����1�a����-��<�Z�7�Ď����_}o����!�%Q�&k��HUx��w��<��xe���U��� F/�+�ǘ�_����������c�0L��h���<k��o�(�إ���κ[��1�\l�v�#s!o��\R���O��\��6F�Fⱛ��{>��U� ɸE����P����#�H�EpƑ=�����Ǚc(��1�?�Q��Y;�A�� �]�=��UP���,z��Һ��&+�>�6�X�ݧ%Y�Y;�8ɴzyڶ/c��0N���A"���ML�ݙ Tex�'b+_���P�E���#L^�+��s�A��H�:: �	���[��(٧ɬ@x�)WO�TO���q����w^Ń��f�M[�����[��9�S�ٹ��r�AӍj����h_F�Ͽ:�e���5�C�R�P���潚i��[1��7,�q4��xc���EX�#oӲ*Ȯ��Z]���dԴ� R��V�=������a���
缸���{���+~�V�t>`DvEQШ&�P-��\����z"��T�2�OA��1����K�Q���Ayꍿ*A��c-�)�e� �T�I�(�8uIk"\�<�����Y��E%���g��]�����I�,���S�?�79��JĢ�/؄j��9����oq&=Ō��#b�bq���:�g�q��խ��>DӴ	�JF�GQ1(�_ǌ.���g�x[	�a�K�r��L`��d
j˽�]��u@��j_"���1�n�݈�#'1�:P��8�K��ygX$�}	��
�2y���Ya����p��L��n5q���/�ų�����*@kTl_h�2
o��/z�д~U�I΋��da �e�6H^����[ee�fr5 �I��d�t,l�]t=`�=��qh���p+@�ǆ�[} �&��a�@��=/�iܪW�V�(��w�/ji�Ur"��W@����X��T�s��β������[��7��(��#�e����b�3������6>9�'O�<��&7ԱR�7H�|@w$xy�:�Wi`���"�)�RVSĀу��l�Q�����s'�Y���l�"%��Ȏ��|�)�0��#��haEC�-�R>�:+̡���u�X:�'ȉm�����3O��#+S�o���6'�
|J�|�)*�T��CּVd FΗ�� k�жT�R�K�����L_���TW���O$�~��I�x��{EU*�t�	��:����Q��?����Os��_j ϐB�)}�k�}mec��9p��MrꯚN��Df����h�6�?�ܡHf��m����9�^G�I+G�gw�(�i�����)�ŌpGx��{5;N���e�s�����_8�H��F�Fi���O�2fV�btz[�A��=�aRf.�L*K�ȀK�0ѼCw;���p&�Q�9�t��m_��W�C��)<�=��r`���!:� g���'b	8����γ�y���3P==\x2]��[�8N�֘�8-)�Fv�L0�."�6������8?/�l����k��)8��ԓ�$�{'6ח�� �j�RBf�.���Z�'�m�F�ՌrT��1��"���׼ɑ��(�0�vh-l����c���g|�j$�r��
�t�l56|��&j7�!��k�]�̱���J��8� � Z��L���م�kb���]%)��>�]��6�UU�"� ��9�2��+ʭCuE��*I�T��(�;?)�z����*��N���"�;�d�x���O�'����x��=�Rl@�������R�*���=! +��%ی�[L�Do�r��	�
��H��Vpao�	]���T�r5 GKj�Z�mZ����(�wʸ� �C:*T%T]�P2KX꺣��&V��ћ��^���Ho�a�������:fl��hM�>��ڏ&L�*��7>��݁�b*�}�Ib��!8�y���|���cY�_�T�Mw�HW�f|�Wh�̪d�;��fv�c�DZ�M��3��T3�$� ��3莰�̝g;�*���D�N��L��VE��*~
��v_�>S�W�u�պ^��%� j��W-4�	;R�/�.�_����۴�w��:��꽿��k�E�x�n�5|�v����
sc�+��+}rY8q�U+�1h_�Ee�6�����95(w�8С���qk��˱$eYQ)�k�����|MFZ8��ҩ�E�����wdl]q���υ�����e$���ۗ�Y�c�C��qp!"'��5<���.����s�M�:�R�Y�H���
Uٍ�d.�r(�3�f�)ˤo\+j(�}��6{[��ٲ޻�
lV�
/��l$��6ʧ��2:��Rݭ�����ȑw�_nd�?�Ӱ�Z�(.l2�9(M��M�db�g �Z)~Jk��l�rò��?�\�AJ��-�F#��[�,̬����I��)���^	�J�F|�H'2�p�P�Z��IO�5�ЙA�z����)����N�`�k��25s�0
�P��s��=W.���`_�B/�|���:jLF]Q!����=z��Z^bڭ|��FI5w�d�¤�E�¦Q܎���ԭ���<˴�a#�-+S}�r�V�!$J���);�o�<���$���s��8AU9��N(QΒ;Y�[�p�On��["ۍ�}�xO��x�����LC>ul@A{�6)gxJ�Ẃ�Z�7��H���z#N	�,`�-9p�m�ix��:p����x���"ę��e%{W,gZ%�*<_4���>�b�9b,CXGf,�����ZH9�s���O3X�BD��X@�8��ߙ�ϊ�G�b�2yp1�mßl�)��<5	>@^c/� e�� .u6�4�Z�;�m��'������u����D��������Opb�~�hk��}9[�S��-���:z��.cw+�R4ۿ,؉�{����	�J ��ÊC�d���6;���g\R�l7	�~ �*c��zx7�������_�,��O$GN�Y�L�+e�φW�Gy�{�Y�a��F�G��" v�5�IKd2�@q����ѽ�n�)WȺCO w4^�Eo)����^�C�^<��I��k��������s�]�l�L��+g�����}ֿ�Qq]i�z5�C]�r8���'��2��i����s�r������'�aAGR�1"���
��ƴ�����:�jt܉�0�@;e"��G�w�A�+�V:�(T������4���;cKN�$��ȥ����T}��j7�8�`�`��"R�o�h��"��ha݇�uDu�a�] �?��]:qz�MMY�)�������o4(?��X/�i��z�20���gL������]1tR��z���1|������`\��Z@��Df�{���F�Jp�����d�����NC_��K��)v���M���`�;�p�)uLZ���sEP�(�l���|��WX9���?�m��t�x��QG�^"�\��Y��xOzg"P�@���;�ħ=�0�AT࿱�[���uߌu]6[��d��eG��K��ۧr�>��1���>	��Zg��!��:.N���J��.�����5��ډ|3�����Z��uEK%G���ܑfŁq�+��	����ٮ�]�(�M)1�����b��g�\ƻe�Kj���>��"�kg�r�C�����9�������M�'p�,U�ER4a�Y:Sq�S��ǩyc��c��ף�>U�/���8b�%0V�� ��A!�Q�M�ǁ����$bRF�ߪ�dL��-(�lc"O�'��������>%��k�I��
�o������=pA�^���%j����Ōs��1�WJ%�L�cd;z��'`�	�e���lb�f��;�#���&��Pi̇yE��G����]��.�E8Ձ�19�~:��ن�ɨ��f�M��qGR�P�o�E.g?�Ϲ�>�"Q�
�����G���>�(�BA�_%��/�?ڿA4k�9��ۓi����J���y�*�0��g��_WT��<�5G-�W=U^��i~-�p>�Q�-�*&a:�ҏ���'�y�"tI���)��}�)A���.���2����k�-�p��6�K���Ԙr2y�����T~�.
�+_�x��X��\:Jq}�=�O�Z�B=K̀���܀�]��t��C�υ.֤X��]	{��'��F�� �5�Ϫ$���I�Y�	��N����\]c��qNϓ3��Zt�Pg^�Dg�fI'}���m�JY�����Z=(��ye�ݣi+(�۟�(�K��Yt2M�ؘ��H�K7~9���̻D�ͷ*_&Ta�qv$���C�t�k��L�_P��V��O>1��k�yp��^��Q��˿?F��n�6�j�Y� wH�s����݄\� D� �b�3�TA�[�$=/��,Z��K�f1���?�O�Nڗ��{����iM�e^�Zt, Q�1H
��ἸXR�E|����J��0Z�u7Q=�<��e۱��M�[r���D�`�%f5 gF��E�Y��J,̭@�s�Ij<׋�5�u(���y�**q�+!���B0����{bP�}
�f�˫�]$����"[m������E����؏���՟�RsW9�'�y���DgsL;�[u�W�=��(_Vj	U_��l�Є���1��\��'}����B�N�tҥ���a���������Z�Z~����`�Iu���&�h���F�w�#&�1�xi�� Kǯ2<R��zɜ���+����,���l���ؒ;'V��ݵ��S�$�An�c�1��Õje�I-f�v�e���"��t�Ht����Vp�A:mݝ�61=�
������x?�y�y�
oH�/XY����\��h���y(���Uo1*N	fi��X��ͨ�]�8�e����YG
�z � �
/}��rN6K,���19�	Z�w|�s0�=B�+��
�7�պ�9��^�d�'5�躦$����r�C��oc���L��v��"�ٰw�����Y`cb��0�S��j6)n՜����;7d��0�F!%Q@>��[�q��S~фZ�왨�-�v ´)����떦;nI�~�F�u�TX	���,I;�n`\J6]!��߽�ؗ��e9���C+H�&�1_C����P���Zr)�?����(�A6q�	�uJW
�MD��w�0d.ܷ;9ע�����|�A�^���7cE�^I'���@"�Q����F&z����WZ
�����c��SD���d�ɖ�Ș�c��������$�o�#�;//P�8Bn�T��6�sJ��&�g�Zn"(���;�:��������2-ܕ <�|�K8.:Qv��=Y��l{�m��i�=u?{[��^ߋ��Ǜ�)��@�Iˋ[H�F������AF
��C{P.c���c�8Υ�;�T�jJS.�y�F|Ÿ�����Ƶ��Q�cZ���E�el�(����$�òӏZRN���˦��K�e��9���ى2��E�grAo&?T�Ʊ��=�H�R���2sq��Q�а��L�OB�0��1A�2E���?*+�ҡj�=�{�!�݈�?�$��ͭ��y{U��K�of��˭�g�N�'<C��P̈́�}B�D�������xbYI���S��Z­
~p[p�x���y�J1)����F��jv����JefW�O��h:X�YZC��n#�rc�R���Vp�``��@}w}�kʲ���B`��e������ �uaQ�;u��p�֫�@�#&(T�N$$ɕ�wo��ߜ]GΦ������73�Q�u�s5�v+}�Vlm���r�ɱ�/�Rb1���ﴊ�Jz�ȿ/0pП�4�
�@������3%��O�@���b�%�u�kTWQ���A����2���x3�Ec��G��D�Wf+���� ތz$��=7ӊ՜���^-4O���D�M�B��?�O�����C�
]!��ٓʍR��C0&�*��U�v�z�L܋k��)�hi ���U��H	k3XW �E�B��E�.j>D��`~'ȣd	٠(���͘��Q��RHGo�]��� [�]g���rO�/���r��szPL沁;F|�M�IW��俌����o��!��ڜ��T��'D��<����U��NA {ϯ�'O�4�MC~�&Z^�|�L��^p��OVsgø�P ��%�������(����l��l�vm���h��|nK?wZ�F�žU��^p����u�j���x�@!��$�����;�(\f+
2����h��K1���?�fd�["�<n4�ͬ�b7����\w�-J^�L��M)�%��}ej_�o?V	�ҹ;^�q����:~ҏ%5��.�o:���9:���bZ�t$:qK��	m�tI��;�gj5�X���J�;����&�R�2��np?�Â܇���P�#F��5�q+خ��	�����6rt��ѝ��	M��%u���ϫ�۪��p`JκY�VVXD� m%�1�_�$@}�������"L�ϒ�L�.�6Y�2R�{�b�B���C�N+�3�m���>��|F�£b�K���(�/�z�:���}�5׭�2%�K�]V�3g���v�DG�(F3 ��8L��:�#x#e����+�����-)q�Y�� L�$B�P�WG���(�ճ���nC'����G�&1�����Qs�{����A��"j�YW|lP���b��r��i\�m�Eϱ��k�-��{�[�(��(ç��8�h�S?R�����!�f�2���iX[U���0 ���5�����Y`_��Df_p&w#~S�ߛ+�s��S����S���:w�I*Iu�RJK�,�7�Ԁ��)�F# ��%u[�y��ʨ�f����5�`����L+Z���:ZA#��)j� ��n�5�!�]�k7/W�S�D#� ��;#<�\�k8C�I����h@�'&��=�GԶ4����!��Aܤ��;��f�W��@iTm!���5%N���Z���Gɞ��*����Dp��^�!AV~�N�-�У� ��^�/�}����M���<(�ׂ�=�tB41�����:v�7�7e�>����`P�Q��:S���I�L����"ԥ�A�;[��b�5^H����_��#�������!�
���֘&�DJ���E��
�d��	�J�������o��{�xv>���4_���M#Ƞ��4����1<����A�-P���C��p�"������Z�I@�����G#ܰw�J+g���J�+3j��Y��V�� �Wꎖ�r�)� q`�W��6C�f�*Mp]� ,Yh�x]���K'�2e-�'�)�6z�5�@�\l�wQ�Jkh��H�f=:Iˆ�n�!vl,�����D�iG<;�q�(�L����cR}s�s R�x�l�uP�MxE�����<*Ŷ+��6	5����vpW�ӏ�qzkOb�y�J`�m*��`՘������@ތ�[�G�!o$q��>�ϝ��G?�Z��5;b����pHYl'.ZU�������-���t��4�]�	�	ؙ4��3�xΤK5�-�r
>k��?�����Б�P�<��k��>�I��P�GsH��pP�(�(��bC (;O��['�B8�~Iҋ&����b4��_��9@1��e�?ns��-G�U�ur珑^�.���~�xϦ;���&�V�����f��JɈ8��{��oq�n�,��+
X�֙F8�8���)���bb>ص�P�<9�₸F�4?\��mL�+ʒ�췯e;r֮���~M32��l|�[K���8I4���&٬)�=m���ſi��v����g`�&řc�k�1i��b����DP�R�f�&�q�:�@�Jn�J�x4EJ�=�mYk*S�ح*����2�-�A3���n����/�)��kMy�G�6>��	�^Ԑ�q�F`x�6E���(⚾��)Z$���,�Μm2nz����Ib^�����=��)��S)"���ŀ�m6:�@9f�dc"Zt�t�<y��_\g���<�'�������V�n�N�gG�n��@V��j�4e��S�5�@Yf[�Տ�X�`�����f�
��w�	/G�"�6�*��-	��dVĮ��O/�������]�[J��d���o�n^ѷp����P�b��`���J�1<�(�)�fq�h�P��ĺ
!1�)E��>FS�
��hq�@5Q�6�ۼѯ���*���T�8� ��y4f�S����Oq_S ��7���s��yxdƸq�E�=�1��6?��Q0��O���Ee�����C�&�� ���3� ����I�r��/[�2ph�Iw#��W@쁐��E��0�}�É�[\k��(���I���Y���>�h���$��x������)&p�â)<��5�D�-k�vt�M���Y���E�JBZf2���ǵTODH�NҬ�*��1��î�n����J����W�Y�de���u;���g��6=�j��M�M�!�6��0)яsW���Ҏ���lGL�F�W��\���γ@�Y!�G��_�Z%Ra���S��Z�^��5�M�	>�E��jV@�v�V��ܸ>P��h��58k�J��"�_n�� �a��G�Wr{[����0\W�;;�"��7��q(�<��Ԁ��c���1kf=����O��KZ��-��X�o�R^ͱ7{���!�[������#~�!����������&SAfM�#y��7�8�5[�[b�����=&�ҼQ�{�J�Q�@~j唅�s�?u�Z¡�Y�����\~f~e[Ac�w�;A|�%Ų2K]�Ȗ!���=������޲/l�qWio�%k�r����$���Ă|g95�C������W�5�d�E`E�2�mV�Q��z"����CX5�z�d��B4\�����-Nɕ�7߳�2��f���W�Ja*o�d��H��]�-���;��7�M�e.:t�&��V�RX�5��L����~�;���BV�`9������K�f���o�����z7`tS(mj��-� e�
��~\�1,�;:��>�k]WڤN�Ko�����x�q�
ո�d,�+�O6Ǽv�E����Ӂ 1��z̔�^����\�1 Xu�f��j��0Fa��o�X�+�����.;i�w(nk���S��}���?\���������Z�$�h�(+}���@AI���S6�@����7����4j<ODN�`d)���V=RX�`2��ա6�Nomt��O^��P2Υ�K�������J�ʑ?ˋ�k��H�W\aY�w���(?�5�<@��jJ�� ���N6�Ɛ&����
��5Z���
r��@�+3P�,��p,�h�(>_��OIrp�)��uw�f�!$"8������y�7"EfJ�C��\S�R�2Y��^����K��4g!+�|�w#1:�`ek��eV7�YOO�pj^ઇ��c�@y15Kv�+�֖*�22�9�+��;����y���҉�1#�
1�3�n?_�{�a�2���?�~�&�gӆ3�ln�%͌Q�`�g���g*��FL��"�W�L���r��C�ڛ9�W)���$�	���f��ۘ�������u�&��=���������Ag�ջ�H�6��f��s�i��%V��Y�+����h@|Ks|���4�2�|�fL����q�j���:&n?�TQ��L=7���rH�Z��b���B��x 㣰GQf8��$��Wr��@��n8B$��c��?� �0�&V&��4K��G�7J�ǛK��)Ǆ�W��q?�	�Γ;e�ʀ�Cg�j��*���_}1�N%ލ \��p�341P��)�!� �C��)8��o���o�X�3�x�4�O�4���_�;?���lT������hW7hkɋ���&{7�D���B�fVu~^B��q'�o���T�@В��
}�J+{��ʏc��{���l
�����Ak+�i ��	�֓��к�r5�������ƪe���{3����L0�u�(�&Xǩʽ�0A��
�
Z��Xh�|Q�_p�k�NG�`�k\tl�|
r���[��>�b������z�\}�?S2���r#����ax�%�-_�� =)Hi�8����2���ڟ���<O�ѽ����"l��lBQ���r,v<���]�ÿ���7�E���<�ڇ~�@��8g ~�1�m1��|��wY�m��Eeނ��R�5�������ӿ����|
����G4/�]6%�H��.�"��ܞjao-����_j�0�D��+X@1S���xVZcW��yv����x�q��o�?bx�� [%��ƌ[���f׼�NN`�/z�=,(���K��c��;�N�c�Y�}��	�^���b4#:���Oێ���CSI�f�X
A�A�uuW�mh������@$����na�Y6��`N����'�>n�у�U�~�`�Mu ���L(��÷��ըb��h��{�3F�PA���Ґ��G��r����6؋I������b�[S�`8�w�K��)Q���1�<�|��R��%�X�8n���3J2;Y���6�����i+�F��Ŏ<0aSXe�?>V�,h�*qb������Z��A`CJ� �>��9R�ps����:V׵ʲhbN�߱��̘9&;�!`zR3Px;*~��} %�R��p��$	Lz�G�낹�M�=qv504�/�-�O6ǖo׀�x�]��ԐLA��m������.7bd��"�O��������w� ��R�!E���\'�P_�������=ol��t��և+~!W��Kp+'�I�|�ݗ��� M�����p��J�P�w��A�@/f~J���N��|��)H� F����8�����F?���]����Jg#���4KS|��}'�S@��N\S]c�9�Ұc5���v.>��c�C+�;�Z�f���P2@�D
M���OAV�	�bĀ�Sr|1���u�ͶK�C`�-��>�u��Q���>��Xa�C�x��IJ�/t�da�$>BjAڐe8�<���-WTs;�r����_Jp�k���+BQ�
��Q[@��Mjs����1���k���W��P1�\f\d� .�EP�鬶���� ,�
�5�~���Y=�\��twwC��r䴪Q����c��d���W0�v�$V�����%DƩ��M��	[k��xU��
e2�����W��ؚ��?�*;�o3z��6R�h��eYq5x�E�'��â신��,=ڊ�y|�W�V&4��w��VSܸHm�U����Ih��9�q�v��.�F���?g�+���.N"�}N� ��4VR+�.	q���������e%p�M�h7O�
c�͗��+O���WrLt#9b�`����z�W����k��3�����������XK����2�X~B}(����\�䜔X5U�#�f|A!�݁�/��$��x��\bȴ�K�[`�,���]���u��]�L(�%� ��	q���v!���^�<>��{��͜�w����U��h��c���qt;��C�[8��s�6k����ȄD��n�=�fx��YX"�-��:�����˒�e�^��ʉ$�S2�S�_OA�9��iԍAO�/���h��F1,��}���}��u&��������T�.���2�ʧ�a�:����\�Y��\A�g�;ߧ�rb�� �e���0@�yٹ������z���
�?P���h1�|��r����b�5W�W���H+�:�+Ŕ׶������ғ�+p<nm����د�aVc����?)A�n;��Ӫ�-�����0)}��$b���@���G�Ѣ����+n��������F}�k[r�����Yz2�.B]��e<��<Ņ��I�y�G�C�wj�g1�𗚤��ߞ�'E+f�Oyz,,7qF}N�PӇ#��jv�����m�.����}�b_��4�My&jc�r�F�]���B�h�[����r��1�Q��i��7̲�pݍd')++r�m!;�5ݻU�2�P�\������_�Rpe6�E���ųà��M����$G{X��[������E��
Ĉ�4�F���k�7H�aSv��#���j<WB"���P.
�n�n�+��Ϟ`�$˺�,)��B����c��2���Sܕ*u�7�Ss~
&�@d�V�2�{�EO}]�/rM�ͭ�,.2��o��C�����7��6k?�R�w����8��nb�M��1"���/� 
���%�Q�_��5{]Ư�>�x�8)W�Ebw.;g�G�qY�V����M�K[��gOx��Q�/�&���B�F,����>FJU���5ߥ
X�̃Q)����@�@�N<00�MLQn+��h+�0����x{����3v7���"��S_%��Ņ�� L�hd�O߁���s6����%�nY��y��r�#�}�g���C���;�����9
DӸE=���b���n�#�rg}���>K�A��mpC���v�kAj�k������,Ŋ�9�,�c�I������� �-���Dٍ�/9v̯����x���P��1{"�(��Ԡ�ߦ��,L|$�G�$x�]+.#F^b�G�7�L�8O���
��k��R��D�:!�=�N�T���9%ߟuT�h#:ZG����"A�L��6����#�*ڟ����s�^5�V�>����T�/zOAP��6���[�C�(E�J��3� g}���(ҟ�O'g�I~��9�D.�WoWn�Z��#0�#I'���5��F��oވ�����%�ۙ]
���u�iX�`æط۲]9?|tJ�-��g)�v$3)���������)��F�
���m���N��-�����ñ[r��P3�,8z�T�c��Ն�~�L�Ԕ�t��_��[��d�M���n����p)V�E����L�2"�}ȑHwk�^�4$z�D��B"��o\�Y���<]�r3k=[z�s��!#���|�}W,��B�|7���Ё�/�]p�
*Xy�d�4A��$� ��X��Z(۩2UW;AHP|�1e�G��L��IHj��:\A����]>ɡ#����{�g��KrJ5w�ra��kA�!2�wW;�=/�4�Y��J��bǳ�;�r���˹	�|��rs�L�י�жp��mH��v�L
���[��/�>���ތz��b5@�zZδq#T����tn�a8#��6x�[�����2��x}������[�z��#�1��U2`�Wa�Cl#j���v�3Dz�>tB=]��
���+����96���C��F�w��W�;:� Ep��ހ�܅g�U��2n���d����(;�k�`�dA!�m�ux�=�)�NVt��&�붾O�5�1�r�L�w.��W�l��;^�:�])"�;,m��*�"��
"���w����Q��)�ԟ�n��f����[l�S��a����В9�֦iO{haK:+�Gz���J�L�`�!�3l���$"�T���Ò��zP;��{��3���)"E�"�v�@��lU�=|� O��fW��&_ۧ��%���A�,f�	)K��Q�숖M��b�t�|�$,"�t÷z�P�f^�}�*n�[!��������<�y$��5�`9y٢������z��+�.�E�ϔZ$�Qa0��~����uY���Xe���U�~͗�9ߙ��Qq!�3�X��.2c�f����u�0����B�"$��#r����)���}�;vU��Q�	Agf/)bqM�o�K��G�(�m�G��Oό�8r2��%��4��^G�j���	�i�H��@1�r��9��;����r�+�cf��̣|D!�#��qT��*"qp�hNs��Pk����+�ߴ��ٟ�CܘL%��}>�KM�� m�
P�&����h,(�,�q���o�����ϑRg�<
��-��+`����b�8���\`�ɢ[�@�^�B�����{�w��]���\
;V�!|9���!���@T���z�D$_�i4C�wU�&��Ѕgn��Vny�  �1�!N���
S�b�[�S�],��H^Z��"��X�v���o�W\�gIM��绔����VA��o����Lv�~E�3�a�����ouh��w�n�^�HBQ�k4��u�W�fY�L����Q\Aa< c2��H�dz{o8u 9�4���:�k(t0p0y��lx@c0�o�u�ܞ�t?�xҥ��lS�n����6��l�|��g�C�í�b���B'����A�v5�����ߦј�>�1�㞈��R��������&!o���Yp�ʸa��=p��5b�+�^nѧ�v��cF�L�f;H1�� �"�*�<�Oԗ)yv�*������"qD�j.G����z��6@cCV0cfpYrfq}5�qV��ʍA��R[�����38�J���rFz����^�Ӷ��r,����ϩƌ���Y\����Υ�ۍ�?�V�V�rj�:Iu]	��HB�5��L=ٺض�R�(;}�X��_��jݕ^�v�L�����6�����1h��]_������d�������P^�XH(��)e$��qDN<�N�tW�>��Κ�?��@ʻ��Iɭ���[[>U������f<T�)�Ɇ� �i S�{RX)��J'z5�e
զ���D��]e*�g�Szd���c��ͤ'Y�Q´����VG�BsG@ 	������\��x�YGM[�%(ѷ�ԝEcJ��M�����f({IQ� ����g��a�1�q�+Ks�9e��I4��^-�ȡ��t�]���W��m���=����VݐN��jŗ�{����֚�ȫ�>(��H'N�J��Xs-���/�Ƥ�8�"ɍk� �y n�6� n�jNՃ�Z7M-�B,�z{.h�3i���_�d�A�e�_J�arj�$+ 8�T=>�Ð1.^I��~�H蘢��L�W���:�H�aSE���F	
��b	F(��ŹP�w���]r:h@a���ٖV�h�b :u(>͹�dU1�C@�
�O�QҌ/{�4VZ2فw��_�;�u�K<z=�L�'4��w������|�^I|6L�Z�� �Ab����>ѓ.���0~Z��I׾���{�4�E��U��J �n×��< S����#^^,�b��?�:�+�y
/�,ɴO�^�|u���g_$(���JC�j�*�輓ݡw�UV�Pn$��5x�5�ty��k�s �a1�
��i�g��i5����lՃ+&���S,+�+O�hN��94������8��k'�W�, H6�c�^0A#���_�d�z7�rx4����=�5o���m�Z"��6��jӊen�H9�d�\{t�(����mؠPK�gS�/�z�Ֆr�VPV�����n���;-�q��M"ޙ�i3��5/�ESq�W��L���