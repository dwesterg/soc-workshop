��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t����z�2w��0W��B'Ԉ�h@��Z3���[�l�jP���d�+C+G��x{���ӯL��i�+����������z�B�(+���B)�/Y�#x�����yP�8w��1�����P��c�%�/�~�k��p�eݍ��wa��؀��`i�%KL���8����h�vI�ȃ�SMR䙼���,���9�7��K4+�ΊxscK�4|g�|ed2EjO��+��}�����i�?�	����M�>'Yt�cܵ�>Z�T�N�x@���h��+��PO#�� �������/��]�!���܁���.���HB%��O����Q�ط��,MA���-s�a�Am��_�v�%E ��a�MG���Dl�nqF���Pu�8���:�+��C��_�T�1��G�v\"%'�+PC*�C�u�U8 ��Va_:��z�(|Qb6=���NT;��엽�%���d����ψ�Y��\��J����"���?��pv�	�$�^�<��Pd.��#}�B%����e�	+bcY$��ձHk�Ȕ�Fĭ�}�cZp���ܭ��N��̾�bOt��503S�;�-�6������M�{4�̒R��ȑ���ڎ����ޤ�@z80i�@V�y��fYh�������rGN
r�w��L�4V�'�폊�{ �}�'�������6��J�I����q�I�	���8�.�s�:8lL�3}vD��P�hc7M�ɕfk�E�y*'��+�E磴���H�E1Xk{�9R��v����~˪9��KK���\�`�L!Em��S��%��!7�$ˉ��X%\�������zvH�_��αƃ� 39�l#��L��_�'-p���^�D[AqMUMO]1%�@��\�UY74��m7���0j�R��K��B�����!n`� ��Z��yN����?�L��پ^�h��h��k8�	J�H X�Z;X<�NAX�����N���ǎ{Cu��Y��Ds�G��Jr8̰�2���$S�+��aM�lW=^|�A<�}� x�B�q��O��2�	�c�޿�)�u2W��<�v����2!��[:���!�gdO��IPŒOy���K�Pn0��nH
�H� 0sg��Ʊ8�41`Z�E���P�~��`�^Pu���W�8�	���G�FW2K�s�8e�r�:Y�?"�?<
�Bw[=t��)X/��<��2�.O9Ɵ�2p����Џ�������()�(T*�2oZk���QPÃD��<h`�/�	^�ō�*���]|*��qȠ��I��"�F����� ��<��O)�Ad����7N��Z3�BZu���&�,4��}:G״�5ض���S)����5?��y�D7�i�u���Ę�څ#���y�,§�N��G�줁&/hB	�ӕ�`Vc`��;����ǿ�ǹY�U���ﰍ�UK����3��"�c�:t��\Z�0ڼ7����.��������F�-T�f���2��"q��ǩ�l�e���G�Z��\��([�)Kx�c���1����XK�0��;0�X��͖YN�AZL�}��Gơ�Mz6e�ԃ`u����E���/�u��o��)�O�2U�Kt7�0S6v�`��f�ֺ�f
��^��0�rT!M�S�)fY�������� �`��=]�PGCܡ��i~��A����7[U�2HL�s�
2}Sgc/Fs��cƇ�F�l�6�Z��U��y�b�QC)��Eo�_i�<�_�D�f��*f En�TЬ�r����;���e�k��A��i^}-���;H��e{�K5��8�2�2�,��2pvkqɜ�<�J$�	�=�0d�p��{���hB�b��5�L3C��*�/xߵ2���B�����#"����\��A}Y�pEޭ��P�֭ڒ*x���|��u���6�߽�1ɐ>�V7Y�K��~옕����O��!*�X�s�h�?��G�W�'��=*�3,�L�u�\y6��Y��3�3%y4M?�O1N�����<ٯ.�(�����U��!A��4Kd������������$�҇z���� �ں ct� /f��h�HY�w�]�8j�J�4	�a��(��l��Y�Ʈ��v����R*����h�<�^�g�ƒP!�w4Q�W����P�f�(e~�]}����ۦ��)೪�DR1�����cE���J�,E��=9W(��BaE�y?��
�l���g�g���j�S7�S:}~�!�0\��Ə�G�f&�fו���@,��gϋڜ�-��%8�֦c)�&��&���s� �x��Os�ɇ�Pr�y`W�x͈��N~aP�$ 3�<��I�߄�P�����9x�� �;����
Ҹc
鞯��T$�0��GO��:�?DK�=�i���"L��tґsl��`�Νl)(oNu�����q�6��v��e���}�@�����+.�L������y�ΒM�.X y���i�G̢�x�� ��O��eF;��0z>s���'�9_X`ʹD�Y��I3qvdO)�!o������ [�O��8�b������
�al:��K�(��.�ii=c˶v�JT-�U>�����wX,P�g4-z��Y���lҏ�~Vs8�����q�7��k7�d�cj�lkJo�N`��F�@�,c�V������da� ��!�k0ghy�P���ȑ���J6y�w�kR�>�"��a�`�3B,��J8���A�#澵�� Zл
���Ki��I˿�L�}յ�(Jk�'�j/�|�.�N�JB�����ӣ�}/YSJ%�����^S׌�����9��ɀ�@dN�HJ�7������A��Q���5;�g���9Pw� ��;��O�v�
��� i�k�%���gV�4&4(l�]����J`�UR0�����t5��xۦ]�DB�s�2��蹲��R��B��bx��.ԟdE1^X��
������4	��Eܠ��kݜ��`��,O�s�8�iEd�l�o���9B�Ra���h	�ż(�����=F�S�?~O�,oe�'o�^u�����K����
h#�N+����KDxS�l�\`�����)� ͝l;=��츺t,��	��=i�íX`T�[?����娩�;6���^`w���O�W�p��%�f�����X��U��Ԉ��Ә��u�^��L�l�����i<)������f��P΅�0��[/�1,��c�ݯ,m�A��Ɇ/Ԕ)<O��Ka���T���^}7ߠ�8#J��όEо��Ұ����l#ǅrG�o&mo��p#�)3Z�Ѧq�U����GJ��.]y@��u�O�،e��6r�֕�(��r�+�Ɲ�W��02�|��A�&��_��kz8T�]�*k7����6��x>7��H%n),�
EN�H�1������ɏ6��F�d��X�|��܅$lVܽպ�NO�*�|,Y�����d��H&�"Ӱ�~���hh�<�go���{��Sh��j��BOK�AԊ�V28?K���9#��Z��+y0?m5؆X*�E�3=��-H^?��V����)v�k�z��/�Z�_-F�k̮�O����&4��j���h=��A�;���WW�L�+G�5�qH1�
�	�������3�4�~�={[�����iC�v"r #�M<N�<���`>����X-�@���r��[D ����ͷ`!C�)��+y(g�Nr����'����;&�!�I~��`=ݐ��@���RГ��s�t��<k�k�1��۬EbA��;�F}*��[	�v������зN��L�d��=#�D_�7BvEU�	�_�s��m�I�k-PN��x����2c����*p4`���o�J���ƻAi�M!c{]9D�lE�^i��v��H��ɺY����6��Ƌ��E�_P���;��M�����-_K��e�0����Kc����by�j�d(��# g�^�KDtL�F�D�z+��k�c��*��u�<;U�S�J��'α"��`��o∉ԽsVH�@�	��Z9 W��j�2���§��8%aKG�s�q�Nj*�n���sr'���[���an��c}���M��K��m�m���9�Q�]~�s1��D!8_3n,�F�w�{��2l���e��)�%���+�����b���*t�;�띡�E7���X&����L�t]c�Wl��c��5®l`���ꚗA2�~nxh����9S�U6�/�ܲ@79��g[�FL�5_j�~��8'�lzn�m��ɼp�PMF�T�0��m�V���=��!Ac��7S��Q員W��aR��-.�w�-�kT�͊&��������[�v>�cl��j�#V�n�u��x�RHo6��5�1��o���uT�jᮇ�x�M&�D�S���$�Zp��� �&�/RPj�i�+�.�~k26<���'��n�����(�p��:�-}�̇�h�bܗ5[�IĂ�?�^@�
> s�I�&�a�X}����S�}�@87h�me��p�<t�/ciY�d����ʧ�w���X��)N�G~fVWc���U=�=��&3��9���5��YP����z<V�_��#�8�W��v�x3��eV���jt�{�Z+�����Gz�H[�I��ݻ%�b-�̊*�/]��%}�2�]�^����Ő@6�`;�=!�4�OWw��3N4#���mkOc/�y��s���8��l�Eۚ�JN�I�aΛw�_�s��L9i�T	>u�].�������i��R�:���>97����`��r8�v"�}2��"�ѻ�k��9��L�	�j�����q�Ѷ<X��2Ě{�M&�R��m��Hhb� ��j��@��]�m ��~%  2v�n�ߤ���vw[r�f���*�;�-d�ɤ�L4H'�H�H�4�;�A���^�j+�#�*9���޵��=�O��ef�X��{1{�*��LQY�椊[�TI���f�b)V���e]�qI��*����t�� �|�
'7�CT���sy�L���lnm	��ֱ
�� t�T�~�M�/)����G��
�5�ɝe��m�����c���N����b�K݅�26MK���h��ʜ;��@PM��^�(�J�2ay���Z��s[�Nd^���|�ep��'�h�nO���8�q��"ԛL���G", �=�1�k��-X0>���a�r���6�0uk/��;�ο��ԜU>~�4������#�n91*���$��N��O�
����WF�+����~(�����E�|�-%h�z��|.J$)�M��r��U�HJ��KRӌ�ɔ�ZX�XD�5~W@ۤo),,}�%�� �x`�f��y�#]V�|v�0"q�fʵP�b���s���Fe���Ĺ��m�
�K��(\�]U�(YA�Av�7�zN_m��\�]	�ToH���2[ ]f�E�ˏ���?��}O���&�vg�dVh
�s��n(S0<A���Qew^-J��ͦ�K�_?��2u?�f�_8�U����t������[�b\�����m����/��nA9n��J���u�>я<��<i�C7!t�I�{�6)N��SYn��[ V��m�D8g<ʣ�
o�;Sp��ȝ"����U�H�vw�F�$9?����k}D���O�|͢4�3"`_���U��i 4K������W�ܦ������P�9L+����ީ��#;��,]�"z����[���j�~)�7I~A4���d3�qbҲ�4����p���*�n�٭vi>��R���_��Ru�����ꇋ�u��8��n^Uk��E���Kr&t����D��d���Ȣ6��6�z)h�{��A}I��+lhps4�g�z,��S�� ]�rw����p�@�me�	�	�d̔c���lw�Y��� /��I�h��gg�tG��n�m�W(���:|;܌2Q������0�/�b
�>R�"HR�^"��4���h���Z[@j'd�4 װ���{�_�� ��8z1��PA�)� �yw����h��b`�H3�L[���Y�^�\�P��䬛T'V��d�szd��nۨ��BO}�M��̖Y�˾�ϋ��;���:c�0 M�cT�n��a�.��>��yh\2���+�ߠ�Z���ʬB��h��@ŋn>�_�2-"�`�2��'�8�П6�m�w��-������&"Q7���^�a��=��iCU��oF����ō�Y(=����S��aڧDvm�B�!���`�2��T�,J9rWj3q{���I+���`/i"�����G��z�$�i��j��D�C�~0]@R�Ş�\S��S_��5pތf�\�Ό0���Ԕ����ܬ~]���(6O��3-�]SK�ɗ�V㊥jp�64��s�Y�vE&�xB�h>��e ��������lu�;f�nu��D�4FG8T�]^�;� <�&���f؄kª�C���8���`��\+��:���e�Z�d� �a�d��֐7i�j���%�2��t�b;�L������{['!����"�����C�����4�(�k�/�We'/_=�I�ܹF9.�� ;�	�P�ޤ�����B{�Vs���z��ڔDwC�>[E�Rgƻ(�5�I���4�����"ʦ��,ٍ��ퟥ�����D'��!]Ɓ�ˤr��J^Ƅ�L�+�sq�+ʂ��C�Sc�4�>��K��\47|�?�Y����?ϐ�f���C���oC�I�ud�������K�ws!͸T�[��7"$�q�e)>M� ։5�̤+mmG���ľ�!��	�[^�S[{��K��E�Wn�H�'5�2�욗I@�z�<���3�X�=Oy��X������6�'�
�����Ԃt�sɟ(57������;�#���=Su��^Dog��ʗ��!xYA�C�[��V}������渒�%�o�aj� |� :�1��x��?%pRl�R�@2������S���A�`����Ǻg9F���h��X��N���h巢�]ީ�(}Uo�������ȫ�:B���)�4�w��1i)XJW�'ӫ��g�P�[b������5����w|��P�A(Nߎڿ%�2!� O6��YD���,���xͮ�dé�q�`ef�C��0�5����8Q�� huB
��*����zC8����e�x�|�g:A>¢�nGa"�d���G�x���o�/����-��S�^5�p(��qYj�z�5Z=%ײ�6�0T���c����Ž�ߵ	9����	��������Y9F�B1/��(��ea�C��q�����`7�K���u?LowXW��An�\�xz�n����O�,K��r���t7�П�oA��a��8un�y��	\��_#_�+�ks�!G����5�K+�Q��x�0i�x���)ʅ;�'�󪖗��b"�l�Mf<�<k&�q�ڋq��{�s�����;Mi�ZτӁy>������{����v�_˂�_�Som�d�#��Cɧ�"O��f��9�L�� ���5��i٤MY���ԉ���.��:�t���(a$�T�DwN�MzA��v;�D	$�ۃŨ�c#��kk�����x_{��m|ϱKp&L��zO�	F��7?���J��(z�ы�����%��~s�ƶM]c��q"v+"��}�1`��A���|��͐�ɯ��gX\˶!r��[�2���� ��[���K���~c�0����Oԫ�[n
�=:=+�bt��ˤ9��FS�{HA�����7W/+[�a���E�����ƒ�/���N^�ܠ�Y�'^�!��d�O�^�¾*H������r�m�4��)_�F��S�~4i������M����G/�Y&B��l!(�7��0���|]��B@4�Y�޼��r�^v�7���eQ:�'�	*$">0��1!6�J���5J��|)��qd��:=6d�u ��V8~�z�K���y�G����M[� Pi��hB��C��"�cu��r�m��*F��I�¥o���a������?��|�P����)��s$N���gUR���"J�Ө��9i*e0pqк`��]�wt񪧷�2�&g��s>_땂����7JR_�f]�����Pf��{Ԋ����?0��O�m�}����$ADT����d[�պ�|��3������F)�Ii� C(N���D4�Ԋ<^��/��H�Ϗ�H����^�!�L��u5U��>�P1qm=�De�)�t�hXkY@f��o�z��J�
�Sp������޸��AQ����Q�4@�����;h�$}����{�-R��`�.�j��+E���9�2���d0���6�b��T.d�E��}*��df��K�V��Z��s|ܐz�F�oWʹ�]N���YH��P�ܹ����U:��-�o���轗l,�ł�E�C���d�{�iI���u�wĮ6�%��EJ��pug�v�|�m��	\NT��*{��6 ��І+��
�ˎ��82�X�%�+���u�ʀTTy�t5�s� q