��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K����i���sFbu��:vc�s(Y�x6��"�K����0'�^y��/�����_����4 �"�����JF��N�)��[J_�K��	ϽZ$�\�_��ǽ�������v�z�[b�C�6�i��˳�6�ڀ3�2GXG�v���o�Zz��}7E�Üˈg 5���:MC��˕|�%�n0� g�yv����93��~_q���27�is�~��9DZ��vr���4��k��e2�l&jN��Rrԥ��̣�&	W�f�������e����K���_�o=��/�y�x���5���H7�nvo�AL֓_��-j�3���9(hEkH���$�u�|@��3��*do@cs�@�����{b�9.yCm�R�hM5�������9ҰM@'�����OR�F�n�h��n:�����R_ĺʡ&�/��y�i�ͥ��{����V����'tn�l�m��b�����F�?d�%�'�������M�T��w���̤�)m�7n�^�=��s�XZ�}>�̲�_ƏU��g�(��%w�P�R��Fz��#��&�q2��k�8��|��U����k���3Mj�C���DΈ��t��Fu�[��[ם=�m++4��V�1�^eh]=;�6�"��Y���H%��ܵ�L:�+Ju�!�E�e��_�z!�.��|,��
��e�������oĝ{�:��8Q�&t!�ҽ�>&��#��^�5�������"ʦ9K���~s�\�Y��&��"��#Z��j�<r��.��`K�I�{�j=Ǥ��<�z0{�|�yZsҔ�!�]�=Z^�h7�;sEni�!����������^�=M�~��C"�J�t��$F���[�X��4��8+Ҳ2��\��ņ��Fݫ�����!\#�ZNI�z��WΙ忨���DĬ�$ir
����1�)u@aO8�v��d��"]��<�M����(�s���\ %��9�p/j���myۿ�(�J����5���
?)�r_��"�3;<[�U�I ��S{m�F�H�:��i"���}|]��@z��F��2��^�9�܀!�x �F�=�/����{�4�Z�A2i^S֐��ׇ̨F_%��H%3�'r��ŝx`�Ù��l��KRi�꬚K�o��M�hXb�K�տE���d�_ ���i��H��������guq��ܾ��`��.&�YNw�J�."ͥ)�{���C;�P۹%�|v�B��ƴ�=7 ��u�X/y��*���`��Q�f�VE������k>��^1�ࡨ+�@�3�����Ž�&����>�8�%Rͳ�$t�WЙ({ʙ�zX�B(f4E7�z�\J��ߝ��7�B��C���8(���GR��E[�D6�MA�I�6�����i��뜘�+$c��1,I��O��st�q��"�i�Wj�}�PK�fnOwk֮����*ʹнo�	��HH�
�2TΎ�'��0�׊��5竬���:�Dr��M�QT�mo���7nmѾޛ`�2H4erŶݸ�"[�)�f��<"q��xFd�B��zb@������+�D�H����J�¯8�9ȹq �&h���C��飤pr�G�ٔh�"w]�I��t�@	m�]MT�)"�B�Vr�T�j��*C���6���̖�� m�RA hN�S!�7P�śUl�Q�*a�A]�I���r�r>t_�M~����#���:�4N�6�q0slY!_����Է_�Y�tr!䌇^���"�%�/�]��A�����_�-��O��~ojE���P��#M�;B�w3xl�Kh% W���>�k;�͎>��@�<����,[��^D��ql.�	�p�]�]2��w^�'=`�\��`b!����fA[��(��U-b����*cg2�Sc�\#༻l� R�l6r-Jt�7���A@CG, U���ax�?�J�-����8��)����i4�^\�)�!_�^�� �
!ӄ��TU��bA!�CJa�A�a��O� ����,�~�9� rzZj�G]�yO;n9���x�i�����'ZL/	��
2E��b�ԅa���,�hq��Y��+sU��gݎ�Q��m��_dz/�<�nC4C���˒k� �u�ꀿ�q���<���%�$�sR��It�$ '!ݵy�%ǎ�yf^ڮ��G[6j�����k����)�l|*^���hhҬ��'Kc6�"�4�P�*���v�<�F<��.�޽BXU|�5�z�oKP�\w�R㿿=B0� V��# *�I��ISZ��=?�r6�\'�f��C�]Tj���y��6e��	���hr��0<@�.ڥ8�T$A�p�,�L��h�/B���RA��6U@֬�jG���T~CP�`�,�`�-h<�h�-�!���R�5.%�7�I����&դ�}�+���7xJ����K���D	7IM
�\f��2I�V~������t�uV�-	oi�o���N�rۊ$��w?��VU�Y��������O4�WΔ��X�k�d��^�v�k�E��� "���v؄���28���K��g������Q�%A��p,�|��0;ܷ=ZsV��J��g���zmG����Q�����y_z]9��G�ﮉ�=ug ��_�7H[}������{�*:U�#jc�]ui{i�N ��u`�#� ��+񓔖aRqth-�Kcx�۝����,����B6�����)88N����Ѓ�l����,]r��)ޏ0�y�Y��VĜW�yU�ƾ(vn�(sL�Iƾ�e�fu�
=��a�+����}�D˝��F�7zg��-+��ڧԁ��&��&��%Y�:�I��b��:���)���wzɏth#�#��;u�VL8�;}�jj�L��q�rEsZ3��^�[�)Ncj�ъc���MK���������p+Qyy�_a�'P*�a?�6�T�Uo/x�U]�Py�'M��	����YM٤��IhP1��w"D��z�I�F����T�p��ߖ{�Z|��1�(_���xM��G���$�k��2QσLl��כ	��~N���,9cw2$+��'�d�ܿ��ЌK��6��L��&H���}��h�����\j/�!,-�M39M��껚���rJ�1
lږ�1wo1}��w�@��43��'����v�N��xNڇ��z�C��^GN��2�=��{�ҥ��oM\Z�Gη��S|�x��-')u��o��~��8A� ��X��1��t�;�O���?�n���-;��+�m����ߧ�є�>����^r�1��1<N��ξ�/��K��>L�q�1ڹ�Z�/ܤ|��ȷތ��r����?�Ѵ#��W%c�O����B��.Ll�n2��_}{sW9,c��f�|��{�kv_C��C�s�}�\6�
+/8�	�g��Sp��k[���p6z�7%�F�h�"[�t J3Q��5�	��9�r4_�ȣ�#�r9e��7��F2���ä���ѥM�Vy�%�T�VfmbX�fg��+�\L�\���c��F�W�>��}nJ�0w@"�n���L�w~��૸��6DȣDsY[�t-��p.2Q����8�ߧc�HDQ��]{m�UX�(���|���c�<���,}�Tł�,�'������z �2gr��&�?8j'�Ye�ꝱ�Cyo�����c��⫱��<��_���h(�S%,\o�v� l��Cq^ݜ@YT�H2���=Ƭ�8SA�i���A���x������> zM�%�tD���Աo���r��nPUb�Kfe��J���$�1Z�/�k�;�mI��qƯ�|ѹ�N����!7�3D6�<�B�p��K���}�V�N��u���g2ұ��(#B��m#u��<W!cO������)���6�
�nr�_<��b��Ք�)�/)z��9�8yy��|<��s8�^�(K_��B���b����7��������%��̨NBٴ0�82D����<�m�Н�b�h�Fd�"��ؽH��q�(���q�������ġ���}�4��e�����P)��L.`�H}62���=�R��4�@�ύa����s�|H�
�Fhs(OR�V(�2<	}k�;o�iC���B�>v����l�H�QA����N)XR������P��_�B+�M���s�j:I	N�h�t��m,7 ���ֵp��a*0��U��U�������Z=�U^T��"N�˳��n6S� �0�f��fR
�@)�I~��_E�容�;�o(�UJ�;���L^$����w#���0����m����.�L��u�R�n���8i$6�о���(Cd7��@^�|�����?�h�����8���(�w��6-�
�-l O��f
�<�N�)Z�E���CcW�#����v��ѧ҆�6I1�;Z�Y>	�0X�]-ݓ���1K�s�{�P#�B�2�l�z \�kw6�>._�dcO�ޗn?+�/}�<�&	`.K��>�1I����ٝZ�x ����i�HՆ'��� с9=%E~�e�>r���DrZ���De&$����9Oi��S��˧` `C�
ӬM���R�J���n��[��eD�/j�{6��%uY=���Q���3B����#������כ�9�s��QÊn��V��YtN}������L͠;�����C��W_c�F\�c�
�5�@i���Ƀ\��j0a��~����"�2p�A0җ��O�T�ʫ�a���R!vW��b�E�"$�R�k
�̐٣�l��p�O�Dk���T7eu�鯇�ץ1pp�	V:)����H�i������)A��)v�y��
�8��z(c������6���'�/Wz�?��f�o�b!�����b�W�[v"z�ei?�,�j�u�q�:
꾊�����������WqAg_�"XN�!PC`��m�uڳ3r�;��3'Kk{ ��]�$惪2��� @�k:(�XS������s���"�[Ƃ�SN�p��;"���v1��i¬��y^��������N�\�k9���9���'�L��V��&����EV�Q�LQ�m�A}�gdu�kUK׎XV���,�1��A�Y_��!4(��qҵ���ar0��d� �=4_k�6$�9��t�P@�sB+�]q�d{^[�|���О��íf�e$w�S�s�"�ݭ,@)G����Q�ʲ2�J6J%���`��|���D���2����xn�ϝ�۴a�,�yIc�\D��a>�qԽeYBoB�%�{7d|Mc@�A��Yp�X�c���o�!V�v�P��n)q�AF��AJ�����Q� �=�W^�N)��(��DB�%$�"��5��jq,ǯ�툰
�ma�Q���۠��r���ɮFv��2|��xԀ�B� �襫�4��	���:�N�������	[垶8��۠'k�]�T+m�d����CW��C�������,m�n���l�g�s-<r��)����Ϋ���G1~?({Ej�^;�ļc*@��]�1ߡ8|����e���g�_��iR������\�
����৖�eնK��=B���wE)���8f��	J!�K���^W������H1�t,�L��I�4��ߗ~�y3r��B�� _5�����0Beq��o�f��-�3(Qt��G�ÀU�Bs����z�8{����[��0:��E�N�Z� =;2���j�c_��ŀrё*M�$)�lɸG�'��D%���MN���K���A�k�;T�A�Y�̦n''��B���`fNǜ�k��S�o�ni��^	�a:1��s}l� ��?�uA���D$���u#���� |,��Z|�[Y�Y��+p����K�	���<�O6�qZPI�M��Uxޚ�Y�ݡ�4I����	�G )r��Ҵ�Z:�c���n����
o!к��x[�����C&^�y�=�|�m]��o"u�Nk�6�-W��j�)�K#�~���TD��t >�k7�!y��p��ex��=&C���D�3�F����(C���֐e����0NSb�f��7j��gd_��������܎z�Y��sg�F��V֜��ܝ�s�h��9m�3b�⽘�cG������eP ^Ѣ�K6Y��e�<yZ!-Au;�(�}�j����:�� �}�r[`��!�z�aIV�fl��0t ]��	������,��j���$іˬB�`?g�'�B�(�:�۟hF�?c��L0Ҡ��[S��g��T��fn�Ђ
��'������@���,�>4
�f��Q���ym��X�y~P�P���OF_�?\zU��V`�+�;u����S�*F$_!��˹}>� �Q.��DBnG�o�_�g0Za�+B*M��t[�;��ME`�i)��2u�I��Ͳ��jx�1H9���R�2��2��h��9��h��х�o펉M�tȷ�E�6�s(�5�n���C�Bj��W��
9�zn�4��eQi�x�,bt1,	ǆk�� IwN�N
�Aa�G�u�_�7piS
UisQ�w��s����='����t�2���.нl��TfB@F	4�+��:�?�<�B�n�2gb∫�H��ioڰH��X�T�!Œ�׊u��th�"�>Ɛu�>2I� �M�q�I5����%-�WjSR+�B�V��&��_�b�,�����>���A��H�>:�����!X��t�Ǽ���yE�56�7�#��7�b���/#lZ�[#e�ss�Yu���W]D��Ҁ��f��1�ͷ$(0��@y(��=�]����(����uzEǑ�J{p#�A���'��K�h��|�`��YNap���c�*o��������El�W��%x{�}E�O�	o=Z�[(�w?�Y��|�d��O��򵵍?�N�� ���c �6!vt�$�}'�AA��U�B��$��B^ �����w�w��Z�Ay^�o�1΀������q�^�{��G��%��Qt�uzܶ3!�Н���2AI"�B���3jz?����\����2f����k��~L����MÿXiJ�Q��I`�N��!�iԛ��~���K�n��a�
;�u7�*'eG��1(����<<�����D�f\8�A��T�	���O�;?bM�N����M����	$!�z;}p/I9μ���qa�̭�Y����0�0UQ쇡ڈ�xb^�絺�I��m7BIK�0�8zD�yo��t���exL�X�����6kN�-�ɔ˟LZҕ�xy���I��,GV���[���"�.xEt]^Q_
����F]dAr���3��.���c�I�n˽j�C�0hl�[�`#��/�������jX��pδ[u��pE��~Z]�)2r�P�z&��S���TN`�r��u��K$�zɽ��ރδ��	~����h��(Vq�\�4��X4��a%%�x�-����i�A؇�k�Ӭ��ߞ��N�A��P��+�
N��
�UA�Y��r�����"���v�z��5��m=ҙ�Jt֤XM��^ƻ�b��#7�<��T���b졚w�(%Oh��&Ĳ�Kpqx��K��Qrt���"��*��������f8��x,*��	T"qKc�i���;���m+��t*_�r��G.��a�m%�T�*Dn�FŤ�O�(]K���u:``����8&V���C�g��i���[sP�k��%��K�_�9��^��mi�G`�Se�wu\����5Z�ȉB@&�� X�
Gp+���DU7�Aw� W�^��U��B@:
{U��x����������y`(W)�i8M�#iėZ3�h:&>˿N��]�7�'�ql%y�E�'>�?����ˤ��X ��-�vF�4�	S��M^����H
��*".��pk�xˤW�4�fc]��z�?�W?)��T&��t]t�Q�l��<n�@^�c���)�r,ȓ!$�7���iZ�AMw%R8�~ӆ9C1ّxşC���A�Z�x�]�l��j�����&�Ж����Y�����K,S���� ��Ҩ3�lfX�m�S،N}8j�tv�V��*��\���0P������R�_[ |&�:w���4�* H`�*��~}1
S��B�1����Xǅq,H���O�1�N�2U�$I�t��k8��~of�z��y���S��Qbz5������0�	#��b���H�d�&�}���C<n�~�ӗ�~?L�v��:\�	RƜ��7��+m�z�9u�g�&�^ܖ��U�2��e[Q���3g8�Ae��QC�%?I{[����a<jO+9a`�Ȝ�S�D0#cJ5�r��S�' @��t���$���f��愶��f�Q��V����DA�nK��f�@���a��,��p�o����'�s�i�]�r��������H���/��OEa���1�̽�"DD pkoB�47��{���+Җ���2y_Z���X�+��FjD�`�Y#hWRrL��?�xp0�-��u�y�eq����o3N��L��\��Y�57�*Y�c�]Ũh ��i=�A��Dp�q.�e��i���p��v's.ݹE߻�B�8(���%~h0v,�w<�v�?s�.=q�����kլ��,��R��F7�R(>`�(v�sN�<[a��^F�J����s���myq���FO�y�f�����'���7��ox���B�+��ļtB��";Ԇ�DH�� �Ne����W�b!�?�l����; )�K{G�y}�,%�V2�|��u�>unٺ��w��+4����AuU�g���j��~�٘� �,g�0���W5}WK����G��b��oX@�]� � 	IӦj�Gܜ�d��ycfh�V`8� �e%8�'[yF��7�Oz�8��2�)+�=��V�ɭ@j,�� �d6:Ҽ"����~�w$U��0�ԣ���F�in]�f1�GIs�=g·X��i؟"�����#�$���Hw&��b�2��XQN��r�'���"ё;���Hp��<{�#�L{����ClV�����)�	o��\H�(E`�Saj2M��xoR�8]�o�oyJ� ����IG_5D����a+�/z{Z�C��Fl'
�2J�W<�&�@ }�����ǬL��,f����� �������J�Z�u�[yo� �z�1F��:�G[~� A����aUnPt9��p��Ox!�l�x	e/�#D�+)o�cR+5I��M��g��E�*SZ��=���-�K憻�<�F����at�ߩ��+��-T��8����N��G�F9��"��ɜFH�-�==�ԁh�Q��^J��	�g��k�����C��AČZx'>�Ş���=Ē��b�(a814�	����Յ���* �{M���嫁������K^+�	1�&\�S���E�  wgI��_�*���q [��)�0�0�>��&�9������H��u_��K��h���J�lIv�vjс�:�9߶]i��*�
��V���
u�O�����語՝l.�ee�SE��&��l��k��ъ@�����X$����
n�C��.,M�����,a�%x�ۂL��-H\,�2�x�5�e��3�ё�q�B��t`�6�BBn��Br;��I%q���ai�I"5��!:�I<:��5��2���C����{H|�m��^J�o�e.��z]ސ���R��Ò��M���bl|�W��!��U�0���ҵ���^�ښ�
6�8�B`�����?��&Q�w�#��۴w��[�?t�H��j�M��*W��L��$���<�Z�*.\cXeR���B�R��n.���i�����>���q��A13ήyp�����5�R��-.@9IFm��?	�� �#1:3����Y���É�#d7��h����G����#��o�*p�V����u��:'�o���q�urv��F���;ʙ :Wñ�v�h�|4�c�h�׹M���a㽳����o�w��GWD/��:�v��3��P�)����0�,���n����Ɲ]�xS�}���I�}��o�.�Y�UYy��������̯6�ni]�	���{�V�m�YO���\�%8��%&"�v�C�M�҉��{�!k��NlbW�)�q��_P�����ࣼ����ʓ�U�Я���;DR|,�����=M�T)l���rq��ܐ90"%�q9�5��v\_��4C�[�`�x�z1E��)y�#��cd>��f7Lu���@� %*�ߤ~��Ŗ�����O����������"�4t:`�zo�Fnt���z��v�>K=q�$��������&T�l}e�����}�:��O��}r����`f�T�<Od�]k=���ͩ�J~��d�
f�,�l��W�����o�?cP�����M�ٚTq�� މ|&�2�Z�#��k��P���h*��ɀ�n��0G��+�8�ػ��t܈W�� �S'h�Ӧǀ��&�!j�k�i%z���h&@^��쒽����hր�*����>�`W�Ri~����Ŭ�������!J
�{�W���a�H�y����aa)�&��9�B��Rp-D�-�X3�ROR'�K���W"�/�7\*8(�?�>�ja�g���V�%�)�Z�ӫ�	���H��:�i�w�U����:��c��≥�#��د�8\��X���13]���.bQ���~jN%/���[G�hC������ߢ^�����w��Ɍ�&Y�~=8N^�Lvh6��L�[���<��68�����Pv0���W[�,��M FFuڽ�ډS��@~�ܤ�CiA^�kkE;��_	�H�b/V3�-E�y$i���C�B�xވ�r��b U�#kf�x��y�M��ƣ%K�B�Þ�b��5��x佛��l�a�C[�T�WIܰ2���D,�	h�:J<��_�������[������o>>�i�,؊7�"�<U7���%��U=�l(�����~�:�7Q���˸� O<�'�� >e7u?_� �懋Wx"N�Ũ�c�_��g�Х�;� c�=��Bm���oP�ɝ ���+���A���t_墿u�0,�S������z�w[y�-����2����J�!9��)�	{-�������*ؼ��F��&.O�C^��(�OX��w�k�@m�>��������+��a����/șX��]O��S�(�E���h��lugD3_M�)�W%�r7��_���� N�� a\W�xl��ݴ�n�? �<���$(0�AN����1��T1 ���dw��"����TQ&kN��)��s�AR������3��,;B���^ё㚆�����$�"�|�n��U�>��hO�fb�G��ã|Î����K�P�oZf�L�a�����o�#��=T��3���F\'�O��/�y"E�o�[9t�u���Ӟϑm���3�����O�z��]u��[�oTwg\���J�ֵ���{����`��������ɘ	���������θs���H-~ƅ��Z�~!�w3qj΢�(������\Xd豯�:A`��^<\mjSU�&f�>����u�_g���3��aF�8�F������36��,�+oYdԶ6EH�<~k��x�Q��Z��|�!d^�ѓZ�ޕ/�w�<���pLv��y�I-�S50 ��2z�.��V?��&�t��q��6��B;�Y�8�Z��w������}�WL� �� '�F;��K���	6F�2�YiyT��H8�8�2�nė\�B�)˘�s5a�4	^�Kꀭ#�n��G��\�k?�_y~¿�*��\h£��U�O!�� d��E��Wv$V�q��6?�")�$�j:��we �U�����,����?�h�?��pA�1��gP�M����L��,0C��Y�4u?�nb�'e�]4��
��������Z�[@��{�2��p��d���猜f�l0$///�<Y���*p��fZJj[[�������v��֪�^�~ ����S�c���#[ba��0��CdGx��uy�j	yt��W���?�����\s;W��D{����&bC���T���`�-�x�+4���;��T��ڂ<"��.�?L�lA��{Y��MS���:�ԕ6�[�{&	#ii��cYLè~�09�0���.ʛ�3��c�����.�pg����>���
��H/�����l��w*#��9B�_
�3�E���Ӝ�f��,+*�;�ਙle�E��#��2�
hW�op��8�2�e�#C���1�Gk2&:����
��A����՜�D�ು{r ��ۯBC'8�t�a2�6�aǲ<V_�L�y���x��Q͑�k+���ƣ�g?���Ӧ+z؞�^a����+1�ǍU>U�=�3X���!�,5J'�|�_\5��<R��:}�������X�j��>I ��u��������?^��yS �?����;��O�"��T�58 f�@M�&�A��8��t1.`�KY��x�3$���_%�[�%�^�es��ݙ���}$ŭP��z*�|=ƶ�&��-���e�Sa|2�;��MKy��;D�FEQ���Ԧ�b��^���8J#���{ל�uo�,?���7�F�A��+����_>����]!�E;�J&J�����p���4�+�-W���(k�Qd&�4g�r�P���_��	l���U'm�:�!����w�6��+!6+)"�]91B��!a�j�f'�d��E����M��-:a�-K�Z�8���e�`�/|jW2GrN�I��.ay��RWSGN"����.͖���ݖ_� �Db��
3b�5�?PΘ~��{@�K��Khpu���l�c�2�rT�t�x/�g�R�[��k���<��j�D@�#�@����Bק%��XG�z'�����ĕ�� �����<N��S�B��`�=�S-���(5��MR�L)g��/��,�`�2�`5i�?Ux.y��q���Ѝ�Xt�W-����]67�Z�$�m��w��v:���0�Q/�܈����q�u������&�oNzÖ�Q�Ƃ�����47_���'b�e�H���Ʉ|�������JLIÚ�=5"4�{6x�.��HM���+<o�]�cBP�>�}'�5�2��q��\�\u]��E8���A�� �5��Md-/�h  |r&0:}��e�A٫��Y�Y��?�[�����{Y ��W��G`҉彝w��	�a 9"�G{�tȽb�Y
m.�1�V ���IX��.MĊ�- y�+f47%�~
�Q?�&V���MV�и�uH��8�����=RCun��z�=ph=Af�h���Ȏ�e��]?���?�C�M�Bܱ��u_}�� U("w[,�	U�B�ֺ}��'X�	g�Ll� ���y��66�$|V;q�_5-.���ɒ��i3��WG��fR�?p�u���ߢܭ�(��,au��윾e	��Zf>o���Ή����O���G���;}����� ���ֈ)n�����G��|6f�缪_�1�U��L��$��&�0�PK+7���S�߾����Bc�t�z��^�流�9�-\�&�B�@$ �������W�T��M,wP� �)��6w�J|��coz�x3΢i]l#�:0p�W����@ �ɰZP_j�v�H�qJ� I`Ό��m�a���%.5$�LQ�;��%RT����C`@���dK"���<����">W�ڧ�Lp��,u�j�vn8�@�m�`��R�?]C�%������2��i�d68���뽲C��,�̿ډ��	�|^�Hs�{ �wשQH.
��[>�p��#��0F&
o`�9fh`+���D-T�9\�*Fм���Ei�P�o�p�v�w�u�mS��
��3*���ZTK���4�#����h�"=�Y�^�!�H%�u�:����|LV&ul�Nɿ�;�v�j�o�&W�^�l�rа���&*5̫���)Y�=�:�gX�����ީ	#��C�)!��8L�< .3��O�s1�����A��h`+]�qb���#s�~Ç�v��H�^�{�b���i��B�����l�kn�������y>m�����UO�%f�%�<F~<)D8?8d_X�̭Q��)T�ƕA��G`k�o�~�.��v�b̞���3��8=52z��Y�ֻ�o��*�O�� ���;ʻ�+fs�t�V�ٜ2������3c�
�J����O 6>���cp���6�@��h؛"��,#N0����):�+m;pܖU�x}�7�q��uNs@�Kx���<y()=m-�(���>�O1�E�Y���3��NڨKZ�>Xc-��[����R�{�nl_Hc�H��#R�Y�{���Ue�T��5x
-��c�h��va zެ;У�	����	>��׫w�]a.����b{�*ք{��8l\E��9$�!����V��%q��q�������1����t��J�����T�hyCRt|'���?ڿ@�`N�nf~����]�X��*൴�L8'@Bk���f��*�Wx1���%� �X������_��W��}�䫲c+r��?^L��m#�R*�᜹:�]�n;(IfF�CX���9�_�}TU7��.��us׸<K�(H��-��p���ɡ�^�R%�1N�_�ZD�j\}L��LMTy�n
w>bA�j�/f�w�̍��%�$�'5#�)�r�����+�
8]�G�MM���&�J��L)zX𫢩Af-�g��]>�>2�+��Ό
3��N�&q*x�= 8��>Лdr�ٿ���	��3�[��5��vJ�G�X�"��
�B,�oQ�ݪ3�KD^���s��$�?H|�}��*��%p=M��FrK~�U�W�?��p��
��<�=s�HV�$`~Pc�s�M]�%n��RU%��|X� ��k�"�M�i*8v$ ͪ��o��/K�z��2b����!���6�����cY�b��f�c-�%=�bF �F3�fv�S�%t�_�'���,����22,��)�Z.	� �-���"�MJnD��1�{�܂h��Y�V(YdK�ʗ��`����n�/m1�|�{H�����~�&cƶY@�y5�nzx�a @w;"gd;~/�_{�`�O��1)r�C���4"x����3����5	c_�l*f�?�D��~��mCI/b�/ �#:؜�yǦ� E.懈_8i��c�)��#��>� |����񨫜$�옯���լ��Z ά�>���y�\�2	!��t��)� ���J�g��+H_1�x'HX~�k\�bm}�S3��;�j4��%hK�"�59�&>�<�wq>�OZ�9�F�Xd{���흏q�}��HPzm��n�D��ĳ����W��\�?��Q3ֿ��q�kZ�J0ub�6��a��{��OZ��ǂi�Lt�E8��>Ϋj�!��'�������F����������P�f`���j�U&����w"����&�8���֋0�0��z2r�i�G�+�������i�
a[��LO��$�-��8K)������Ns��
�[D�x���o�_�VJC-�W��:�$��$:�Y�A��65�ޒЅl����s�9��Z�v�Yp�h���f�v�&�f���g�����h�H� $:q���V�?��W�TbD^15�9,Ƙf�R��y�Cr)L���;�-c�o!�}��,�>�lc;�S��w6�_����yg+�	�2 ��4�t�\/5<����鍅~�"E)f��Z�������]�����h���p��Ł dpA=)����ZȚ�6?�U����Ш1j�6���ڈ��w�����?����AS��f�^��y�w/�^ѕ�Ls�ɖ�[�?�H,^�fe����i�9QI��߷QM�Br`�J5K��.���~re�C�RR�������ft中²'o�LF{]��9|5��ڑ�����6�<�*����;�����Ti3��+Vr&���3�1�|^	���l�s}��n�~
=<��
brp@��P�d6��m-!P��E(��ouUF���%[�Q�?P�T��&�����tť��n.&]��f9�l@P��w��;���m��X}\�q�ľ�s�P�
�.�^��R��%��,�����Tg;u#̼'ć�E2����J����ˌ�|@��\ϩ�Y�!�Rq����G���tm�Y�-h v�R:��.�?+x�I������4��iT)�dN��7�%�~��r�^ϋ���u��m����
�O_#��FBn��/�!=��BMņ��Q9e�FAٹ��*���#�Puڦ� ���sd2xN+4g�1��T^�w �/����}<E`��ELϤ��QCv^xԌn�a~�Nҹ�>X&����/`su\�1%���=k9i|y���t,y���N"6�;��}����}�ʽ��oyo��tV_����u��W�Ʀ#	��e�j?I�'��V{��(��^%���`nKg��z��)�b�WVLZ1�	h`$����е���;E"qTLA�R)�(G0Z��[9wϽ\]B �<[C,A�������4�4i�b�����.
�%����
��B�������:m-go6)��ӄ :c_��xb�Z�A2>��Ρ�����coK�0�B&P�/J��̗Y�����O}D�k/#��L�)Ws��)���oz؎g����M嶮0c.��Fi�"�����ۯ4uBy���kd�)�ɛ;�$¯���r��^�S��P�uj߆	��m�?�m'"�ko��	�a�*��K�ͧ�Cݩ��Nc����&Q�C�rx&J�gu0�lha$݇p��X�L���hrTȢ�zQ����3�,�BU��������A9�o��Oe�qƲa9�1o�g�ڵTD=�����n6�U�NȤ+�ʚ��y���tWq4�WG�{c�t��8��C��;��@��2"���V�v��*mbZ~N����P���G��0f�#�ĕ#���	~ 
rĮ�v���ϔ�M�����u�'�i�>��B�}�D��SE?�t�{������7���4U�-Q]\ͿI�E� �r�\v��K�C)=j��{K?�i�,��24k��2B��ev�DsE�{!����h�B�6��&mw���� 9�g�|G�M6��hsu���wQ#�%�Z�iv�d��p������$G�G��qS����� 
�ו�c6�˂t\����7s��^�t�����x^�N�t	$Θ����Ȓ{	72j̡��O�HM?��5.�d7q��N�a�r)հ�����o�
jHTgє�3Fwp�"����~��w�a_��/�i�U������{'K��6�X!	"@��'?n��؅/Ӡ6�$�9�c.?O6��Z�Kr�����݂*�O��g���P�$���t����AV�j��Ԧ1�kL�_�f�| )��u1��e��y�/��I��w��ysedӻkǢ�W	�´�>K�iΘ�A��Z��_=`1���GHf'ڌ��)Tv��C:v�$���`���<+��w���������Ǚ��_D)�`�`Ow�d[o[M�e�^��6{	���~�����`�BG#~)#��ʊ��4>����2�'`h�f��:�5�/��h�"��H"�e��HP>�hR�,���ŖnHs��]4cm�@�(y���Pn�i.�c�iL����f-�����X�l����Ǐĉ �8,���h�����5�����q�m|+��0�qz�n���r�ڨ��3�v ����w}*��p�6H!��x��5H�����ճ��_�gڜ@DL	�wb�T�B�-A�w�y��b�����7�U٩�wC�d�;;�Q�d�����J��]�s�*U�D�#�S�����n�gB��&#���K�Q���|�;�Zf�D�C��V����G�k�o�͘�RK0w����ҙf	_1+2���=����}���`Lw��n3r`!�Pw.:p�!���u�]>;���(�>�;�]�i$���mƝ}0e�B�Ȧ�g6�z����n��t%�&�t�׫-3�?��l���y V�W�����h����s%��E�kl�Fu���p�6E^ {�pp�|}���l�k���6�d� =N^�FI���K��_.d���x�G{��C5��>�$��f�Lf%Ɯ{��,��m/E��=�����t�N\��T�i��T�h5K��]u�FV�WЯ��,���K?��C=1�+qB�`�k���/�iqݺ
�B�&���-c��&mi&M� �ps��Vl�>.���!���so� |Mйް�	�E#�4�϶���KZ\'����7�߼��ꍀS��O*��uZ��f��8�{uZ8s�;_e�S���"b$���ɗ���a��m��@�Ip�v [��e�ܺwɟ6c'��'9�BOK�t�,P������,E�����}즇l%��
N�'E��*� J�ßD$e�}s+�m�8:8s�+�]mb�-M�Y�d�YYM��+ق�#wvsya�=�0�8ow�:���8v}/�E9�w��ϱ�`5���_ڇ�U��!	g~V-`�����/���۝�l�:���qc�\R�ujg˵!~���Ab�t���tؕ�ڰ9�ӷ�x�
c���@"���HU�R�ALƏ<m7g]��3 La�e�t˨�.�Hc�$M�Q�����&�qayZf*����shp]�ନ�d��(.-t��񀽕�/@�S!���*�+?�>4�ػ]��Lv����e}D7dA��()*���p�ȱ#��Ư����X�h$��A�O��b�k��e؊ �����$楢s@�"b4��Aɗ�]d�(:�i�Io�]/������W�:���ް�]�\��)!9��=Q�vp��S,�
��wl����;崓*
�"��N�HR��}�q9ͤQ{��;�ܼ�=�&S@��4�Bաؚ^�l;�	��o:�`E�m��'P���l�b��w���S���p���+ 	th|�$��dB�|���^CL,2o��X�/G:rnTϏ�
�9���!��N}0�S][�6Y���1���^T4�7�bj�u�϶F�`·�ͨ��w�%-6�*��p`Q4.�%4��4W��ּ<�/��0U^v��q=0��!i��l�P����Ǿ����{��PO3��d�!���L���w�4�@Nl��?��#��.�R��"����Ճ�d��9��ѹ�����i�7��F�^\��yFN�<�Q;�t����ir譼N��!G����Zn��D)^!���-��Pyj(��A�<�A�k�}���b]av	�xױ���_���_�g�Z༆\^U$�^�p��$�ʌ��Z�g�]�.<�p�T���`|�oI��k��a�M��OVچ0�!��ՄM��rћ��]���G��eźC< ���[��̪8$r�Qm�:���;�ge�8� &}�H��)�'2w��9c`t>�C��98eB`�X����hP��$6�*Xx��dڂV�KUvA����֚hZ7B֠0,9�Y"�Ӽl���F�9f�گ�!Z���k���ʃΛ��6{mҰ@!�S��6�6]!GJR�Ŕ"��p�� 4�n0FJ3���	�dl�^��z�n��W��a�,�*�vT��][^��)��w�\�SC����j��#�R(uD̰�Q��a��l�X�`8i��ohl ��yG�j�w��QD䞵�#���u�cFj��0E[�?m-�j�]���N�� :�ϤA��B�=�,(Y�P�ԭ����E���T��m	ַ�9�	H�+�z���sH^�:g}T��6�)���,j<�����rS��K ����g��=^��G�d)Q��q6ܰ�c<��,OU��~��������ER<h�u:,0ӄ|���J�'����,�roR��}�J�$�݃K��Y�n��T����.Z���g����������jU��M�!�0��UU֌�m¶�"=��*S�ū�>d8�jw���Q7�
r�f�̈́�#g˨�Y-`�62��E�=�;����A�!���;�4!�����vx���܏����-[f�Ӛ����^=�	*�j(?�,�E0pf@じ�zб���#I#�#�D��@�l�߄k�T��.E,���HIPc?D$��D����0,�,�	�V�\Ժ�n)I��߻dڄ[+�Ƣ�����Vpk�MOB0�_K[T�m\.9�B��y�L�{�mru, ������=��l)���?�(���Fl��͟�M5I���q�3���g�q�FHj��ԏ9�1�ӻR�vmf�][�3� l5Ti�0��l1�(s>f���=�5��̃�/�"��S�E���
��������_AV�J��#)ȋ�x��pR�8*�@p���(<��%� ���y}Q�iO��vXk\���ϔq��{��9l�ʾ?����B*��m,����i�"���@���mzLV8v*R�^�Wl�F��	��y�P�h(���&U�ٞ���ǳܗ���������m��]���w�\P)w�޽"p�x�P�s�Q��]s��0&��y|2�*���X�8��};����w!�B��`]q���R��0Y����l�6d#[���~j�8��ׯ8�ԹM�"�YυQ��`�ͪ��'�Rt����x���b0����6����pw�s��6���
H�Z�1nv��� ՏFT��8wUi{�咔�r�� ����2����>r�������L�4z�ly���>qr���o����d@�K�(��<�[7�bW���IG�Ȼ���EQ�jӵ�0ڜ��T�S#^�_�&��NJ�v?�0������G׺�V�x�����8�������`���HLkX����LЎb�����!<��%�*2��nny��e��8��dm{6kX�C^ҝ#�x��5�V	����?Ym�N5C��0="���x�f��A[ӕa }��9}�r�"�k'���|aJ�d�b:������fD��k���Bέ�s{��P�l�z�
��f~����D����{��iq�?�S�߂�hR���f�J�,e@��O�����/�5@���B1�1�U
�ࠝ<�E��p�rKYJf
��*ڤr�ʴ!k�(��u��<��QE�6��K��x��i����\��2Î���q�c�����{	�K�V�9����M���T�4è�H��B��&��z�e
r3T�P�?H	+��s���@�Z�s��za_�81�6����E'h{���Zҫ��q�6���Fo�Jc"U��p�2�љ���,lG���JgT4-�Z��W"�9'1���Q7������`�)�w��]�Z^ ��]C��M�T"rZ��^5��:���3ݡ�A�me�)�Ȅ��d�<��ċ-�@�#�
�2�D<�+'.G�g���*��C� �sy��(22��u�= K�W>���N?��D�J��+Wh�G�V#�q�[������E�`��ki� �����ir��a4�>��Tõ�����8nS��I�_��3���1�6Ǣ��(��P���ڙ��ZI`_Lt�4�I��a\M�>�nFtnSq[>��'��Io�sٛ�H�6���=�x`%D.���<I{rl6�!�b��:a�n��s�@T��m�B�x�U�-�Fa�mv����v|l�P^�~K�5n��ݪ�'�� GDrχ�Ձ$N��s�����I�
qb;.�EX`r���ܞ��=z�X��s��F/a��d���G���v쇁8K��~��W�o���+��OOM�Z������Å'�r	��l���H�nRCT��+J�2�׮�f�׍{Ew�kM��W�fp�8�����Y��9xNF�b���!�'�����r��^0��Ɉ�\)�6u`��
sH�~�fl�р�T��hܰ3��y"凚բ�h���Mo�~5bn<��i��Sh�K�S���l��%�	܆�O�]C~��7�C�eA�k��a��������%���*�30�]��n��F(D�����r��'�[�����,H�L�1X@E�Eh�Z��g!������3�ܱd�ӈ���jz�ʦ�0ۿ� [G����̥W����۩b��s�` f���W��j!�7�ʣ�Q2�e���� ����Z��hv����nd
u��+R(l��U�j��I`m�	��x�zUcNfc�G���pJ� �F��~h���͊])9h��,��dB��g�>4xm5���]$���%�4�*K����jy]][l	!k���&���k-=���Ff����"t�Lh����O�$�^���簢!���y��~P{��<$Dن��'9A�m9���'�+��iwTƟ�0�ge~�Zly��L�_��wL�"�e�ؘa�*[P��%�����%It=�Np��~�z�9�u33���,$+�	<eΌ��S����aBӲ<���OB���bp#���-��J�ϰd��j%�.���i��>� F��>�U�
ش�q����r�>"DY|g'_�i���h�ʔ?%{�;ճ%r�����W���=�0���lջnG��y����Ce��Q�5�|g`�׻עh٘(�!~7����P_���@����78�
�������>�V.Y_�<�Ւ���j�<���`�%$u#����V��zw���v�����Rʝ(�����W��g/!x.����a�i����%=DH��T)�G�1��.�cW���7��.�L�hy����	��>ދ4�)�J��?�\7�7��B�@�v��Ja2�ֻ/χ�lc���@#?6b.EOq��yM�_�
3�y�z������A�����}X��++5i1:q�6++��7��_�ڙr_3����Dec.I�%��d��\���'+)Ѫ���a~���:nF��d�^��Ij��G��F�Hgr%���Ӻ�t��CGr���O�|�*�g���8J�O��?	����@u��N���,�b�K96�J�.�K1%n�8�:��۾V7�����c!Do�<:��ԣTB՛��ԓĬ[��)_�j'����;ۀ
���5|}������9xР��<	<���)d+jܕ{m��O�s�j*-�o���z��,���w�xr���q����E��S�P��O�M�R�#!�7k!���&�Xk�8��!�Y!x틉E��oϐ`��X��'wP�_��(�0��ps�,�F6��IQ��FdDT=x*(��0J*F'\巷.�-�u�[����X�D_�Fc�����k�gM�r�M��5(�	���@R�ԝ:�H�Ɏ��hGw�߸����%\I ���H�z�_�~��y.;�:��S��2�%��=@[��h{����2�j�Ӛxղr���.�q7����?�Ҿ���A7r6#���v��̅3��f�
۳X�Kߵ9�q����$����MPGqb��,6o�cV�V�pC�D���5jU[�
�aBLc�|;�ԛ
�m���Gd��j�x���uՔ?1W{�U�M���'�_f<l#��{S�G�Z��G�t���Z�f�>�dڸ�Cby8l��8�ܽ"ۻ���!x�g��[7�S�R���Q�Tۦ�$�����P�L&�^k�U�ש�,��W�Dq�se�3y�{uo����9T�M�a�ųi�a�F�����NT��{�+)m�E5V��ky��p�	���C(�ip�*�rI�H�tR]���Xl�؏l�t3��K!���T���.�(��yqOy��%�����΢⊓C۲'��tĜN�[���(iD8���8|qI�o��G�p�B�9=���G�'��*.�m�Y��#l�Eޗ�������(�ꑿ~�\B��sy�L�����ր����ظ�M��\��R�y�3���ŚV�t�k3}!����iq����ag3Y�Tu�+t\w� L.��cgC ��`�$;�lA�j����Ԩ0}
5�rDQo��Y��rP�Ng�f�?2��AE�>�I�������y_�q�w�_i��(����NH�*t�6S�i|������&�����m��h��'L�#r�{v��Sڙ�&�L�G�MCL��G�����ȒV��U3tZB�e#Y�Yx[���VG��0�2���6���F<ѥ�yi]}�<���܍ב/ԥ��K���]v��,���^j��"����%�9-UgD�?���ƭ���`��p��+��������P���ތ��wB%�B��Q�6��dtХ@�[�{�/���J�e��I\�_͜?>�l�C�<�	C��o �D~��{���oZ�k[�am���r�{w�P�k0�L�g�O��������ѿ$����Zp pD���8�'�z�����O����m��^n�߷raW�J~B�M�Q��7N�9�C56$����Wd��!M�ɘ�R��?�xEF=�
���{L=M�t^}&v��z���};��ꬵ��3^Ѽ�I��əjۉMf��ë��!�B0�u�\�ŕiz����/�5�H��VSS�&��m]ȵ�����V��D��e�Rr��]B�TV|�� n~�1K��2{	�T㬱���q d��o(�Eq�e������?IE��zL��ό��w�^1g�DW<i�bI�f8��F[�R�<?���_W7E�/�ZjK��)b#��R��nŁ]Z��	������;w�"�f�6k'�z��hӺ��SgԔ���d|VطO�8�޶Vi�u/L�|)u{�6�:`�hxq���vh��˵S�<w��1 @ �{�y�K�h~>�;��榭�_�dpON�l���K�z������H(+�fI� w�]��!�AgO�}�..�%p?:z]��S���R1�9�6Ӈ�$1���3�,ƽ�&pV=�#����i�އ��DDх���	�zI������NQ����:5��$ںO"d��sWZ�q ���`XW����D$�^臤𥷶/������1$a����{��<�)�t�����k̸ٴ����@��W֟A��B�
l�ޯ��+�*lP4C�!�	."fށ�O�0��Y�5Q ��UJ�h~���]K�ī:���<�.�KD��^f�-���T� ܖ�&(3����	d�5�F��aY�9��Ղ������ŧ��U9h�kQ�M�������^#7��h!o4W�I9	�ŰKF����s{����
�7� ��,���$��x�fr!��m�?��YzR9��N�H �G^�o7ֳFuyh��)�k���q�P�����;���_>��������QQ�O�e%�O��Հ�8	�^=���,�֋@B��Aw�]��h��ًf��Z�
�bn�m�S��/�?j=>^-��]]7?���%����KeC�Zh���z0O�N��h�GR3�'�ǟ�1*M�$'G_�Y?�K����r��3��K�HL���x!�Ԇ�ef�/9����I)Wnӟ)�G=��N��a��85�qּmV��3+�E�K6FDǡ�{ŉ��bi�q�Ӆ.�o�32�����ҫ@�_ZI��q�NI��� :�_L�E1qN���_$S46�&W[�;����L�$�;���h�T�-�(���K�u$�#p����n�@����v!qA�=��C�6���֙=���nG[UX�1�bR�Sh�b���2VO�o���0$�`���AA=Y^�V#�T6���-�i��*�dM�����vQ�gw������p�
����V�:���+ a|W�X�0�d8��rN�An����o�3(�xx_��j�g��v�9q�+�� 4�,�h���{���f����������.'i�M����d7�����xv̤�E��a���m�Z?̀:}����4��J� %3��IgN��D�d;i���{��Uz/q�w�N֮6Y�OIۛ'�kv����t�wN��4�Wl����]p>�⤷�5;�&�c���@�E~���@u��'`�'x����c�ۧT_cvj.�f�Y�o��Ť�»���(���E��&��?L<q��5�b6z�ۿ��xڂ����XJ-	FI��C_�dC{B5��힑5"\9?��G|����\��~`+wџ@ฤ�$� ���I��FNX������X.<3�2+�/,�`ژ�V�B����3�����'����3�E�*'�e14P�|vK�w��tU7q'fH|���=����˙�օ(M�Bo��Ԣ�F~S�n���h,`�����㛱��-]��������� 	�<����s8����L�?�CS��:���S�u�iB��V���=�X�� |/��S�����cK�BlB�����v��S��OtCx��r�b�͟%��x�Ks����՚=�_&�ά�]{c�^�Z�f���v���T�Ϫ�說Fl.��/�p|��/�?m{�/��!���F<��*I��c�O�o/���u�9����҆��/�+���_��:�&��
$�rju�3��)6.�V�-�(�"��ֆ	_|"�`��X�j�:�Ǫ����*��Fћ~�i���QS�g��`{$|�t�@�����$;�P>e�T���{��H�y�.ЮS�9G����˅uc��s�Mq{9�]��ʍ/���$쫒Հ{I�9�@Ĭ�x�Ɓ��[���' ���qx�!+a�ߌ �6N�@�Z>�2�0r�v�A��೿���,����/#4��wY"�SoY����
O�%-�Y�؟��z�&����Ľ��.@"HX	k�!Ŵ�h��?�^�G1.Tkn@Ԕ|+��=�3_�]��/پA�����]�?<�]S_�d���bj�2:ruEm;q�ͥ�%^�
���{$?�Q��Pr�-����ԧ;*Yּt$����
���O�t\%%zKp�\��o��Ӭ*��E�q��:�t��.h��hY�rN��P5ԕվv�޴GN�7�w[yy<�N�>�e��BDe^����k�_W�uƪ��zT� ��&IeU�:Hc������Ni%���4���쐺�[�@��ļ30)��"sV�EgPp_�s��	`Ǯ���Â`��9�u��dr"L����c-�K8v��NVb���?�5���H�2s���n�:���|B��ܝ!ЋЖFr�0�G��vT�p�'ؚ���l���ս�6ag�#㨺BRk_|4��|1V��/k�s$��f�S}�h�k���-�ĒGN|g'���f�z� m����^\<�߅U�dǑ����x�a���wo�h\WӜ4q���[8�7D�;AbK,��?UCמ2�ϙ p�֊�~-��`�H�u�>t��,�4�L:�[���z�gQ�V�f]oW1��n�����
E���a*Fu����-3��!����|�ﶽ��j���XJ�7�f�S����.�{e@p�1��/�WA����)n��>�\���v�=�hws��N�������m,�2Y&m�B�> zJ��g�����6������3Jw�6��pd�2 Ċ%�2�GP��*�ކA�i��Ƅ���f�spG�'ŋa/#>x#`W�����Ă��Ŀ���q�h�'�L�/�:&ڇ˭	�J+7��;��.Y�+��$L��5���d(��Ag�K3˱իw{x�5
�=|#�7)з�r���S}Z~73m֔�.���F۳�|(�1��2	}3�K����m����6Seq�ogB<vz���V��ҍ,/�bM*�����]��_f.Q� oU	4D^�
8��G��G�c>W�ŏ&�s�^�jqŁ�& �-�&�3���;zi�$^.&��� �y֡cr�|υZ����3�T19������&�7!!�s�ͻ|7��`��Q�����<.x�>-��x�0��ܮ5��yz��[]TI�n�U�E��G+��#B�o�^� .p1��+�c����OMP'l\A�a�ͶB�M
��e
1�f~�SC�� "�R';�h�C)����)�^�m�}��wX*�d@��f+��g��>����g�Vw������qj{�����z�fh�3��iJ�g������`�� 
�P���yj�jX���4�����~"Pc1?[.U4�^�㴖oÚc����sｰ�	��]����o��Ѯ�p�^���^UZ|�J
���1z�6�QqbT����>�/S��8;��C@g�,j,8�������6!E~�w�{���N~ *���#���g���L��?�JM8T��*�ƙ�wm;{�U
�U�Fo������$h<�f�u���V	Tx���T�e��}No��O��gjۉ~�F��Z#� �����48Yf�b��֒��f�x�w�^�)�����k�.��pl�/�1�lg�G�&�z�"�=��+!oG2�'-��Q��_Uf�Ϭ�U���J:Q���_���.�S��fާ���z��z�J�3Y�@3+A�yЖ��:�B�3.f�Fg��>H�sq�j��a�⬝'��'@:E��q�YHl-ך����N�<E�&n�E�f-�A�u#|&>4*�pZ�*�e_���FW�Ē/VG-�vm���XE'��&h�µ/�����4B������o%%�!Ί��~sv�����]�(o�6�tD�\Ƅ�o���8&��2���ѐ�0��m�텿)8�x���C����r�X�y��B����:B����0�Қ��U�|z�S�^w�\�FDr�������:���wv���H���-�4*����'i�j�Y� �����Y�Gt�i����U���n���j��ݳ�gR��\��!����Jـ|���Vʣ�-����8�$�銆�!�le�ҧ�5�u�#O9y%9K�v0ˬ͖������@L̅��B^���}�9@���hz!�kn/�)��i�J�=����S)��wxS�0w��T�~��d"A�K��!�	%��M���ޘ�B��"��OD[��]���{����&fwiT��5Ϲ�S�0�v�"f[�������
e��D/+����"Y���9'�q�dw�6b����=�բQ0\C�-\8��F���{X����-�U�yJ`�� ��A$W/��]ؤ��{��)�x=�mQ���H�2�-��UX�2���ψ}{��??|���n�`�����K4x:� �ku�ε�3?�)Y6�r/�b���#倫j�����i����_��
=���T;��]�H�|{�E������<w�wl�6X�jƎ#��q?M$*F���>Tw��!�RȱY�>��3�q/��[�w
N�WbY�'�m����*���c��2.П,��K�C�Č�2�z%��WL�T��m@%�V.�v��T�T�n7um���0}��V$� �Jr��CM�M�KO��w.�TS���<���(`w�>�֪�XO0�T��C"fg1r�|����U^Č	o��g�Ъ�.�;ÒZ�З� niG8��i?ݕ�'܈�����i.O��ul��&�`����\�N!�[�^����*�Ĝ]"�v%�X^X���>����?�t]�%-�P�)3%�G7�GS��$��� �:8f���j�"�*�����0TCO5�C�~�����"�y����m��^Qg���p�
c&�, L�P����*A�`D����+%�J��M�Ğ�֧�k� ���P�c\�x�^0q��E#Q |oN�O��� -MJC�yPd����� Y��j*"�0����t<Mj���%sB!��k�4sx��F�9s�䗬�c�#�O��Q� �"	�-\�M�����;�ܢ]l,oaů���x�����nGUl?��t���* �q�K���&Vz�ݗqڹA�a��c��laR��?Zb��U i��b�����杂����$�f�_�-�;�p�u9�_φ�x�2��K�b���4����������v���T2�ޖO0�ͯ2㜋�DU�'/0�k�^��m�'x�Ԛm�C!#��y�
��Z
� ����4N�R-�e�_�ֵ�lr����)����<��P�������O�.Y�'�4��[�TdsD��4ճ�����rDJ��}����%�M~��s��D�Th�{�L�C��U�k� w�bY��@�_�=�0�G�z�'�ϼ<�h"mT+W�_�����)�����}ytRs$MMǽ�8Is�r�Έ(��OM�T-S�M���s(}���c ~m�£鬂��ǭ�yۻk.���Q5�A�\o���MLI}-��s�@�w5���-���7^jќ��\��SK�pز�-�`���������gZg�Z�
-�\I4M�V����� ���>ז	��ވ6�m�
�>�r���e��DǙ������G��u�/ϋX�ɱ�"�|�������q��>,@�&uFo�E/3�b�Y��p-Ss�X�L[5�����?�ክ�ç��$	����[hG7; �h���'�۪e��L���^��bʿ���a*qN#R",J���ft'��/�p*n�n�?U�Kz��O�#�y��gW`p����,1'Q�t}a����B6b��?�6"�1RK��_!��U�0�E� 
�=Y���}Kq��A�{s)����Bٲ�6�ͮ���PGN>-q0�D���)YEp��(�u6N �[���`A�&8��o Ko��r���P��=.y�jk���k2��S�(�\<��s�ʄ��jm�k�E՗�=�+u��_���
�1����҂�f������W�h9����U�">{^C8�Ht�:1��lvE���t�:���5��:�_�~��%��/�Vh`�y!��l�ŃLQ�O%�U5 �����#��w����X�V㯈�frN}��U�h�b��׀�~��/���(��M���z� �1a5x�4�̠o졕?�xv�M�:W����^��2ք�S�;h{ދ��t����@�Q��;;|�����62��Q������H�	�L�au(�A�ȫ+�h�,*yk��^):'��|�a�u��q�;��1���"�9-���R9`L�.m�y�G9^~��v�����E��f�rs�9D��j��j�!Z��BUdK�YI��`�F*u�aR_�X�9�eѠ H��s�a>��p�i��4���e�,һ�/ 	҂ȍs��ѣQ<��LE�iQֻu`ۤ��A�)Ҫ)8XI�0�/�A^�)Xq)��&PX�wl�W�crN���@�@;�,�ߔc��vL�_`�_#�(nl4cA[�+_%�p1�������������?>m�U��A�-��;@&���v3P�5�:r~�%���
���Ю�{��9U;��g�s��2w|^fG�X�t[?޿1�dq�MsM��^�}k���<4p^�lG߅NgD܎������\�p'8�zqJ�5��7��Y����Q֨�3�9x	�B�ar�S�pM����ȳ&1��4X��g�J�]�����Gh���Сz���A=���Ai����D�u@ "Izy�N%�3���`?����bo�t٠�c[�%�8�Sa"�^G�a�Y�Nn�`��ZM��IO_4��Mծmw�]QC�%ѐ�y�z=8��a���%�ucH�Q�������g��?#0b[E�%�G��k�ygn%
-l��ל)Hŗ-S���*�ƣ�n���ۼ� Q$��ۖ�a��
�H�^��k��;gr����~�7�zϊ�~�EM �v�c�G��`~��/�E�g�w�xjY�[<~�e�Ό��9�(����͢p�K���f�!��F?Mli���������<��(��f��-�Y���u�q6�M�Q�w���i���6�L�/�u�\��^PWM�zu��[�/�a�� ��1"�!s�/<Yj�ם����VE}�Ud`P�̑�ݍ���˲�%�:����ׇ��Ǩ�|k�B[��cAF�L��]��Н}[V�+^f��Ev��{+���������L�U	kŚ�͹���Rv�O���xX;v�FQo6��C]|M��Í�K�yhh��Oә0B_����>������{��zC��V�[�哻�6~ m��2��MG��$�2k�&]�֙�]F�Z�z��w�ԧ���lu$�'��r�R�ؿYUUi�|F�;�"q[��Yk���s|�/�]�=mD��S�-����!��4�^0n�N��Uk3�YR�(=�q�c�HB~�&P%�Rv���~ZacG )+�f��� ��#Vz����`D�h�����%,s5)����z&K&��ي�_;�r�����Yr�Rٸ�妦��Q��F��E2$q�_I��aw�I�8^h)�!Q��W�H��X�n>Oea��G����:{� 8Ä3�x9kC\c�b>|j�ma0��1g��@HX+B,ʱ?L��2d;���O1o�+�����?����R�C��+޸�pO����$����=Qt�y�ƣ$F���$���x)���7Dsf�l���SN�L�[�ϼ����r�/P�*��}$wH������A��P�8.�{n�iO��99�g���e/��fb:��jﾀt�&��U<(�wM�<q0s� C��kC�ೖ���%$�K��<xI�V�:��la~r"]�}Q��J�r^^ ���w��l]0����:NߩRN�PǭE�A*���В��Î�gG`T����ΚhDO9J�W�yD��t�r� �$"�$�ZU���Nk7k;�L��"YԽI��4�!M�����P?��N��cZsۖ ��ӟ����Z�������mX�Y�4,R�S�H����ݨD���Ne��Zyj�#��Rp��w�C��O�G�����_��Î��������h��Wl���CJN�ˀ���:���]BM"��� F�No��������5b2� ��9�*�^�+|�h���-�G�������,$�f�/���^�@M.�i��sb?�H�'_c�9��'��rƩ+EV��oP���L���1��(�Q�*h������3%I�U�%p��,R8��)�
u��6��M�ъ�T	�;�d�1��l�ڢ�2#�]���߷�7�5��0�?���o�' ���آ�`D+�?Ʀ�Ԓ��3b��`,|�%;]��9䴋�j����=�	l�<=����cO1�,�p�E���1� �C�u�m��u�p��{ ��.n������eӀd�US��'�`n��;3\NoL�	��Q:BD�?��&��c�|�a%��i��[���˓�Bvk�	1��/�/�S`�����2�7E��9�(�i=ݹ<���g�]C	��m O�i:�&{}���[��2��B 8�c����Ey���:�L��_U�QذU ���˻�*��n�u��`�3lsߣ�;������>}�99K��=C�J����B��!:���J�ؤZ��m���'�����=0�^9a���V:�����n�n~N����e�3�V@��߃I���^?ȪKe=(��Z�c?�%�����"����eхľ��_��(������dn�]��F�~���x0�/�s�Cëj<[�23�Ӓ�\������8p����|��tY�|KiDАu�z�cr�� �������=B����;[�����1bd
.����-Sf�i�oZ�1ZקVd�^�'��/.v���!�2�L�����x0������ct� �
a�}&N's�7��-��؟�*�Ǭ�t��N���<�*�/J��NZ[
�o�&##�������}���y���l����%�dr��A1���|�u&吏9�Tт���|�@����@b������[`R�º�5��+K�h���{�]]�&RT��	T�63=EՈw�N@x��@MS��O��p��鍺ul��)��Jԥ����WMT�;�O���kt��[���#�/*�F�z6�;�m�D����̞�}@)��ef��;*�`��v�������8����S���r>�����J�J�A��p��[��S;CX޶�g���!������W+�Va��:.a���-�U�A�D��U�:��-b5]�D�g�D�'$��\|�1��������y��/���y�'�-�y�"���{�I)��P�	�2W��Af�z�ʵ���}��L�,c8�ߴ�$@��D��@K�q[>���,��-�'�m�����/�b��:E�f8L	7�ݤ����w�Y3��r @���r_w
�qy�v>��?��k����p�ٜ�I�=u���S{DGܩ���2Ь&5C|�@�ܕ����x������c�"��cOd�1D<[@n��x�J��9I�f�����Dm�bv1q�T/��~�Z���{�[�a)?�������,"N�t�2$W��Lc�ډ�/58w��.�س��������ƣ[2��'IC�� ����y�,�W� zz����1ï�E���,�VQC�ڷ���9�މ���됍��\�p;�R��%��K<�t�`4�@�ȌLjF��h�f�|5���)o�������6� ��˃X��	�A�/��+~��d\��!�f)1�E�Z�4ZU�ksn@h���rh�������b�������`��[��O���z��T0�kt��!#�p�!
LUI;ChdV���-�S槭�cf� ��Ȍ}G!!���v a�������w��q��B�}��e��G������VwI���%܈�X���j�E�*��I$P��`�&�|1�6��0��brT2��.I��<�R�}nE�4Q��B�d���Ё�]&.S(��2�W�͵N��v�	�6�y8!ʾ{F*;�T��x���#\��!+�^��2�]�"Txo*���R-���u����-����?���*��3��.��Fv�M���35��a��܌�4'Zt����4i�2\7qE��h�]�?i�|�0�D-�n�*�^�k���� �^U��v-�K�w��`��w�J延5� W`�|5��b�c�U��F�c��_-Y�t�t�>�繦�����1
6�51�Y�r+ߟ�x�`ZS�5_�����	)���L�@O��E��[]����F�������,M'E�K�g��h�=53�]o�;3&l�����2l�r���N��!w�i�Vbk7��w�Gǫ 2Wʲ�&&=2��Q"Q��W��윓�d�-���3W1��e�7�CͰ^�j���p|TL`�_]�h�\�aT��s�X�������Y�wǰK
0aw�C��GMO�ׇ�8i%,6R�f�� ���ے��,�x�7s-߅�b�,�2�`ϙ&B�u淚n��<���!�F:�S�1y�:!���*��5�|I�WJ|�}"z�����.�,��t���[�꺴�������D��i�����Ӱ'(����9���F�q��⁋`|�s�T~�`iO��!��_����Η��u��(��"��wA���{u�p��vu;�'g���6�"5�&�6���w�t����"��_�����.܄�����X�6w�,Z�na�g6��@���>K��gD���#0��,}��-H���s�.��2���Q�ԏ� ��q��:������D''�a��!|E���<�\�@tf����S~�1�L��/&+jvqN�Q{N����j�R�B�E݃7�X���,Onݘ�<��'!&�s��;��ܭ�SSe2;�����e��:W"��O��ݑM�E�WR�>]�6p�`���!e�Y�����g�N#���d��"�e[pﻪ�zw��d�A����4�F�F�Y�?)�;�+2��2��N��ߚ�e	���՟���ӿ��d����Nc�L�Q<�`��C�����$�y����?�:u!Sw&X�b�\+1�����Ȯ����,��qJcy-�-P�Ox5S݄���+u�+f��:�/ǈ�,^�*�)�ZM=���}�B-8����#���a=V�	Lgg��7HY���8��Y
��c�ܽl��˛bk$4�5]�X���%¥��լ�ё���%f��:~�L��5�W�A��%�6�E0����"�m�@ ����� ]s�����w��ʋ��]80bQ��ʪ�<����XE�h/�� �p�7 qF�̎A�'>d6VRWdɀ\o���`�T���6���=j_�ݑ~����;R�K�rT���I��	�6���}O���o�`�-y�[r>$�6F����ĠȬS�Y|�?�ʂ�I��1�F}��R�,C���H�	������E��^�[�Q<.��x��D_�&�8_��Ml�xT�v�1�-�d4��&�~T#���]����L�z���C�% ���@��FH]��'ɑ0G%����Q�ꎯ�)��l�N��}3���:O�.�Sk�a��K����2r	��%��E��3�xf�Ȼ�rݿ)�k1Qz��j�"e���{U;ބ����i��$N�T���Ō��$�l��� 8J ����S���*_�E�K_G/���ь��l� ��G�;#��Z�v��I4q)Rw�[­,���N�~�>{�܂�ksq+(�+#�&�x/88n�6���8ʽt������k�b�Q�
�+���XQ�y
�Zy��F�k�G0�D��曃��W9���c27z�9i�n)�����	c�Xt$
^&�Q";��WcL���;*�Hd[�Jo��?�AQ��Ztt�D�� �U	�]~>Y�M����a��E;���`3�=��5A�vQ����/����%V�Pe�Q�n̸�dk_���WM�BN�! �R��C�	�al׷���PiZ ��5���ɧF���G=Í��}�]�֒{�l�$�5�"K�uѰ���R]���aG�d�gcu�C5�c�pQ&����L,�Qhj�LR���L��]���%����W�ļ|�"��(_��ab�k����d=t/͑��M���t��Y?5oѢ��8�a�y���}��w��������c7�1��i	3�j�u����^�2n���Q���_�j�7~��Z˕�>^��7��z�[N>�̍X ��:��h$�&�3f��X.)���D��l<"��@�(�ڕE��C�^�jW�����*���9��$�my&�ు��wN|L�Y�!d)Ip�m�E[p�ik���/���� ���"��	��pUo��n�����@s�zǰ��-J�	C�/��:�g��:��X59�k/'f�B*0���A+��&��������d����<���%���ԅ˕Ǚj��3�9~�Z��V�;2mf�nҬ�S��ǚ�`�����Ҁ�E�V�eE̲�m��[Vg£VnN�u�E)�=wS7��9vS#FX'U-C�Qf*r3�/�F�G,�h��q�1:
�g�Ǌx���#ӆB��m��W����E���F�勴l�	vV�{n�����%���em��v��k�c	��D���jF�������1�0�0�XeO��x�G�Iz�*\�?��O��<H����#+�6�w�̓=v����Z��x�J��}�Q����q�{3[VD�%)���P�͖!�q%E	*br���}W�v�c#Yb1�-Wv�f8g�W&P�N<vF��G2�'�mNs�}�/�g+��W����?�y�������y���̩����,cC��f�6��y�������M�'�#D��&r�I4#f����Q�v�w��g\�*2s�juU y�X�y���b�$J��.էtc��ڔ�$�����9���LL	�R�y��sמ����2l�<'�q�y�&�{�E+P:φ:�ؠm;�#�U�#��E``x��sX1�v&�Z["Oc9���3�O*�bB
!R]ҍl=���)�+j���S�w���\���LE�7�+��B�M��+�7�����Q��?��CK��OA�?o���śA���@�ā����a�S��I'%#7�-T{{��`�6b=U!tC@'1)�mn*?י�#ߺc8���@\��!m�]��<ͧ|�Š��Z���u����i����p$��$j*�"sĄ�J�Ԍ�K�әE��`:ݡ~(UF��Kg%�
�-ǃS��ZQ�SX{��c1����p���z����D���N>�?c���4wӕc���;��fit���_������hl2X�*��U��G��]��&=�S�k����&�ݝ�Iø��U�ĉ�t���Տ#9��� ߄�4���~A���Y �@T���S~&�|����6��A�70kG�	�!s�x�YvaxMD���c4�	��0Y��\�f�	~7�CiDl,��5}q_�7��D�4��A�Bc5��O���s:sǂ�	Im���]�qp�:�U+�(ܙ�4��ҌOQ���1[81�#��PkY��΍���Io�R��&f��I���۶+�|[mԴ���w��?Id��.�F�V�n.�R�`o������0���0)�	E2 �d���Z���칪Ѱ5@h)S�M����u׶*�C��q�e�������7��mP&w��~��^�T���+s������)b55�]�����~�I�b+��0�!gx.@��1F���3A�{/h��6��c���ޤ�T�K�M��g7�eQh't�̚&߂�N$��;���DX��� H��}�ѢR���qF�� �E�
g���֞����3w�T��ޛ��bx~�Ԃ�,ڙ�����0-D�������t�u`�U~s[>]��Y/��d�V��:��$zȧ�����[�,V��5ǻ	�1�]�vo|}��cmR�T�}��N�PFL� \�N��~K-�|&�Fw1y�h,0�Q���F����*�夙�������u�q�I��c�ROm�n���o��I
�	�f��+";���k��Ȉq~|�'a��T
\�$־���'?4o��%n�Ri�iݔI��I����F��T��:;2�ҟ��w����+=�>�>�O.�� i)
���]1j:���s�*�2°�F܇�ԞY�`���#�H��-���n���O(���W�cT��:�GL6#�1o�}�%|�-��z�4e��[��L/�.^�6>�@�sY��@%�|^?#zLL}�qů�T��݊��U:-&gr�3��i������yG�y����Wr�#�?��&�:��P��Z[W�ua��X����Ep����J���cljܒ�B(�ヌ�Q��-�� Y�1�����KN�=�y�B��ҫo^��i�sx�@���\0wSQB6p��3�=���1)c�O;�&�WO��z{_BUQ/}m�����b�S#�?���=��������s��+���W���fT[H>��yބ���� ?lg;����}�W��S�����N����:�.�w�K�a�9Õ,c���8�7�� <��H��gn�J>*�	e���4��V"1��ܨs؃M�a-bd�<�>�����d�a�����r׮$�R�B�*�MԲ����bC�|n�}�:���F����!H�ރ�=���Q)W���4�rD8.�����]s�T��z�1��.6Š��!�H��$�.r�%�>���ݪPt/)h��}A����'��>sL��VQ��O�g�IZl,�"u��d��>k z��}-+5z����1q��$��+��X��!<*�_�\�QҎX�_�^�ъ��]�6�z��;���6)��G9��$�D�P�_��������
�nG=�r�j2�Z�)$o6�Iƨ��tU18�n�P��S�2.�lu����^�<�����;-y� �b��S���9�o��0h�Ft1vS� w�Go���j��d��	C_��R�W���v�䙢8cA���NH����Q(c��D�����Η���./���b�p� �Q��� O�SPG���v
��U������:k,;����`]P��Y�3^?J�(��=Yݚ�P����T��-�Ѹm�q:IH�-c_�� �u�%�����9��2��O��Ǫp-/�����P"7t9w�I���,��5r�'��lɖ)�آ+����R2q�	��/o|lZ��5��S��qՏ<h�h�ڤ��ar��&��a�/�"g��"����V��<Am�{�j����`c�o%4��%��֚�L�79jjŘ�]��]�� �<�)4�M�HuЉ�"��B��e�b%f0խ�y�3���o�Ӈ���5Z�3����������؞���	�h��KW!T�Y�w6IdV-�ߘ�Eű���������ޱ��4�!��Ws�O7Z�Y�	w�{1`��2��|G�X�'���pE�CN�!Z�j�B�s��y���#�6'ҡ���&=��9Iw���FGp�%��5�f`��=5Y�Rԏ�s�g�J��ߛ f�dΒރ�w�[�0'�=�L��3.�t�&U��xa�KĆ��?Z<Y��� ���Ə�`�Jͨĸ�sJ�I�VV�~N���G�#s��}�~[� ?C1�J��̼���a�M�2q�n������\5T�W��H�oj����Z
%�#��tX�mU��-?!���6���e��6�=��1^�@I��4mn?|��/��N�H( ii����!ܲ�����-n�v2T�}U� n��T����(
b�Y ����L2���.�Ro��>���#��?�Y/ �}ޑ��.��N�!�!
$�"j��l�(����RI�QMq��r�P2$���[�Z(k�q@6��m��4��<��<	<����p�<�`����[���%��&����=��i�Ue���
�e��L�/Phޠ�8�,)��_Eܟ���{��h���{!u�픧]��w]A�M���� {�tG�Fw�t�$v�oZ����yR���׭/{����"�ڶ�q��3��P�Ǣx�L��^�v�22j����1#�	�fBv�22�����6�u��$�Gl���U�����^�!�@?�ͥT��d�\z��;�,�D�)���zeg��QO�=�e���[�B@���f��_ޤf�>,�S�7�<Ҋ�?���W�-�R �3'̯�q��fگ	C+U9�̭-����m߇�d�����h ���M�] ��Bv�6.����4��C�J��Q��RpZ���RU3P�c	�Ǣg��h)B*e�Yj�"`�r�+�����P�_IYIT�a�'U��D���C�o$�x����c�}�)wr�_�H�z�,�p�fxHPK�Iy�y�K ���M���u�!�&'��8��R����
[�)�r�^^'&�&$�����<u���[o������ҕڅ���$1�v�#�ӣ!���(����r��e����U��w�t�*����Q����V��N�O����Ȧ�쎅�OS�i�T� 5��K&g�A$���(h�)�e��k_��axG�.sܮ8E����Q�|Pf9Xg53��zA%�?k5�&���ܿ�bC_^u��ir󮥝X;�8YK�}R�m�2vxM�$����d���n�V?9djER��<9C��\fw�ݸ��o�� �΋�7L$Z��M��Đf�2��6�?ϸ��7xp��X�eI�=�[�f�T��\ :�k��3E��U��q�A�!֣OG���'R9!���1�B?�c(F�8�������+2���� �Sa�4^e�������4nmV�u4j��8 ܫR�ޓ1)	�Q�l"4�*���sY�(K�8�҄Q�b���46����#py����s�;�mc<��D"X�Rjh N�*=\@	�1#5ǖ��?�	K�~�!����C�sQ�8ɶ�q�c�Jt��lp�/�G��� ����r�l�es!��/��������N${2�5ګ���W���S�^��<�V�� �����+$��ȨN)��"��z�#�Pn����h��t5L7�b"�@����%!6k�q����k�A�xjz�(T�!V���V�����-���)���\�J&���w� JNb6�r�����J;U�kq.f�<��ʔ�3��}t�P��0"||n>SG����K_�D\�x���Mw���ke�SVB�π�y���S�u���(�w�A&��Ї��?�����D���A��f���	ٶ�jH�({m1:C���63��7��ڞ�/ж�`:�vo��e�n��(g��<7A�'�R�ZX���Icx[�=�Hғf��b���]���KHn����BV��'��(��Il
�=�p�pq�N!a��*�q���d�y�>GQ�N~f��-�g�K��NV�e�u�/�TK��á}�Q�՞9�t�;�*���w�?Q}�������Ѥ�292zjx�,W�,TDAc��=�V��z�pd|��V,:��	����m덕HH�q���]x�=u�l��ڇǉM�HX�eVa����G��!������9Cy��s��'@IM��P��h�g���9�pH��U��m�1R��1�8a�R��0��,^j�B`(�Hh1�.;��ȳm���tU�"n���V���65�����'0�^u��41{��j�?�k�pTL��z]�*��Q4U��W�V�й9�w�r�y���O���y:s�Fy��8>����-Cܗ��^@���|!�{���C���q��L�=��bwW�9�i!�b,w�B	�a<���m|��xH#��s�M��'�_�� ��5z^���-�����$���G&�C|���kʌFS��m�~T����B�'m�tx�I�㼫�(��}��T:��Kc�bU�ԒSh�B;�^RcF�P�
֥�b�Ĩ�M�S_|*{�3�����5?�a�7�e��8&��:�Jx����ɍ>Q'��sf��Ƭ��X�T�� �1��07�Y�� 
+=]�ñ�I�[V���יU�����1Ww�w���� 8 ��9g������K��p|����xib�*'�u�����0[�^+�k(Y��|�!D��]TmBz���s����:�P}[CԾ�T��ߎ�j�"�/�1ZP;�/����?Qm�e�/:
�:�sǶF>�vTW��/pS��a_P��j+(r�r��G�ׯ����1^h��������G	e�s�k��K?��ķ�)��8A� ����|�������p��M��|\��e3]|��Vm��qN�0!�ga|��sb|M�WN�Fl{K�1��,�;��Re9b���nt�����"��r��+i|П(������p؋ːaJi�;I���	��l��FŃ�1�Nn��?�˹������M���c�*=��<�p�T��& 2-���s�g>?X�d�]تE]Y��<�]o���>i��c�w��f�'������
?�]�����c����y���EvF<�EVQ$�ZN
I��Jѿ�������NU���;������D��=� B�H��	�v�mO'��~�h���)]�')��"�7��	�ڭ�:ߛ:%�s.���r�h��J�\D���� ���&�����g�H�-W��%��s<݅C���	���v�,��{ ^v����ȣ���9�=T5L���Yi�X;�QP�5;��Q��9RU�5q�4�e��@ɠ2��@~�6���c:��K1��ȥX�O.�N�<���/� m������ـ�Iv�� p���E�d��l�:�h/��^�.��i8i���H����6�Ki���6�����R��-6Pr~�e������6P��m���NH6�м_6���ᐾ�j�K墿�c̳��%\�D����tB�J�G'9)�	��R��Y��~���yeF�k��y6Xd��%�a�ҙ�kWA�OK�9�'Ն0�d~��G�,�F_����ka��RL��G�P0Y�I�~ݩ�K�;��Β0(�qj��N������ �H�1�i�J$���׭��*��g�Ń{��K���i���~�� ['K�R���2/� Lk�1J��w�G~��^7� �� ��Z+���9#oN��������^:��w賯�2���[�"�M�9MK~�aP%���g������o���2_y��c�%�8+�vb�R͓/'�����@�3)�T̀.��V�p?��)U+k�:D�/�$
'�7����(&-r�4�]�A����|x[T�9�dAecp��T-�J�9l�����^ �2G��J5��K.���4��l]�D����'��ծ�B�{ p�{��k����Ʋֹ�_��4<�X��|
'��|���f�3Pn�}N��k����FЊx��_n9 	�1�r�h��<�6�R�S+�z;h57�2�RF\��=<�l!��M��ɡ�B��~���7N�@/ɴ���N���ѩ3k�/���U�&RNz�������������3%>P����흉Ά�� �{d55����gr��o)�nuC���Vhp����Q!z`���j֨�����'��-�0C'���M��-�OH�2Bt���H�3�l	g�}o���h��%��Y��L�k7s��o��LS�,s?D�o�iK�5��;&|�j�}�l��!�֐(�V��航�5��N&�IҰ<�8��Z��|I��'*nŊV�G��⟗-�k߹��ʳ�����PVX�� \�/u��}� ڟ�f^	��P�v�����n�����0��r��e��:��s�&�.�>�m��HN��_c�/'��>�t���	]������F$�)��ދ�Qe�����6}h��A",8�^�!�Z�qOp>.�7=��)B�����+����$���Ǧ�zp�KA7u�z(^��h� ׍�O�4[UL��x-��f��������/e���	Ԑ�$aj��H���!t��<B����+��s�R����~1w7*ڧ����;�W�W���w���e����wT��[S���y|�驹g��Y;��Ǣ��|�J�j�PSi���A�<����L�9�Z��	��Y�Ä�z��CW,B;L3�3V�j�0�q(i�'bv63��`�l�)H:����5�iǑD:F���]�)�ܝ�]e7�<��gi�S�W����0�z�;�ܵ ��r����\��ա� !<!չ�;�O�4��%�b/R7ޠ�]��tz�Oi|7��9.C�� �2E�Lf`�(��ޗ��|����U|k1�����$��\�y��/��*��Z������A/x���n䇣1�n�H��"���A����5��y͐F��!m?�r��Iγ96QW�1����1������XG0kR�L��/S�>������;q�im�s��Έ@??�
0 ;�S��@i6b�^A�G�e���*���w�u��0�@zb�Pp ��mK�����*���6�ۆr>�
�<�ӔSҀ^�Qd1�	���EWa�l���C1��r���d��K�Gn9�ϤW��{�c���×){�ܼQ5V�B�|�ā��$&�D���L��v��f��/��:y$�����x������?k\��M,�F	5O|f��(���Ԗ!T��1nT@��nHfv>D�I���P�$��g��x�1��r�*��ܣ�T,Ē\T�6��X�"g�zU5��S���m��)D����!v�W�q7���h��H ��kcr���� ޸I�Tΐ���ȭ+���K��έ�.H�H�qK��}K���Z��*yC`�l*�ƣ�(�1�	QR��e�����hk��ilá�p���n/�{�Tڵg7�m�
j�N(���Ѱ`�<���$�}���٫'�ƻo(�p�I���^��RKE, k��2�D��WCX�0�:t�F� CAW�ۤ@���N_��3 	�#9������XΉ�\~`�Z0qd_���lg!V]<ǫ�G�oB��=PL�>9|u	���}j���U?J�6]�Y���G�U����Kc�QUW��� ,��+���$u���X�qI~��&CX�zAa�Y��۴�k	d�Kء�V̂��i����p$�$XOm�l��(!�R���{c%�b�u��-�6?���gXF]�N�u�q������{Ń��x�Q�2Q�,
i�т��{p��oE˖M�O����u�/W?��u�<c�Y�g!�u�9o��o@�3�Aw2E�N��}�{"�O���גf�������fY0]Z�Sq�Ck�؟~�-@�._!��g��q����m�Hp�h�ٗRb��|�]Q��%0G�����%�w��Q;��H�+BSJ�Y��<a�z����tW�r�V�����~��Ɯ�^�^9�e��
��$�1�8䧦��̇���ivy��$�{\&e�����Z�F"��6��&#O��#RRdHeY���w7@'��Ij��h\~�45b�v��>f9���!8����O��t��#�;��_JUhfg��lՆ;�D�N��H}
��V�fm��������/Џ(�z���R�	8��"�T�ur����_�|)9��uPC�>�;r��ky��Y�8m�TB�u0��Ef��4;��T9�xy��Tb6�v��F���~$iY7�qs��?9�_2J������y�>h�:�|I���nώ��~R�r�*�, ~�BL2�KmI�PD,~s�R3��P2�+�Q�]6ct�Q�q�;�p��L�}�CS��G,�����#p;Z�)&�-��$0hr�ݭBD�?�����!$�����&��.w��岝�\!���kn&��ߎK�P��ܸ>g0�����N�4&A��m�Zr�i�I�~$0x|�s	�>��]{�x��B�Ұ�R�qVf/d_�׋�z��%�/�XEh���������e�G��]謺][&���!|��	���	�5HUk�q7�s��p�6�o�@���}����<��-�D���'w�O�$ݞ�Nc�%�Dy$�RU�|����7�DCZ2~W͝~�n0���ߎ�͎�x���Z��sF<Da7`O"Iġb~;��I����eˁ���R����L�|�ve�h @)��j?�1�o(K硡��Qs%�/4��c��L��������>�n�c'
����E��p�ltR#�4�wz�
�}�9Q���?�ե1�����h��q�$����
��r���L!�x2mv�h��i_|��ެ��5K;�!m��U��C�����9�>��R��z�R�0����l�hI���7�&/��_N�߯hv��`��������"����1��4�xZ�v�[L��}N��/4��1��O2�W�㔛�� ڣ3�yx�W��k{d� 2��17�ʀ*pf�bZ�Q:w�N3f$��R�Y�;_A�6�=�z}�� ��^fK�Æ��������܃d���}$�Ne)(cj�Pv�,9�%�R������:��%�^ט��x����l�b9M��;��E+p��A������$�E�be>ID�c��L��3�-;�ո�P+R����ic�Μ�Ǜz��9s��Ѯ�jPIB(M���6���ٱȣ�r��9��^��pŝ��a��f�B.1ԓ�����du1,i�8��5�-.������i�;:^�S_�H��9n_a���Q��H��R������>
aK����r����ӝ[!7*�uxKh��I0K��$�_,�gJ�ʣ0fe�=��S{��r?q�9�V<��A\��^��T���J�E�@[�񮷫Z`LH�R� s�:�X����&)���/՗&�A�� �N�,�b������X�=��M�͡���e6��t:T���,(<+N|3rr�Nv��"�g��\q���m�J���m��1ܒI&��](&V�!R��n��s�(4� N�:�)	��\��I��'F�����s�K�~��zq�uV76}�>��p�E{�O�)d6tswo����}�1�!0�g�Q��|6�a	dH*���Cʏ8�b�>G��oS�%Qf8J�v�X�x?�����1F⧏	�>o~��i=�/�z��pE^(38���c"������G�lrd̳�JSkY9�Zw�~iX'�^z1���xֱy���J�ఘ�_�ݎ#��#M+���[D:S�*��S�x�|�%��:����|�����´{t��σ�7������4������uډ~����D�%��m�s!��
�8���z:%9a��� cW9֚���;�u�f�N��J Ź��_S��D~ ��j�11ز��6�>�"eg��v|�7+�С@d�g6j��0�c���Li��q�_��4��r����8d�T}\x$m�P��O'\��L^������[5](Ҹ���\��,(�Iɨ |*��o���k�� �������*�I=�Fs5��#����FU4��e�L ��(Ik�Dt��@1����
� ľ;�����5�i��7��Ņ���I����(���!�	rua��C�m����?��,i� M9�j1��[I�fi��WCj�|��<����뽚:~
��|��I�O�>
�+��%mGb��;���6��KM'�'�@�j?���S�>�����X��A������BI�JO�9/S}�����X�b?X�[zfT�P����Y]<&"B��,��kR����A�w���	ؗ9������ru�F��x��0k�� sFV�2��<f�DҗЁ.�T&��8Ԝ@n	�Z���������zT�%�1�N�,Vf1<�ב'�r}l��0��i`0lU�B��ց��a�UBm2P(f��������A���t� �!f^/�_hR��R� MB��&���4��$&�s.���S!M�T���Ŷ��F�5���_h|1�����^�1
��m �D9����<�%5��o���ub�̛I�:*�4c�;�_�5����kS:�ޭ-�"�Нl?�T!8R���.���2w�5Dy��+z&��;/m�UH�BU��6��w��JQlZב�"�M���˗^{LDՙ2/jM�	��'�diQ
8�R���E��c	�Ae��Hh��p iYTY�o�#��:����8�ӑ&�AG���!��9~aӶ�,˧�����F�Z�}�UH�88y�MRR���Z���!������Λ�0�FT9M��w)�����~Bvi�,���$		������Y������O������PE��0,�w�5� �0�:D�n\Z_i�Tx�����p����w�h���ȱ�=õe㎶o��y/��5t1R�lD����(�cb'	8�9�Ap�;L�uP
>��u{l���
�U��tB�����j�Vz�bJW�lJ�����M��]���Փ�*�ey���(�F�1���D�S0@Z<PGrI���	"�Ω�s��%N�l�ѯ��u�2>��c�T�c�r��6��:�"ϏJ@���eׂ>:t�3J�U�{q>�G��� �lA�%��q�qĹ�}��~p�v��{f
�d�O�FJ�;�RlF��il�>����� 	�^���p4����ZW�)<�?aOU9�ȹ�?��A-X�X]
+<� �X��>ൠp���_�.�q&���>�4J�B?�b���K��&�>p�Ԑ�N����r��[I��������HU������(ZJ�$"=S�麢͓��L����x����k����Ifو �Dd��Z�}=��Q�	݀�[�/����5���տ*�Lɀ\N�<����>�O���~��P�&�J�����$'ǋ٦D${n�b-���SU���Hf>+H��+7��C������������gWbJ��$����c�<;�l˳�.|0�4�����|�1�e�N+�4�j���`xO����`���d7<��;�WKoҤ�$0�4�h]=�_�^��%����k8^�"(�q
��3�}GO�e��b��u����W���Պ`�iN�'A�geI84S�=�L�{[�Xm��Ɓ��pNW���̯�7�-��]"���jvd1���+mpP���h����]�).����X��fڂ]�����ßlQM�`4`����x������k��HH�4]�]���tSVA��?}wH�l}���ca��Z91gYV��=�}([Q�*:��|��E}d�;F��U@ʕ�Rlk�ؔ��p�����D�QD��절���Hď[Yёf��>OOV�[�*��S�oe8R�7햸/����}Q�����bb�	.5#�g�u��0�yh�y�{�L̸P�t�M<1s�(p�_:�k�����><_���A����D�D��X3M@ѩ�5��u�6�ؔ���L��򢄥BR�*�93,s�Ԅab~iD��x���u��ËI��L�e�WQ9�R���N#��T�{!{�3~i�b�Կ;/�12gG{]��Z��F쫿{�˟�Y�S""��e�x�4�9lh�lw���Z�I� �����
,Vè��q+Ծ ��G.����4�;J����s��_��w�N{b[Dw�\}	n6;	�%뺮��(%��m�t���N0�[@C����7����������B^����U�����T�_���<���_��UVe�;
>\8It�U�*��MJ_�S�Š��*H�2��˾E�&��D}hcőHr�m��@�-���/�J�w���Ӌ�wq�OJ&���MLW#�J��#h"�h�(RsoB[7,���{i� �6(.���ƪ������"��zEC���Y���@�M(�,SՄ�#ޠ��Q�X1Ъ�ͬ�� �t��d��� ���x]E�C%�?�,�2崠�V��[E~%�L��5�%�ѣ��'�n��y_@8|2�Ն�a�ץ��P�]�7���2�ᾆ��"����G5G�AvlOK�`
�hY�z#(<�Q�昵F�xԱ�+N�)�uK�P���j�5�G�&���.�荨]�U����!�Q��M�����~}O6£$�X��wa�z��xʛ	U��_�qr]W9Ƶ���\��6��(
7�t�����]���$U�Z'Y�0z�J�h]�CQ�fr4�:(rN���.c@��<:!�]�����@9䂷�mZ�-��cz@5��[=��,B<ڑ NK���(xB��~ߊ��J��3���Q����O���|m٤�ߞ㤀���6~���]AW4�h�bB���C"d9	6�m	����r�?w��^Aؔ��
H�r���  MO��0��g���{����� d�'6�w>q=��&�h.�p=T�"��g�w9�@�"��{�?$�H@�fE�xw��*�O_t�������w���`g}X>�1�G6�d�SF�|��X�n�y"N��+!~Ò�_��LS�S�`H�GQ��=�k� /w������n�bb@ت��V���`sy_��U�bR;/:b2>7D����B�E0A ��"�e����8nW��T��O�d�ȜO$lXFm�5(0���0 ��p{�e8G��}h0�����7	��=,�Yο(���}g���	 2�����E�uJXMx�K�fa"E��Q��/ͪ�Z5�������ϖ�R#������wG��LQ5���_�%�i�Tb�F�����z#C��3G"��5��CX��I���2{������D��z��?%D:���tFvV��/-4�dʐ��۹�#�n˾1������.T���i{A!���6�LC������O;YW�,�t���R��@)�M��h����;���wk6���9�[(n�x�_�����w|��Gx�>���Sa��7����̫���D��~���yq,����#E��U}�K�=�\�o������)��+Y��`փ�Îz�<b5#+��R�{�>�~>���o��rn�jG%����L�f"�r����Ae.!�Ն��Dmy�u��f6c��x�;�u�*3ɟ}�.0�An]�[�p����騮ȕ~?j|ݭ�Z����;�v}m�yQ mV��M�4k��;?:j�2-�uҾD�zo:�~��^��Pk�����or5����w̒�0�����!��P$B��[v'㷟�^uO�szں��׾vW_�5��G\���-��G��G��Xi�>rq:Z8#�Ѩ�x�>�Xp���X��d��q=����~X�l'����٣�w��BL>�gQ;c����!,#�-���즁�*V�\W�c��M&�HD�pQF#�����.���E^h�Þc�� H��xmFҙNޖ�q��"��i2 ,��.��� �$)��M���tV��T�w���$���a�{����.|����4���?{������ba����S�$�>�=��+��N�
F#7�]zn���4�����>��Iģ�<�Ҝ^����%�E���E.2먏�X��Q��M�P�!��~��k���������,�<�
*���B�ӱ6@��Ҡ Ԉ�sWT�q��	[4��U!n"������Q�E���N+r��3mc�;Z�Z�#�U�
�n���V,X��\�JD4��"Bu�,�M[�	I=M����sZ����~u���1de�\6}7�g!3 ��!QT�'E��J� �^#�mQ�v5�S.��f�<C�V��\u�h3��!�hv;ㅬ��K�4����2�g�C%۽I_�S���փ�|;����/ ̺�p�xh����Y�?����a�DI�%����}�Z~��칰Q��#�x�q�����\����j���猩mt���-�_�թy������G�@�k�m&��0U���Y���p㈋�='�I\��Q��sm$1�=QC?��R.��v`E�`�vtHA�J%�$�9?���w>�í'g��o�$#��=���M�~7�C��$�7��b�~�����Z�lsO��v��y�_ )h�f�2�C�����鳢������X��+f��[^�d�<���um�4��k�qS_�8�xb`���<V�"ټ#�o¡a>=b6�y���v����-�5�� ����1�^�[�t�$0�qE/Lh�����(w����@���y���{UQ���Ž-�vh=�`���e�����a��:�d|k�.���4�j �L��,pӕG��/���I�� mS�`T�"uJ�'�?0�j��"-.���g?`	vIRD�2qS`J����V�����;��w"��?���¿zd������Ɛ�Ev���ZMے�;'~A�k�O}�{S r�o[G�0nLQ�Ht�uD�2�g���R��oD}��&Y�8��� ��=�̩A�h�|QAI�](����M`!,��	���������΅}��m�B��p�|�Ov+�\o�^��
�n�@AiA��c�ą|��| r���[^����?EHP4��C}=DR��=f#��CDOS�]O�G��@�/�%�pv�1Y����~�k/UX}��Ȓ7A�'}�
[+݉��A���6p��`�3�R��4OL3���y�E-I]nGw���&*w�w���b++��#D^��������g��	�ϥ9���2�Ou���`�jG� �Ԯd?���F/%�� �=�.g��:����إ�����=3I�y�E�)���2��PX�6S|�r��|�}� َ�40�K�;��~F?V��$�0��8��Y1͟ǿ�Dv�X�`g��H�H�!��S�X��0��?�"igQ��x>`�?ݦ>.ceW�sE,�X�x<��A���c�b�s�y�U[7fv}gD��fZ�iL�ה���K���g{"��Gx�V�(����<����La�$=s֫�&�dֿ�.I<��帾u���.���ǯ�'6��0MA����X+[�"	w�;�I�K3�x���t� �4kD
�7݃��^�xfʴ��r����9��η!W(�}�S*�k#��������f��D`����tg��=�k������YB;0��������ۇa��	��+/Iq~A��%���X���r�m/�ٍ=.-cc�M�H����0��jO�_gի�Q JJyV�>�����Eu%1+M�o�VL>0k���O�X=�y#d�A>Z�/x����^��3O�&�b��W���I9iu��>�\@X�*�gy�7g{�(�L�U��+�~@ 'g&�?(5���[��X]�qW�Y޳�G롹���U�� )ܳy�ksK��<��_c��|�3bz�ɩ��T�����q��C��� ��)�& �37L���ᐚ����IųG��5�P��2d��?��eGE0������gU�`������Rt;�)�1�]������^�۬J�w�^�Rϰ���>�^���#�`cQ���𺢭�1SKǻ�־q�dZu��*�_3��!���	x�!��+�[/�bH�;{��¤���y⁭Oc�L>�#�K��q��B�>��j���pO�Lur�zʿ�d]��Ҍ�{�d�F݁�u�8mB�3o���o�cQn��*�P�pOYA��v#���+;Uج���@k�/��cR�R�>%��uE���[1*[^/ɣ�P�t��<����c�'�L�݉��x�e�:�;]������H���)Q���uO7�]�PbVϠVs#.m�Zf'�Ybc�!.�*32�P@�c�y
S;q1j������sJ��J�*6נ1Yw^�u�nR�����E�4F���w҉�N�
rߊ\ ɠ��=�L�{8�]����'> c<7Ɍz�l�T̑ul怗���mvkN�
���#���3TKY�����`��0�iN5����{`�J�h���۱�:���l^���x(H><�Fo}0�0���ͶB{��H�9�mV@�H
+B��/�A]ϟ��q�%��ڋO	N��$��4E$����GLW��_bh1E�l����u�NR�|9��׃�)$s��5E`
[_��[�<W�I�P�}�Fx�y*����A̙��z�dx��#7�����9�0&˵B0�hi�R�
$c&N��9���L�̪��G0|���llcu���u�`��l}z����M�PkU��C��9m�,Ͼ��^�&�:��c��)
3&w	��^����V,���GO�VO�t}�ɣ�J��qɶ�?x׋s7-~Q`��Y�� P����oɆ��=D����[�Rf	G0�`p�SZ;]�R��x$�o�k�{V�ꮍ{���Oq��*ɀY�Ș��6�Whdw&<�k0k멺���8��i�	w�R����|��	��������[V��B�Z�$# ������@��ai�yb�׭�m{|�&�G�5�Lr�l�� ���2V�^5��w�'�$�g%cw�ˉ34�í���*�%x�1���2�`�wȈ{��j�[C���m�`�{�YBQ&%�C0c��Kڙ��Ɣ�qgn7$=2a�\h/�� �����v2���v��C:hU����5�N���������`8��א�C�+'���(�ҹf�oC��9}Bj7\�;�џ��y!1�W���&��}5?⯖�����Ǟ���	pUo4�kH�&P�J�l��| Xv���$�iK�?�]��+1ԓ�\g�#Ju�ׁ�t����+6#��+&�S���٫v���/kd͎Q��O�%��
��db_f� ������� ��-��d;���&w����w����
��y.ޔ�����,�Թ���W��2,��Z��I��\] ̓� r���:�/�a&�o��pb@�_ �~��XVn1���bV���ȑ|iϱ�[�0�S\>�����f$��o��o4 ? '�RÑv���A�O�{]�N� ����>
#�1;�N�G{���^q�_��ԙݷ��y�fgk��lL!1MՎ��P��zn��l��5�*r���OFF-��I�4n�,e{j�Ot#>��1��@,�%g�G��Xs԰��0&���"
ų��t��`ϊ�9����)DoǑۡ�+G}P����[�;�Dv(�+����5���&300��B`��x[{�o��L��ʟ[b�A16��uLT�>7�<��(�o�a���CcMy۟�_379���j�+�*��l ��e7*ه�a�՘���TH-$g���N�&�-}n-�8�!��͜�n�	XuF��Q�gD��K��/Y[�Izؓ}�+�9��KFw@!(6]I�V$� �{[�ˏ6Y�|w��k8��NE��r7�a��-�ۖ����q2F%&�����G\�8�ڀ�y\�
��@�KՑȗ�,�a�8�V�P�8\Ay��fх+�=j��Fc�v.X��4�Q��eω�ɬ��b`����x��E�i��21��_�Q�Yl}�)�1:��?��֎�m�P���/�;e�T���S���"V��%�'�����D�+x�(t�SD�n��uF,�	#�S��l ;J�?�
nSϲfx�q�j3�Kf�lo��&/�@�� $����i4S�#$�d��{�K>T�#�0�RK�K>��5�)A�LH�$$� lg/!SՑ��4d�Ot��i�}+�M����P'Glm������N�Ӟ�ᙯr-!!���Ӑ����\���qun,L�#��P�p娶�봎+���g�(�:����:в�aւ�-���{R�QAr��'Qz*�+U�ջ0[G�'f����akR���@�2H̑h�zD�NZi�N.���*X���VȘf�ݜ���ǜ~�qˡ-��Ww3�YR4ѐ)U_ 䃎.7�ǂ���Ԅt8��3�� i}�����s7��z:�OB�.��m��Mcak��`#�L�8�(�3�A�����9n�J^���E.A�&�&��;�we$� [�x�Q����/V�T9�G��H����Mg�W���l�G h��ܻC�]pjf�L�^br���4�.7p�$��H���ʍ�₮dem���8bV-b'��N�FY�m���(@��
Ԥ���n���E~�v$䄳̫O#ԧl G�;���㫡���O��x����2��-բ��!قN�IO�Od&^���Sl�+$-y>�4�%N������'��Y�T�$���[O
GL��3�fh�%{шa��#���#պ��$�j�bWFq��ҿ�^�f�Ǉ~$�P�&�-� �.e���L�q�a�NUlj���=�$�}6�e\����DX�Dqω�0�2���` ���W]A�˸}�������fH.����nO�h�&x�0���E�:n�MV����`E�ޥ��������;�|-�O�Y?n���Y��"���g;P$���b�ދ��"%b1�T{U�M���B}�̓�4ln� �$`��>s����
/��GMU�9Z��Kf��t����b�s̓n��/\� �Ǯ���\�ӌ��+��)����7��%�������_����@R�DG��/U�P�D��zSn�4�(�b�5���p{��ty�-�鹉�6��(j뇷�\E�[U��}	&c	n��ˢ��,��c�ս�h'�2����R��a���ud��9��s�Cm����� ��Ѹ
(����ܤ�#���a���<�3�'K��-��}����D!������?J�l}�*h��sUR"���]��Y��]~����T3bktws�2��U��$��d-"'7N%I��S���h`p�e�Ei�_�K~/R�-��ov*E���z�m*�=c<�B@Rq���;0���:�rd߄}�?��"*�Qme����9� e�#1�az�K������~F.JP��X�H�̵��&��TR���'��V��V�1���g����d���n��٨�y�k�ل�&�f��&r�����&�;g�*���vp�w	�3���9%o�ݎ�t�o�����N�]��;.�_�+��K��,N����/���;{��B��&���]�D���}^�#�y�A�2sx,�s����І���Vs��+P��!Ʌf;��a��k3Q�"0m�h�e`���7� �ϕO`:�}?�6I��յ�����D4����Ⱥ�1l����&���:���M��::�f'�W�
{�(��'�+/Ūn�ZK�V,�,Xe5��}%�J�i6�$��ƘǑK��W�ǌ�ǵJB90خ�jq/�у����{L١SĹ7 �Z�LLG|C[ڤ
�-k���/5S<�jo�Za�Yf͛n��*R��GU�#2J����R�}�d�_+��������q�co}������p��K�v��^D���;~n2���4�`1��,�K���֬_gԜ���`�c��L.L�U�R��G>ךFq)	ݳ�9�ø�xo6�L(� )l�؍&8�P�\��A�\p���XgqA:JZ�ᐆR��u59�3J��
���sT �� �H��"P5����Jc;��������#������y9�j�ɣ;��%s��WPΙ>��U�ȭ��'߯����q�� ��d��[ Z���D\�_��U��;��#�c��n.�h��ޕy������jm�Ϩ��V6s�$��Dɍ9�a��І�t��΀�U�r@��e��ߥS�g�U/�H�]3���հ�Ir��;�"pB��b��`�\����n0�x�[��aw�����5*m|����[�]���U �\�iY���-��*�#���c����6��G`ᣮ�!%�8����fBsJ��I*w�=�<D�8��A'KJ0�e[[��Be&	��ֺ꺹��sgaG�+|C��_	�ޯ*C�ȹh��l �y!�������p�{F�ɯ��]�y�'����c�2�������j�Ս��F�3����Z��IY~Q����N��L�,z��� �s��j�E�>������p�Z___�4�!�����/(G��?(FP�mw�h�iM�.��W0�`W�Sn�Ϫ��Aάa�qõ��)��p� p�+1	$g����k޿\s�0�i8`��$�00�����{�bmّrX}��nW̘����B�r픫�����=����jE`�&YM�%]�H �"B�3����j>i�#_l�;qcD	1���#/hԽ�p�AB�t\0ύ`&7�����{@���fu�
:�M6��
�`�`����N�)>��5vo� $8��Vp\~T2¬�W�*���d���z�:���JP�59��.a>1���f� n�Mcҝw�D�w"q�K�\&�-sU|%bi�qS\��hD�"��0�[�� X�赕H�[s�'oޞ]mF�8Iysb�v�Nru�b����}^��v��zh�q�2���("�eU ��+Aɋ��Q�)Qe������βVu���1�h��዁��V�u]�SU��Y��$\��:��`�q߲�r�༧ˌ&(��ῈZ���u`�]N�P(WJ�`��r5�]�]��l!�0���c|�쮂�"40�� :%C�y�'��a�w@|�~2X&ߍ�~UM˻A!�@���,���5����5�&���lXp�- hN貑�z,�PT��]1�Byf4����-�c�N�ȧB�����,B� YU4���X�x��ʩ)���a��#�8��=�/~���g�P�K�#z;c-ۦ�+�0�i��u���q�9<>���.��yy�����d[=qhĹ�˻�����@�\{��`4ԝ��}���P-�ۑ6��ֹ�$N�ݑ@�j�r�ʤe�� 7���f�=]iG ~!Ҙ&��U�@y�o^R�#~��?B͖��d�u	
��۷[>��2�2����9�N�+��~�Ֆ[���"۩�YN ��4���s3�2���-\3�竕� ��O�F�<N ���������e�;Kn�y0�e��սF�6��8�z��%C3�&������qAdC��C�W���j�?�I�}��T�ȁ"vsB������S�e�Rz���KXP�l;�GZ��|��o�M4�9\�{�΁�U��5t����.�j�q�tYJ {����pKU{�&�y�A �s�e�בE�� 
�U��a��8b���)m4ϼ셕nq
�_���A�(���>��G૳�9��u���n���t��-�[�����1Y#5.�}G�Y$��"J��T��.Gx�D�����<d����?c̥��-M���,��M�WR��;(ޣU�S��,.��W���rr�w Ғ��ͧ@�TЏ�<r�@W
|�9�Ai^�B���;�Q1l��S�T�ȋ'�?/�T?T�%��h�o�P�t6�R�����7{�VhvC_gӅ!E���Rw[��o���$���x;��-d�KFS��͛�PXp�P��4�'��c�C7ʶ�Kv*X���,H� L��{���dk��{ҩ��JW, �fpOP		CB]�P� MTj�B<��Ǽ�!wM�>���r���	�g���Jݢ�y�Ϳk%�5�����tx׶���We��� ��Z�ʃŹ���a�zH���M�E9&p7����w���!~�<��F��p>t����6��5r
�0����ʊP�����~[�R���N��sKj�2Ԇ���na:��?y&��k�5}�RLeПŤn`q4Qe0L�)UY�Ūs"ՔZ����� .�����Kh�]�kО�eD]y&�����	�h�a��J0� B�W+˄}�&`���1v_�ffUHux1S! &�e	{Td������!����F}�Uoiж�c�y�=��&W��&�&�O���Ԃ��: �!W�NI�&f��N\��������=��Zy����ggp!e��9��h��D?��0u8�s�5��z2�2���׎?��>�S+����&�Y$o>�m8����)D��XƏ�\�/@��w��(ۂh�����?��`���Ý,�o
 ��x��QA�TJ��&��L�^T� ��g��]�LzHx�_ C�8�SQ��+`���P��0����S`l�r ��v�Q[@�(�B2k�Os��+�S+d���p6�;D�3@��gһ�"�d�#�B|�3F��.5���vb|����K�I䏌�ha�7Q�+�"aI:B�	�W8�ڞJ�B�SaA#~Q�H �`���Kq�\�^F\�L?d�!Z�X[7��
��Ƽ���g�w�[xɎz�&yC#Q��4�V�G���-�|i��!nCU"M}��sp��I�����T�T�
����&Ȩu����hT�w@%
y��f�?"δ<��� w;` v?�n���1n�={�\����Y�V�<Gd�b\��G'�5R諓e3^b1|�EH�Ω��l-���ǱQP��:��=q=,@z��k�y��L��ݛʬM�k����z�_z0h�����jhV@*&q�F��y�2�IY��ϑ����#j�JQ>s������_�<y�/�g�� ׶Ѭ�:�����bM4F�ڝu����%x����x��#��o���	��gxef�h���ZC!�SG��Δc�FN��B���nч�G�ؗ],e����ݏ<�m4���n�?j��������:�����\�e�1��f���+q}?GP�P�D�bK*�g�옱oOw|�hZ0.�Rd����f���q���������,���vǈ���A�������T��a��~lf_����,M ID�Vks~~N0 0\N�V�c�k��)�B0p�_�)�Z*I��Z� o,��kŌ��63 ����$���]y?�۬T��Uj~���]kQ�+`�LQ��['g���Y�W��E#�C!�T�0�K �.M�.�N��Laѓ*^��W~ao
��1]�j��6����k>�8=�35�O�ى������Bȑ�r?疶4���g�Rc���E��uu����E��GE��ZHWN����MA]�H�#��E�h��z�W��n/�����5�nw��'˼����'d�٣�b��p~� Y/�bb�������yø�p�&���~����/����m��a�3"X9����S.�����eۑ��'���H�M��`4?�~{��I��K�c�[�����X,d�V.vP�HK�_���"^�n]Ʈ��	�d���#�Ƃ{ɶ΃��6N��t�@�x4����,U��8tAyE��:�c�X!�,��n`��R3z D{AX�Z'.�V��
��X��×�	�+�yET�8�
D���8�c���$R형3&�}ܦ$X��}S̽���_#��q�JfM��U3e��Yx=�v*Y��m d��}���7�w��|���%�{V�ż���-mL��AG�����#B�\u���k}�Z)/1)cfKc7�l�/ʫk@����5_)6|ם��ұbu����3`W�3��|�Q7*o��s9Nگ�H\w���L����/�%�=?�0�J\�7�a�@_��'�ɉ}��u�Er�8,	�$���!�޼w.�5�7���6�_
&�@��=��N�t8��dcL�ui�T��O�[e0�9o���V*h�8�͜">`�t�������� CL�8��:���>8/տZ�ug��\��@c��G���)��s�Il�c_j�MSgF���<�MB0�+F����V+�չ��.�F,�*o��68pWi�1Ry��Ӛ��щ�I9|kjè��l�л�4+�����S5/�16�Q\��U�4��.��~�
�u�qy��|ﵫÍ
J<���4@*�G
x�v �/���h��Y��K����J*�z��Pk��Ct�V����d��	oۓ͢�Dh�Q��WTu��_�R 9
��)�9�4��&�Z׺�%w��s�
^JH�VZ^�i�����B�M�o��i��r�˲&��ϼ�9"���f�7B�������;�D���ltOr�m��:����/���S_U�(�>�>k
7�x�e�I�7
�.�]e3��%� �Y�W�QO~�^����G.����:=qoI��Z��wN���c�9��dveȪ�IK�@&�����yQ�N	���$��s�X��&��B̵�k8�<Ŷ�Q�W\�:8�$w�F����R��'�Om�x���fTc����h��<���k�U=�U�����iL��|FI��g<�{35��l@�����
�i�.��	��q�^���k'E�^4��{�ym�~��+3u�����	����I���#̼� qJL ��3*�=)���`1$�w����A�"����Jnhlx��gف~w��66�X~zNVH��#h�ƾ�~�#H�c�H�$
�[�k��EZD�'�ޓl�����v�[�"��-d��--�����"_�>_���B�{3�n=8c�p���!G�@%�R��%�!�V�r`q�R��l��R��EVʥ��q��da��aܩ�!zӵ=j�#�J�D���ysQ��ݾ��M`�k�w�&�C$@w�Cw�+���e�n���@N���P��P��dw��(P[�^S������b_h1g�8lc�Z6���.p��31=�ü�~���bi[����e�����纯��"T;Ǯg���;�@_7�ƥ*�����f2ϳ��VeLY������5��c��g2o���#:ժ|��$�Ă���p���y���?b1�Ј��%�C;�)��5m���F��i���C��y��Y5�J���aC>DC��=��0���OJX�j���o,��s��o���z�&ْ?|٠h��j�H���M2��<i\�I���g�<���v���ւE��xu$r�����yٺgt����mO3^�?Wuli�1�Y���=�`t<z���͗�)�V�8�j�`�x��6b>F�n��~+�����g�����"~Ԣ��������hL֥�A�]IN���.��λ,���k~k�o���4�ކ�4�3j��*=���E/�?5WM�����?�/��v>
�xk,^�{�p�)������nv����9�G�M���ߝ�����*�0��3#*NM
h�l�{:�h�6;�U��D��Ue@�J
ُ���
0�U��^�ʽm�J� ��~�g��N���M���ke9ߨ�dN�#Z�ן�'�&D��۾:
C?�<랑�99�E���
Y2/g[D���v�0�% �N#�[�F��n��$���`L��h�׆z�Tg�
�P�#��.�d89b��K	��@cϴw��� -"�G�_t��Ҭ���JL>���Or]cĐ$���*�}x'���`#5=���W�����\�] ��q&��o����7��1H�̬jP���	R���S����Mr�X֚:(����5O��"����9��őj
��&���͵@�m;�Gʊ�� �d�KZᬫc,W.��fI��v�l+MT[�sf��6�v}Z$�n��%Xڵ��W|���Չ��pV��ñԷH��[5ti�_yKd+��]�W�N"�^�\Ɣ��q�į�:��_7WLڄ��t)�R�B_@�n�s�Fl�c6�Jm.Ftܗ'�ۄ��z˥ٗ_��o��p�&֭�SU�r�
[i+�Q���o��]�(�s����yX��X���+�v��8R7Q�$���������A&����"7xj�7�5]B�\���<�u}0f�{g�Ƶ��L��l����ZҔ���'T��mW��^A`J��<7X���F�q���I��o�t���ߎ�u�S�@�!�cUm"Qs�Q;�Yje�>����/G8���`��b=]�§���<��~�Kxr3<Mח����?�
������@:s�i����]�5��4a'	�	�K�$~%)�qP/"6��&["(���z5^�^67cO`?�sc]H��kR�t�|�S��܅©'�d�Rʂ�c{ƹ����p�"dg�I��2�p�����7���'`��x�sE����l��׸�Q4v�Yk�xs5��f;@��Q�Y�%��/�i��0}����`]��2��Mޥ�%�=�:���y!=�_Y�{Q���(Rr
u9^0��&������xHm���bB���t�c�[/��,,��I�bKt���ydQ�[&1�-�P��B_��m�GG�/֪�C������	�Ժ��	��Q:m�[8)\P���h��3���x��_�%���	%&�%�*DzXm�\�4�2�8N�g��1��K�p\��\��;!P����Z�=�cO�E�쑨�r��ȫ�6'�X�$�H�Jm��-�MW#lc����+��M�'�VTς�Q�}�u�����Q~����%a�ڻ�&���X IZ)?9Gb]�\�n.B�cq��N�!=��`����r��VEM��3Aܧq�#4��LeJ^ć�>�ȕ�8��,e�J�4���^ b������+v��<Ua�E3��uI�|J�_`t��Ҡ&r\[I�pM��<hU3��'\ʺ�8�2Sbw�´�8��#B׬�ia����g3�-� ��!�Ώ�Z]`&������e���U�PxJ:����3�{���)|�6�M�8۽�$˿��e���`������5�ݗl瓛/ԣX�ڡ'e�1�"S���V���nj����@�m"�F2#5�}
��N���]��TkK�щvAd���2kR���u���v)�sw�}����`h�m�����bL�kY "���G����͒�u6K�| <�לּ����@�85_^T�z6n&V�����n�ŒլZ��(��/��E�*C@Ώ��IܣHJ{e`��Z�&d���R8VG9���6�D�(p1}t0+�����-��/��u�>G���因��{}���vgi1�1F�٢�XG̀1rX�����;�p ~�"���t�fi�.e��f�u:u*����r��⫨U�V�ϝO���>I	�|6�Z�8�T�V�l�䯤v��Zw�O�9��8�ɹ:ޢV5�PIp�b�|r+��Ce�˔�-� �܇�e�_Z>��[����R��=@��\hQ[=	v8�g���@��?�--8c��I<�.2H-�8��>0@_���t>��M�eU���\M�V���n_��3c�6[��㱆Z2�礩+�K��4d��s�F0���4���E��*��h
H�&���Bk=	��g|�`��c:��q���;��&����OyF���9˞�J[wH�C�˧cUSQ�$�皞�p���7�BK�� ��I���/�>���{_|哺�Sr��L͆�?�J��h�����H-@v���}�U$��K���ȚhW]����^�fmx�[�ͩ?�O���/�{d�S9"��Z�;�iExw�c8�~��^To��#����Q�NP���%#�����ol��$�0:5R���	�P��ؿ��[J
���$�v����_.�-�.����X�c&����;Uh��[�|a5	�� �?���ܢٲ�����Ӟa/�+S"=��P�&Һr¿!���
 2vРi	���*|ߥw�H�Q6��4����T�zV mۏ��]��1�MAhT�2O+s�?�{�><���&Њ��%��$��&���'aV�$�*e88����KTq�%�Q-�]��"���N֠�gu�ۮ5��~fYc�7���I��� ��4G�{�{�Y� w0|yEGIn��t{3l��p��:�	sˮp[�^G�iN�;��jǁ5��f+����ۦV�i�1��&�,}ba�!i��n=M��E�Q���X00�!��8�RG-�am��A���h���,o�6����'-J�*�1����d,�)[�Q���,�MQ��nţ���H�ה��
ɋ�g	
��S�;�����o��h��`ysT���W�k�n,2��g7���K`�R��J�I[~%�� �`�L�0T��5=�׀�a)[����BE�H��6|}�NZN;q֌��aS��ௗ#��ET�"P���O:J׬�3辌�=�� ���L}&
zCAoS�$L6�!�HM�L�8�?K�T��6igS�6!+OV2Ŵ�i1��,ߊ��g���GxZ�f�Q)�5h.) ���Ծ@�9fԳ��r�M�)"a/��B��2T�
�ԦR����:���o��t��^��V��Iq\-�,�)��M�Pp���V�OaЄ��I����	lp�w� ����H��HY��R�_\oܽ�'-��+(&;]nqX�+��hI�_�� �M��Ww��dr~�t�:�ow4���{KCF;?�I�J=
���Z*���]�'l��k�ρ#�ҏ-��潅M'�T}�W����[��a�d��*0p}����S3nn#I/Չ5Iuk�T\�����������k�� ǥc�3�F�4�,Q"VY]��?j"�0�-D#�6k��F��}��l�6��hO��<l���&:�A��.�(���Ee�,)�׳ fڋ�[�Y>�RG��1�)���U�^n�SOՔ�L�Y���0&u[w��F=��uf8y���&��/M<�F��R��G��T�k? H� �t����N����vѧOe3{��1�Kɤn�
��a�]�CV�}�1�:������J=.�
3`�^ �mROf5�
]�F� �@��� ���<�ѩ(�[9���`0=��3?Ig�v��,���cᣲ���F�]���K�m9MD�&bs&�hu�tZ\�` ��� �uA}���E��7
ޚ���aN���=��N8�S� ��Q̨%B��OF��2��R~�§Ƈ2�՗j��hd�mgƧ� 9�����9C�L}h��wrr�e�\��N�#�)���O�*1���D�.�cP����T�ߗ,�!%�8���Z�?�4[o��f,p�tp}�̀�D�NG��	�`�`븟�
^o�GӔ�Z3�;~�^�=	0ڿS��D&߲����U)�?�*��)�L9i-1b���$Z�0[����r1�'��1� ��D�j�z��ޅ�X2����p)���O�G@���| �@�����^�~� (�3� 䮰a�SM*J�oTV�)=��NL3�W�Pa�"�Su�R���s�(���t;�E@���? ��4�L B�x't��l�d�r�91FV�T7�'!H�*L���Gv�q��O~K�U�ڵ���v2�ҋ�l�XL�׳�߈�q�%e1î�):���8��;(>U�'�L��1�^��*�!38#4�Y�㭼<� z�b&t�6�n�9�o�$W�i]|qnUB�r�'^�� ���tc϶@�,y�}*K�ЯO�;�>�g�=S�M���h���6j�Z$e|~�AH'
풤aq�L�����3_E]�D�2������'�.1R]��=_�2��"�Hp��.(���ݥe��f9x� �ZMZ�����i�[��L"5��D��F��#uhg�r�=���Q�+eq�$L�y�w!�
;q��k2͒<HO'0�c��(c�ś򏥙���j�3�%W��'��)t�b�m!�j�(�b#g���Ơ�+����p�����B�e�5#�)\�tW�lgy����o�w��Ԗ���>+��&�~����a�lLӄÞ��nK��)$<U����Ê�T	�	N;��ϓ����L� ����
*[�UkVZ�����6ԧ>����q�����'I���[Q��'����2���ml��������&V�� >*NC�7����E��� �
||	=U�oIHRy#�F��i�rɄ�mfU����c��̲RÖ��&��+�K�'u<wa%yP�E'�o���I��<��l��z�,�:1�+��د7��7Z��@������\kW���>�D��Ф��p�5|��3;�_�0 Sj���5��6��n)L�rq�݅*{�B�N]�Z��"�Y���!J�o�� �r��c7#�/\�^	�;\��W���hB�͈�P� ��[��^ۺ�R��֔���x~b-�lŻ�Q�~��%��%���A*��K͈��'�+�=tK�~��~c�9AÑf
W	���t��L	g��v^��}��V��&�Ac�����_��l�Q��ٔIn�AJsE��O���o�v[�Z�=�����^�K��1Ӑ�&Z����������\N�z	
�=�u�t�5`��:b��y��2�f�V��#� ��b�Z^љ���7���[��O��ǁ"��|�	�A�!T~��J2�i���.���g�
1}Ue���O��6#ÛJ��y��qPo��^���1_��(���ys�9l�R�O��s��p��.ߍ*��šGL���>��j���T$�U��*DQ`�HP�t 
�������wCk�881�JV�J�S/0x&6Sd-���V)��.8E�؋~���*���V��/�y�!���g��W� ��8(��>�}��x�������생'C��w���W�����p�t�Oo�h�l2�����i������)2�3��A���T��E��]�]C�������������GK�`���$�yj�Ւ��I�!�Yq�o�.����|�@Oay]|��=��ZpKd^�C�	c��s�`(j��%j�ɏC�:��$��'�|X������*��k�eϮB)c�S#ժ�{d�uEh&���{���ƁV,q{�礻��|vQ� 	�q҉��o>3$I�0�]�SUwXu� �/"l��u�ڛ�=(��,�']�`��Zj��K�A��N���̪�!S,��j��,�����W p���Ry'��(�gW�-�`{ =�H�����.qH�J��䕼Eeد��RJ�FBM�t�����[	�W
�Ȟ
���'6�:���0���ms�7R����{�#��&�TiA�����/�����Uɽg��['
��_�)c;���=���?�� ݩ
1]sO٧.�);Z�yC�yx��!���{�pǪ���^���sh��d�o(�
� T s���������0��ptcY��dq�U6��Wa�f���B�=:	��N��
q�]ȅ�%{��ο�c~I���$ Z2��(2M�~���zJ��l��]�������-%dGL�1u
��m��*)��vǾ�����f��02H/oP�/��0[��I�H��u��l���i�M�w���F�f����-B���� /jOZl`q,�-Gݫ��A�TBy��$�]���&#�����g&�r�qᭋG\�%d��Gl�(�Ȟ�|��,������MQ�w���~�$ϙ$�u��l��/�&"�k�m������ZR�W=���U�r 	��ꮄ#����y�*Ԭ2S���3�>4ϲ�ƢV�1L�e�V�܆�Cs��'��WR�58����K	2i���eh�u��{�'G7Q���4�]4yΐ��Z�&���@Vi�Y��j����u*uI�Cg�*~������3G��Vy�	s�����S�!!U1Z��qBj+���2߅�"^�I��
���br:�`�R������j�d�̠��TE�j
�!@�qN�'��}�@+O��K�G�1Y��D��\�$�F$��/E�'9W0UGXZ��ң�A􊜢�A��IU�zKb�4��
m@Q���V������kz�;ji'���H�q-�Q�9c�]����I8�hֽgE�"k�2��Z<U��#D�4bj�b��sc�:^UFr`�����>�e�P�	�\,�f+ҿѱ���o�p�CdD���&�r[�@x�I����DcJ��L� _��q���o��]ѡ���#�v�|�̐�|	%��Q��L���.W���������BRe4�PZ���T��������=���=`�"��AIr�o
 ��!��bV���|ǽ,ǯ�����ZE�@�i.�kV	z��%��.�Z��jMƬlrd����\YH��߰����K�@9ҿ�m��P5@���F�ӱB�Oj���X܎�B����B�ݪx�,���t����yP�$|��cR�f���j'i��:�E<F�;a�]�ɏ?#�j;�K�5#�4���.yܵ/�^8*Y�u<�#�H��u�SEy��9XM��2	���T8���SH	?�I��1�{�ɺ<�}K��'�����9ǉ[����,j@�v\�m@Xc��ZV�j\�_e�ɞe��q�p�F�n<"9B�c#8Y�XPhi�Oy��'߭�tG*˽�"�6K�B��!?Pd���K�yA&��pиF��_T�i���Ϡ�O��������T8S:����%�W\�4�8u,Y~�J
��M[ �\/0�y |W則8nAڦ�Ϣ����SJA�+����;1ʒ�75$=Mry�:�B�F06�CA�k�C�`��*�k�)SM+j|�S���8\%���3 �p��NsP�>�-պI�uo�{��t`�*U.z��'�/���M^�h�6��J��vg�ўG��1_7y����t	K>>�K�����k(�S<cشw�e9��}�c?�-�c؞��������Z���ea��_��e�z�L�
�1V���=�o�h5�/<�(dX͋b%�k1�H�й�6W�
@�},O�.���W���.Y��]�^m�����K�����L�!E��ϡ��Cpny�
��r5�4��J�i%�^�8|�w��F)�H^��, ϛנ��&M�\6�����i]�e�5(n<31GEb��X�yG�+�70E#!$+�8�,���/�=6$��O��@8���'$v.��4�U*���n!�I4��\f�̻�i��F��1c:&�-� 0�ٔ�~F�Y ���;oy�wW:]� �U$��J�5��NՄ�a�4<)%��5��v9'���Y����m}H���V!��;9X�:��i�F@_5sD���� ��0�\z�ŵ჊�uE�2.j���ˆ�|C?m��0��ryWO+��f�6a�;�c�d����2��YOگ��}E=E�i�.2"��I���!�-�b�?���=�J�� ���ku����g7X?�9�&ڱu-v+�z��ׇ�\�#�Nf�埞��WO��
���	��4=>NSCa���(�w#�\߹B�����í�����j�J����yD������$(=�%��8��3�M�ؠ�ݏ��6���O�A!��%߀������ЅЃ�����������۳u e��=q�LF6p���%.���C��{+��<��w�~JFАB\��=��4�(�J��ݲv"�L����'��?y�Ï;��[e���	gS�m��z+�ObX�mI�D~�Kn@�a9���^#�[+�r\Tp[:!U�ӑ(�p�B	���r���<O|a++D �}��S�fͷC��k:�S+~�qa��<��b%׭^���#�xȪ��1>,8����u���Ћ"�����\��>h���ʓ5+�V�/�7��/�ӵ$��`Δ����@��
�% P�j}"�X�w���ۈvj��YZR�Y���&��ּO����,���z�&*_h��`����m|"�Ѹ��QC��T|�~'띓����K��!^]kclQV@�s�q�.�I��άU"Ӈ]A^�~R�B((�^��K�f8\'@؋"�Vvf�6ܸ ��[��� PC+R�w�Pw] /:ۢQ����q/�M��?�=�a��a�V���Hd��\���@�v	3�U<р�8@�H��|�'����9��!-��wX��7:��&_�ir�X F�4.Tn���������0lQVXf��!ĭQ����� �IN�Վ�舝���@�;c$�����XT��{q	;�iU�Qט�\i
���h�_i�uJ?K������6磌N#o�)VYxp����w6	�I��9���e!�W+����0^�Rf���/(5:���fo�T���vLHX���w��8j����N`U{�{sj&��H�c�&ע��ɚ�	X���ZR��������,��]�W�����H<+��.-�8 a�9~�۾�P �cEӣ�x�J��J�x��!�~�0�-������<�hC"%|K����d��a�&��F>m
-�U����OK}�v��p#A�"l&���6�qD�K������Y{P)������.q��M�b�B�`� rd4��K�8*������ҩ��p��f�'�[7l���P�����k��"��ѱ�op�rM�W����G����t�ר�i$/�[�����5��_zp�����r3���!�������*	�x�u��E^��m���Y�*�9�D���3��v��[�*$��7��a���A��.l��`��m�@q1-��:����p�F{I0I���d:B_���O������AV�X���\Aߜ_CG^��V�ƈ1$�#	y�s̸k�v	Px�1��iw��Z��_��l����6�9?㚰J�+{�������p�{q�I��mߍ�BX�T�AXO�n�uM��o��:*&B�ҭ�Eڜ̾���V���gI�J슇D��%}�O~�	�a"纖�C�DQ�� ����O�?�+#��X�/kd�N���'Xfm�J�bZ�\����3:	�6	�K���q�-1G�(A�����5fl�!�7_��k�_�p��+�?�'��H�:H�'���m�'�,q�\�A�$��'���ыC�F �5��@7�I�Q���G-��� 	R�}���T� ���BUc-ۓ��U6�f��{ҙ�~Fθ����_�e��d�D>r@�҉!\��� 杂�Q�����o*s=<�l�=�LS��F;#�|P؆Ч�h0���HqZ�jՉ�,����x䋽 �/�؟X�CwZ�Ȟ`s�}`k���D����1Tjd�N�ƀ���9ȔM�ሗ�"���xo�ʹ0���:�>��i+\��O�+����ʨ�p"��S�X�/ce�o����}�7�����k�Y�����,60s�-�3�$�n�I'�>���6�+��Q8�������S�M�^�4p~sp4��ϩ�Ν ���|��p�/�"�`��B~�F9�O<��3nB�?�`�9�0��h�Ƴ�Z���R�)@d�"�$�����'d���cO�'�4w.��z�s�ޯ7��_�hpch�x��[!�\��\!>Aǌ>>,49x�S!���h��oo�5��b:}�~��Su��!�Gx������x����Ds�P����:�۫F �����l?�U�fWԋZ	��~f�\�	IP9�����3�l�ci��3^�:D}ɱ���82�k]Eoe u���v<���Ii�g��_y�T�ĥ��j��u(D�,��މ���ɭ 0'x��#�GU��E�Oe��<��a�.+kzR1����8�@����0UT�/	0x��	�׸� 0Q��7m�^X��?�4�@�1^��v����׮�Q�u���YB�������g�j�S�ڿc]W����9@�GG���|.���U����9� ��S{����R�
	�������=�T���L�V/�ol���P_������Vf�u
�"����"��I�QW��qN�VўKD���5t�,���5J���[���a4*�N�vd�-wȅ?B�`ՊN�������.N�k�w�8�2�"�#5�mŴ?Ȗ��3?(Ψ�H��W*�BD�7��e�A���?��b�%X����Χ��!?��hAh� ��Y/_A8/zvu��v���#ڃ���^-.���	�W��E3yb����p���!��ĸ�I���Ś���؁��E��hӭ|+/$.�*0V�ji���i)"�{[�@4נj"-��Y�q;cW#^K����};�n��)���m���Є�jE��	�%�ŉމ�H8��C�e���`�:9�iDL��B[]���:���z��-��N�I�d�d��V�@�-�B|w����b�ty�jh�>����]C
�����zU6h��i�%�D��Ri�R�7�M7m֊�,	��p؜�H)1�sb
y4��M��}�o�(���t�GRx[g��!�2��@�m)��o��z�X>)�s�]�@�P���Q�5���ܬ{�
� A�jW?���Hg��D����1�F)9����=U'��j79�����~�lM�O�n�|�6�	�f���u�gE}]�-N��S_,��>\%I��2����#,S���)Q�Dz�7�`�ڢWM��������8�ަ��j�=�b���%��2�W��Y}D�	
ћc*��;�]������&�tw�!��*�I~>֒��Y�#(_�]�����+j<���R��ge�l��kD&?�ǒ�\o�E�մ2����Px�-�'�R0u�������1|�����;����~N}@Mץ���<����$|_�ޟ���/��P���D�|�Q��B�w����O�נ`T2�ko-���l;GҀW+���ֈ��%�y�`���{T:ը��(���V�2B�M�G�GV���·�!�^m����F��ɕ��/4'�j<�~a�V�|���o"0!T�3n��eN��g�E3���.��f	�\�w
\���3~�ֆzk����%cUA��9��ҿ$Z�ԨE�}� ��B�0҉)k�=�+�H�:M��롍<�y;nS�����/�psA�goъ��0^��;A�u|���Y����3���x�l�j֭��ʪ�Gp[���T�{Y�W4$S�;?�����<���y&O�n�������w�~w�RϊxN�l���bi=۽�'�S#�Z�u����Wtҵ#3)��$h���_Ms����W��d��8�K5�k�$��`�Uv�m�e�}�|z��)i"�12+��FĈw��ub�%t�U��9f�r1�m�)4�+���O��ꪛ�%���z˲ݦ�������p�e&B�Y3jF`��Э�(|��H�C��?�wT�$��/�H��t�9q�	�w��B�^�W�[lo�l[I���܆��%�KώV��Û��o������4*71[�N�4h��*|Ly{i�e���~�d���w�q�S0�-2��2ڔ�ʞb �/nGv�v�31�2Y�S⑴��R.�����>*O1,J;D�ZN��o;c#��z�S'�n��v/��lw_/-�ߵ�OfK��	��C옩�[y<4S*�Ϛԉ�P�VZe|%��x�뙵��S�\Zza���P�p��8���|
�l��y���m/_a��L;'���
�M(m׼�ߛ��ĵ;o�~�����m��]���4�a暵,�Dd�/��ֹ/�}�R�|=9� ���w�+�r�^�O8ft<A4_iaC���r?{%.d�o-�=��YdCʎ��� ��FR �Yl79,���6O��ݓs;J��l����EYlz�����?IЛ{����??����NW6�f�VY\Fk����CK\���D'��2���Y+Â���Hz;��� �MD9d�ʇ�,�MI*��%t����l��;n�-�^ L�$���K�+��|����Y��~h�J���o�?����<
�9����PK#nJIRW{+v�M+P����	9*H���%3L�U��O��[�3�ٕrT����uMP��*^}�Q�gեqM�on��&ɑ2���Y��r�@����:���۱�S��ǜ�A�1�%�,v,���+�X$�;+����X�oM��v${��ľ��x�"����K��Ph�M��H_��;�&�e���+�����|R����Vf߶%TwZ$��P;�n�4i���g��k3bu	K;���gk��-�h�������ҥ{g/ Gw�-W�5ֈ=R\��(5��	����x5F�C�_ܟ@����ʛX�|O_�f�CW��"j<.r+#^�$<Ω>�P���$�� e�D!�/݁Kb��Oj�f����Q�z�N�鿔q�p_%�ґ���Q�S��>�Z�c���/|����Yp P�4M���Kb!�9�7����aD�b�D㣰���?�)��mVD���PϾB\�윌W��n013� �HBN��#9�`����"��';����Ȕu�g(uXH$q��hD(����<Jo�#U��� ���X9�����ۗ���	�㎲-�� ���zl��W��+$aWrŦ��Ld\S�^���Ѷw��R(��@Scz��/�N��=H�S��`{�A��pj:��H�K���!�%Q}!�O���D�ƛ�x�̦��x����$�ץM���Y��ѣ+j�S��M����jU�@��G�(pa1����I1�%���(S�R�\Q�"�l����V�Ћ�J�.����Γ������ߎ�D�BvI�j�ƻw���t���+��H.\�����q�;��SC��8 6Z���l��s%}�9Q>�Xq��Ȥ��.��:1�����ɡH��͹'Q�4���,ؓ����T�Zv�8�aكU��+@pF��l(�E�]M�ț�l��*X�ӹ��D�V�Nՠ#�%={���K�'�[5��A��l�	i���8���̴O����M���t*��V�5��߁%�g��y<�M����-m���g�o fǌ�[Z�_��!�@�e���|��4f�H��O/$>0�����!��0y;�UN�����P1�f
_�y(s����W���m?9��~�����ᷨF 
�_�mڔ�7���`���K�L��o-����(	��I�= ���^8��̀��!-�{��T̼-�;���N�5=��9��oW@���Rtd���v&��0-^�������i��|[��M�"�u�X���X�@��U�	g���X�@��"�Q�ϖ�Ԫ�6�^6�]o5�n�@c��^ŧg$�[� δ�@�Za~��k_�@Õ6|��{������6�VK����t���h�9��y� �0Q�L`���/��4��Z�}u8�G��!��(E��7=�Pc��>9'��v̖��5�쇚�|nQ�Ϥ�0բ����	g�� E� ��|ʮ��L%�Z ���t]��� ��a�2" M�c��[��3�a�*���T����&���!�=�8�qJc<��e�d���.�o�s��HfO��@J�ʷ*_*iS3tH{G[:��,$XU^����C��I�՗}����n�(`#� ?ʻs��-刕������D��Y��'�Y��6҈!@!����2_���&:ۻ8�&�֥��7��jWC$������h Or����9L:��L���p�,zF+bOOĜ��x��}�$��4����(�t].�?:1�~"��V�����K�$$jɍR�ӀI�r��D4�[�lN���@�����P��>��{8�^���N%V+ ���-��}��O�B���_m-C6�֖Jv�bUۡ|�Ko}d^�%�<��'��3�2o|��t
�Hh-���B�?i�9bNl];��H��6�>���BU��������7�<�8b�/�Ӧ���]�<wV��ή�����L��F9�/�^_G�k�ɶ)n���g0�0.���B�'�p_~������g>�uhh
#�����%��̛$���!���ap�m��=���tX]^B�:m9A�.ړq��A��V�/��ߤ	"=�g�E|��ֱ��`ËЂ;^f�G1�q�r�&�75��&V8���O����E1j���Meuk��g3RG��,]�-�\�AB,F�t�
��>�;������u���T���@r���#���j�V�}��B�\!��	�!$�x���S�N�"leԓ���H��<� ����C'�ꜟ��55Bv�˯}���}� ��b��T���SX���h��1��t/��+~��HM�t̰��k �gt�;���j"�Ԃ���Uud�[����]���8�4Xo�;<{���O�e�·E��p�,���L�+m��A�Id��R[)�� �zuֹ�~�}���dS��Yiջ�?Y���.^�V��Z>ˍ5���3V��<-��wߋŢ�?��w%A�