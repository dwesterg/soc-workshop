��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>�����{I��v:?�BÅxJ�B����f�d���n�,o4ʣ�Rd2V��&����q�B��$I툒GM@�m��O�+N���K=��~���y7���{<�����(�Q�4�.�����BbLS�K�,�ݡ�&-��-��L.}��7I��L�p����U����eT�O`(+0�d����GK �<V"=����)��*������/����PY[I����n��l�è3��ML����59�ā�#k[y����%/�7��� �>�Ĕl��U�v�^oD�,�iي%�R�o��|��A�.��4s�����>§���ق����J�v�C,�!k M������Ѱ���N�.1g�T����)��&\e޶]ud��cY`o�j�"!�"�9��I���bJp؊2���ٳH��{] �G�
E�*�����Y�D�RpȢkB+��	y`�jP�A�k�����L9��0'&v�x���ي�ݲ`kȨ>��m*����9�5���Y[�K��;ďH�a���O@o��)V��$�V�W�/�1�}n, ��Z���R��1�F��{�Z���Y��{�+���i�8,	�/���\|k��p3J����epBfux�@��rEq�np�h��s�	����^.+#k��Ȏ��b�����@t�z���1�Tw�T��	3�a {�i�-g�z���t�,��x��򟛔�(���0ӇY]<�u�����8�y��q��ߥ!�r�4�	%���b�IꅟRY�Cd������h��ZR�Ԝ0�C���p�6�~,���!L�v`vCI�ռ�%�e�e�0# G�u��9��P_&�w߆�@�^�\�g��!���� cp/�5�����v1������ �h,u��͊��߶F4�IV��%g}��R����jBN]�4"�6&w佌�����kq=�a/��2y�2?�NsC�Ա�xvRy쬜���u=M(����p���@�r4՗�x'#3�">�#�)��~ϼ��A�rq#��5�d�<��'��
�+�R�mML��Ʊ/�~��V���X��m|v�N�/S�ڱ���[�����.A 
�ВUЌ�j�8�O�T��B(�6�u�~Ț�g����`�$�d� �'\���<B��0����������9o ��3N�>�ڔ�H� ��c�5+���E��߷pÆ�)rFb��
w0��d��z� ���a
��]ٕ��1 ��!+i�gY��P���Lz-�E��}iE��ڡ�nQ5&y�I�O��8�(C�T;ƪ�v�>�W���ʃ.P�At�	�e�05�'%���.͈�����j��� ��v,&�ihC4X�=B��NϧRR���Ռr��MWR���w��[hq�2;Zp�𶭋(.M���2�-��d2�.^��׺�#A�νcn���@��`�T���������H�h�����h'�C����ps�i��?t@�]��5=\&��~j��<�{���}�@��5��!�i����˂A=�U�젚s�$��-1����*G�/dXM��.><(Y��DB)�c-6�f�n�C��q��6:�W5Eg3�.-�B�Î�)��Oo��V4��{^A�m/�CK۲2�}$�-p��fU����.�������/bX���юM��*���^�Sl8_�"g��벗�e�+��? ��KJ�{�s������|%�R�l��	�՝,ϵCh�]�)���Ž��U�(�O,���;A�3�"����a�\�z��'LKa=�����5�4ׅR\�S ������t�tۅӹ��DpZx�&�m���D����tIF��_�=] ��{��p�LѬ�'�3G�=�a[�{�A.�(�1� ��c���ИQV_pm��ϝ�(��)���:]�Vr<?����8p��J�˞���!؁de��}�o���oz����ئ�3I�~�
iY��`�ZR&B�����CT�Uҷ�e. ���>�,����+C����]zɾ���[���oxh7p|�8'=���<tI�v�qN3�����h�LpfQE���u8�T����_+��%��L���Q�I�X��	�[��XJ��6n�*�ĉ� #�~�?x�5vY9�Q�>�;�r�ekU5)ba���Ya�4r�7a��!h�3(��M����%�"�g�X<��}��6����G���5b��)P͹�kI�)�So�m*��H���Q?�d��:^�㾰/�!�OmK<�q��6�@��#Վp	�9���d�V��\��I��(� օ.�OkB��d�ΡK�p̟����x�qg���3M�c��'�������$p�d���v5��6��?���$ �4� ��B-?��J�)���ڊ�H��b��g7:_���3�=�yG��V��q�O������e�S8EY*�F<�nl�ߍ}..�v�|����F���}�i��*��9*\1�W�=3��[v����x��2�վ<���qKNs���b�]8�[ɩ��>�h�[!��w�,�_BL�0<��@�)�x9�Ǘ��2���Q}�מ��D��Шo��n=s�n��"��|Z�,ȿ�%�����С�/�2)��d��)JX|?R)7ތk��R��&�هwMT��^x���`Ĥ�sEj(�"�������qqxr�8.<��s����`3�9���a��q8�+���Ն�/��h[܀.xc�jmV�W�
�-�>�F�,�V�����#��+�?��z�{�)<�^�7ui���P��>6T,f�l~;���B�p8mOJwd�NҾJ��@[�� v�8`��ƻ�.b��V����x{$��d��r_���P!�`�&X���]�U�9]��Db����ܪ��l����8��G�3�CHk��P���8G��fr���n{�&� �d���5�m��:��T9>�8i�GkUV�~>����)gw��9�
���2澪odm�R��#i(VyX��̏j���hE ��� ?�=�gXS��輫�E��-+q$߭�6�7�� �ќ����<���N��A�2U�-8$>����6����;�%��ݑ�iF�Ws>Q4*R��j$�Mp��M�'ƙ��,iq���y�G65�?�g����*���Ή�(6�s�.�[�����(\ՒQvV<�P	[�s�,�� �Z�vb3e�&q����{�;��:�!�.?�崼���!霧��F�J���_����!:��N�*�IQ���׌��X�A��(��j_�ȷ�4�b޸�)Ŧ���W�ԑ��\�g�#u
�R��=x��2w����`���HBn`M��P<�%�]ॄU�.��Cf����!��&���Z]Թ�񥯽v���z��Y�����߯M�#��d_����4�Pd6��j�NԃFK���#��|��>j��
��.?q����xm� �3����x%�����)(5k���oo�j��H
��[R��#LJ������H����D妹�$SK�U&���wt[��q.R���5=P�4K�G�C̫o5��%��w�S9��m�;/3Uj��ڣ��
G���EB5R�)����pƥ �p,�qo���������
şY��/ �D�K��ٹn�������5C�e&�=�]��� s��ߋm&��Ώ��qxC�T��4=�ߥx�O��s+��TO�������SU��"��=�g�j�{wd�I�X�?�:C��Q��a���*W�/8s��;��O��y5����H2 d�X�/���t����N�xO�Z�A/�H���ڮ�Z�q�r�ұ�]l�X����tR�^���i�Z8[u�\�����BF����	�75V^��Κ��3aB8e����W�AZ(e�8�m��V ��g���I�ȵ{�i h�?�����r�Z��׊]��G,`�Z*���Aj*�b�4&��~[�0��Ȱ�����loR��as֦J�Ό�a
u�r"��]��(� �/��Ŏ[�C;ms�̙9ﬥfPO'�|�W��1GTV��e)��ϗ%t�S��0��� �������d����~o�x<�$��5�jʿFXn�P�0���A���^j�ﰏV��=m",�pL��&do��l2�_���=�`�U�$,�O�)%^|v����w��zq���C�V���HAi��f1����ߏ����#x����'��:�u�����!W�� �q�TL븳��K�.��CK��i�&������f�OT���7,�&0tU"�()�#:�Dm�}��!SA�(0p�h�,9�b9��vA��<��H_��GUI�:�,u��'�xU*k;��h8�z��<ͦ�	������*8� ލ9�g��KE�()u��*�$�u�7��oVQeH*�7���Y������)|��ʢ}麎/�_v�Ҕ�BP^�t
��xw��A.�����py��S_o��|��dB,k3xh�>BԸ
�a$PT{����t�[]}ӄ΢�JAE�׹]���-��<O�0_M틩�3B�c�C���(2�F�/a�>ufKb>�s�+�|�W�ϟ,�=8��o��M���[������/Į,���h��=c:<�����>��l��e�F�M��z�`x�q�JK�?��˦����o�P�H�U���� $�]�bcļ���g�k?��ۭ�>���(}Kk����{�޷*s�A�M-������M��^�m�vye��5����$FZ%/#6b�:-�H� �W���<
���iuu���2�Ts��l�kk��b������T�+t���e������n�ͭ�,�q�J���,934���~����A��RnwI3b�0�`��j���R�:��cpK��4�A�u}�{i&�7�3p���p#K�&k�~���ވ��l��������5�Z�J(�Ö)���*H��Eꝲ����#pH�q�w׺��PsAL��~*so��$k�q��+WX"��>˲Z6˸q�Q��CB���=��	���>o�7G}���2p�����wA�?ۜg��_�udp�I���"��5c�ɥ���Q[� ��t�+L� �}-��x�A�E�{n���P��P�|�+��;(Q3�g /���@�U�����&O�^�-�e��>���n�DSy�*�v��o�pj�Y����*3�e<6����FPۖ��e�ƛ��Ewh\�#���?�֐�������#�Y�8��ƽd6��6���ۘc3��ڽt�;r��[�d}�$��!~����B��o!.{Vі�8�ԡ{h��[Yas"���PK��8��ڟ�ې��19;���(�I*\��u�|E]sZ�5���&,ڌ9;*<R.J0��KŢ�5;8�O�8�<ߝW$~������}͍��J���s���s��09ʲ���zm׉&����4%��?���^��,���G�DcU��DK� ���I�)+9ji�h�����f�m۾��/�H�1ݿ��o#cO/�H�V����k�,uJ]�	�h��>���\.�x>8J+`bVΒr�����V�D�n�m)2�����ޤ�֏\�)��z�O^�-��o��k�}���g���߈��Wl&��~��EU������.<�.�2"�8�H� .������m�8>�]8��+m�5��L����$~Wz��j������:qu��'^�� ,k��;���@8�-�:�īu��_����d@x�(C�Nq1PG�g�˷����)��Gm�	�rN�X�<������_\(�e�E��Sdl�LZ�]�^Y��QZS��Ʊ���_`� ��,�?���m|����cwjy@ED�pe��@�5u9e�Jk�?���k����YN��7:�/g8u��P����o;�P�?�*�'������_]�V'W�O��%�摝��2:��?���:�@[�D�����}O�JF���3T�8K��$i?�V;��Ŀ���4�$����_<����u�дL�%�Ӣ������(�8�h >VT�ԈGgABa,��qPA䏱�2d��	�>�~���M��� 8��DC���	�p=�m�R�ne�8����w�P�'���o��C��7qu���кI�i�e�n���@�qa�(�D�`͖��;�*�m�]hx��s�	v��� 0���T}{�WIǚ��~\���m��%a9^/�
f4�:H'?���.��[��qS�{����&����:�8�c�}�ѡ�$-8/j���ƉN�Q�������.#Բ�+��Ow�se�_ː���0�N��N(�_�_A1����y�/���Pn(�������Ȫ>�Y��z���V���J�G�4M����{,��N晑�[X�8�#���=�G�&���Iř/�vR���g�e_����p=K b�\,��7�4�WO����8��~�O��	J�|�c�% ֢�� �m	T}N7`/�m�M�V��B�Ӂ��V���
�`�3�_��C���6�ɝ�!�;���I�ӊh������&,�8����T�n��I'b�c�Wq�{�����D���S9��D�[dY�A1����!w8�W���}��h����Aǹ}R�X�!��O�o܋&k�|�o���5e�P6N�߾�E;�+�Ɣ*�]�fhOj`ˉٴ�Q�>��F m�4���]T(P��=)
�R~W��YPF5��)�?�=0M�Ăsѫ&r�2��'h�K3��+:��;	*�l��K��vQ��,sU��Q��<H:�ui�4�.r�p�C���|:�n.�i�s�u3S���6�,5���� �����z���@�j0��g��Q���z28� c5M�n<��7*2��3��OU.g\i*&ˍ�|r���[���)�����4���,�׎���&����stIZ��q��_�:�f�P����MW�|���~ڞ��ȹ��7}�(�����E�n]6�gI5.Q�r�%�����ƻ�4h�^TNp�,�B����w#�j`�swD���K$~/J�e\a>����E���&0~X5�F'���/*�D���k�mg�3ٜl�*�{˙��ne������F&LwH%0얇�"͛��; �^�m-0sGڥ�b^<�r[����<v2��G��R<En�E�]!(�$��JÏ}�P���-�lg�5��`���iP?�>Dq��<CƲ����ΗſH��)�咠�Ȯ�K}J�G�^71��9�*�8}��tEӔޯ�����`�,����8�����p5��(��������=5*.����b�i�X��9��JA-֟F�Sp�� ��4�P]�	1�W$f�R \�r9+~��9�i	��C�zWb�{c	G3��K��$��C2�J�\��K
]�r����^TG�۵����:��f�rm*O�? b%��w��0ؤ���ȧ���Qc�!�@�|��t��c�)6՘�6����W�Y���J-=�N�8��ˢ>�o(uB��Է_��~(!\w��g�<�����q!j^p;��N@t0�S�H�� {�'[���d�$lm� q�N԰��%k�8��@0��d��F����V+O�
��F�
����u8�ίk�$zht�-ԗ�F�B��L��/ޣ�q�P�*�Q����E��xq2��0H���l�+z˫��cൡ�=��_�҈\$S(��^Q�@�0�8лBgɕ�Hʄ�m}��(��zc�-;�.��J0����NF�]�A\}p�)3�e����+�VR�1���c�V��^�V��Mc�Ӏ�o��7��-����"���g��p�W;���P�������8�L��9�7B5&#��1ເb	-��>��"�LB�w��{R9�yj��[�R+C�	H��.�|��"=>v:0�����jV�v�,�>��	SԐ/3�L�:N����8Յ��V�a���4s[A� ��(,�ֿP!�c�_�V����`'�j��bC�;�T���-d�����O�8�3�ڀi>n;�RO~4��=<h �x����b>��� s5q�?a���麃K�] �tE���$�wo�3#*?`o����nv�i����u
�D��x�����F��4��U�{��þ5�᳐�6XPxG+�?rj_D%�\nb<���2��<2�\<A�A޺�#�e3�ĹQ|B�-`P��I�e��oj��N�*1e��];7��In:�y �;�_J�݉P��{X���Ip������K��&�2�a��"�`��W\��/��9 �@�@ ǈ\������<��YP�����M6}A��>����4���M�I��{�Ց<���	��ȅ0lD��|E0�t��j�j�
|w24��*Dch�31B�$��U=��1A�`��O[�<������M�2��{��\虒���&�Zm|ᤡ�ө'�=ڠ��v堒�"fj�T5��� ��&�ܼ���	\|�m6/�{mna�m�)`�z" .TE�Ҭ�;|rE�e���0�f-L�ܶd+��8�뀈�VHq?Qa�<����-���@�z�e�e;�C��/a�������k湤ߒU�𔭻-�wߠ%�S#ǆ_�k�|h#5�5��ov�J��Ȝ�V�ikCX#<�6�����_UJMօt �N��M��tA4��N��z���L��
�1%)�gC	P��}̟��@ϯDJ<=w�'�.��h@�A1�e��ߊw�P�����͓,_EԬEK�����������@��gMi������cS�V7.������o���P��a�Trt ��t֠��
���<��Ŏ</�l/�I{�n���z�b�P(�^��,����R}��t�ѲH�w�A�A&[����<:R�c��	�k��+kD����S�"~��1������-�2�1�fp��out�AD-�����W=N�����zk��1MS�ZÄSwj�/�ly��R���JœNr��.�~J��������̎b16�d���aM�o��y'��3E ��������^��=0/������rb���\U�ؕ>��|z��X:/[���hX+u#9�7ú������oc�-z5�tF�-�2�vM�-ռD���%�	n���@_�'��kMa����w��Ap��CinU��;?�L�Z��*�XQ��z�? �g��fq#�\�����2X� �w,��S?s����i>2��#H�>edRZx���!5�	.�0�o{[v��^��Vk;K�\����X��UV���}g3!D��?�q���]�Ԥ�F�#)p�f0�
$�e��ފ�ְ��}T�`��&����<�O,O�+�I�9w%?�؏�hg�uC�P^{�����W }�ȈD��u�@����� ۨt.�cn*���EI�o�Y;s�l��@;M�Sp-k�}�[���.D9�'7�5��V&��>/%.HAu�ٺ5��3	|ֻ��=���`��`f�"����6�U3X�'Ɲ�]-A:��|ou�Şꪏ݊���2�ވ�"�x��u��̥�z���#y��|�����n��rʷ&�`����E�2��UƼ�|)#n>T��7�y�3t�g3��	M��V��#8���3`6bO��Αd�_������ ؟�X�](�Z��0]N��~��W�y��񺧝l�ķ����v���������������x���lNl�kd*_��/�o��N�ڿ���%V����7��&8��u�Wsӛ!�\nJ|���x.�E����J��Yf��xs\�v控,I�����!;��v�n����X����Ri�I=Vo��t�3M�n�t?�@	�Pl�ʨ�������«'�P��AH�Fx)'�%�� ��!+lg���>�?���'�~>��]yp)����������<�_c�p��1^�h]'�4�"?E��o�R�pKع�E�%�������t�D�8��I�&4��Q�w�施!~D��h5q
:�H�'��9Q"�,��V3�d� B���"\nc��^�H]N�#$�H��#�y~����[�#A���[N��Y||�7KۙJY��B�� ��
�C�a���Y_����CsL$�J��O{H�$���X�X����t=<�{�5����f������-Z���#Z@nE�������71�˿�S���� (���B<��5=�p[0b����K�F��$�@�*����x�z�t:��%αT�!c���h��P���8�(�1�p�W���CU���k�|������Ǒ�x�Ł��2��Y�,p�d[\"��)iFC���C��Gz�~%�+��r1�'��N������P;������_�����F����|�u�J1����F�2�X�x��,ZTMb7�rܜ�d����s���-`lF�W gLi�����;ߚ)�e6b*αƘ��j"�1:	F�gs��QF�/L�"t���x�)���.�n�A,竡{�N6��\x��!�ޭ,g�����y}cF�9��r�L&�'N�W*c��!)$�K�lj}�bʿT�8�8��ꨊ��F�C�����/k�&s�����xV��U3�K|�4`�@���
�t���C�U���?�[:��.���c��Sn���h�s�?L��*d��ۣWh�P�����&]He�G���j&zH�{ػc�誡��^��o2�p<΢�2�	p�g��&v
�"p1Z�5���.�� V=�d���U�p�߮M���9TZ�5Ɂ��b��{�g�B���H�*��Fw�BM�wI�u�>���H���S�D���_��a�{r"�6:�,ÉRKly����@�ٿ$�����KH-C�dɋ�s��4�9�����T��$�f��$�)�D@��se�!(�/���*;I��8����;��������lԯrf����P�p�-s;L�`&�p�f�a�,�^'�П*	ǧ�N�̇C�0�j�~(����G�@�A�7^V~a��O�i���Y�t�"���̘�b*[	E�Z�-}�zߥ�"�6���<�|��Zkvl�8qb�P�W.-����?��|zG~�?遥!s>]_��};.$�5��v�nޡ%i�)�Lڭ�^'?��f�����H:����j��A~�DB:���z�$Wfh��o4%�ʣ��J(�'H'�2�^t���|� �I=��-Pۉ� �
V��t�ܒ���A�T���;�֐�`����<mC0��^�D	� �.M��A=st5��-F�k�*䳐6i�W\��NT��H�t��5��D,��c���7���L�Kȝ;�/����t\*ۢ��$	�$�Z��p��e��������PWVO�כ;��q`]ۮ�	D�65^pYE�LW����e�7gQ����z���⻬U�L,����,��L'�/Ş{�8� ����#qd��׉7:��mL�M�ҙ�!�R�����6�j>���cۙ�ƙ̈́	��IlP+��2��j�O��5�ms~�{��4#+X�{a(\���_���7H�$�}">̷ǎ����.�E�%���^�������ߠ�#��D�s�v�%�#Y�@ȁ���$~���h�{q ��?P���!Z ��*z �3��;ku}��p�Y�&�)V�e�~����4�L�P����j�J�9�]Cњ �%E2������R�A�RHZO����M�yIZ��D�s��I�-u�U>fM�z��x��5J�M�ܾD�#Tj�!)��G��u<���׾�hU�Yە���J�k�!4�`��6���@��?UĢ� <�2���>�0Pq��g%p�R�R���1�`E�A;��\w�KZ�?�:,+kI�ڄkm�^�+��Cn�X�� �װ��q̷��
���IA�Z9�9�W>��� ���Wg̍��BIx�l�����L�ɡQ�a����"x�����$G�b6�yee��:!<L��xf�[���e��=qw;]�v���H	E'���u�[�-05;H6@to9����z$M	�T����j��L����廒���K�����R~a�^]�S������ ����-s����;B��q1l0����[��?̂�8x�D����p� �F�?#��E�6Ɲς���|����ɣh\��ǭ����՝��9q�����/�Z@j*ǌ,���&�X\[[���޾h>����e����[o0��ל�x��B_$]��O��^V�?��!""|]�0����CRw�k2A.7����z�?#R�>��b��cǀ��FC�Zm��Nk#�aL��E�X���&`>��q-�Fr®QI�i�>uRG����k��=�M|?`�*�8B�� ����uiɓ��~{�%c�-�H�`�� g�����w�S��ʲQ75�?��F�x���h =��������'�d�1���r�����5�\X�������o�+קNJ J�����ݨ��K&_�������K�^cI���	la�Ӥ��}ߎ�`������>���Vj~Ty?d������+�KP揥�k3-h��ͤ_���7�]8��C�����T�t�]���Ç�|L�U��.�� �Dq�%tٞ��P�~����(�{&/�	A��cg<Z���؊�ײַ���x�W��l�<�Tn�B��1-��Z|4x�A��� ~�L7��(QF�	�����&��S��6l_\��}X�X7%�cn��2�֭���/Ȧ�5����h�FϨjO�<�󊗟g�^���nU���IE[��m�<:�Vd��{���n�4h��������\�5}ꄹ��k?C1���^��v�tH�,e��#��7��%���~�a��=��N�"! �-�l�d���� �K3���VcyC\��RH���9��w�o{�,cY�7���(��X�������-��* A������0p���@	&���O	JE��4���=@^���Hisk�0)���g4�e�!��r@]P�P�`�u}?��*�6��ِ�,��,�u�W->t�玥,�{�/\y�\p�iSFo�����ڂԏ0�<��Q0��j-b||mʸ3G9L�~�D�l���$�o��x����t��v�J��x��2/�)1����+���qt��D�ĺ�5r�zŀ^�<o-�)�U�"�O����P�����(w�
�&l��d��6�X�k��&�w�W䲗����᪰<G�@����vYgΪ�C�c�<_IM�"L�>?.<1��!E~��p��$�/�9�҃S�*4��P�b��c��3�54�\�6�H������=
�&�8'1�p��f-� ,f��ಒ1�4QE| �Y.�ڦ�� ��9� �������.ߩ�p�{o|� �����^k�w9���탬2�CՅ����-�?�u��/ĵ�Pj;x�L�*�A#���{����d�k�L�������j���r�5e�Ź��[(�_N�lV��_޵W+��!�j���y�H����u+��N�*�u�+��Τ6�vm��O�˔<m�ϝ�=��%�G�[n�O%5���-E���([0�	�܄��*,�e�%��f~����Ε�6;� )�J�N�-�7�)U�~H�w�i�JO�qfRM ��:2�	�ؚ�;��H@*�K3Qq�bJ�r��u-N�tDfU�������ӽ�w�>��!	zv�a���x�7�LF{�
��;��.뀅&����w�o.j�]�snN2�C�i��O"�N}�'��4�$�/��ײ9)}�@�F�5w�{��Fc�OX���OT\�*(�7G�-"B�\Zw���VK�q4���M�<��xӤT����LxRc�����3	F�(U�
���H�
h<�OA���	�����������~ҕ��/¥�CG�j� n�.��2�����7%��w���h|LY��)j��]�m�K�����5jȝ�
�hZc���zG���!_
[B��x��3ۡQ�8�� �]�{iC�@��&Ն�߿��s�������_���G����n���GJ�F~u\�S�*ř/xIx�`8�(���5+[��Ͼ�Nqlk|�jǻ��3���U�!U�����T���E���{X��m�W|�s��V2�eU�S��Xm0�8��i6�e�
Ł���⫨����H0�
j|�xڑ�@Y�a��%v�̔�.�\x%�����^���F��:Wu��ܮl�bd�cMч�
��P��QZ=9�j��9���r5rM��+�e%�@:nW���t��鶭�-rf%He�a;zLRAU��uv0�G�Bp�V�����ND�)GT�&����p�AZb7���kl j����d���t���#��@-V�}�>ܔ^q�����q�h$�D���@��k.u,,[b"����/��$p�Qu�XN'�`-�.Uh#���Q���T�	:���*$�`�>sqM����`-�.�*�]�3����փXR�;I�]u�C�%�vţa���!�3�n��/��~���`jX���X���R;Ҕ�1��H�`ҹ���N6�����ap-�E�����G����6'>����{��ǹ�5���:�E��\{|#jUM��N�{�rK��
@�YMYz�r�Y����SG�9:�T/OD7ǭW//x.O�U�=�{o?�|�ZX
 /�t��%"Se��Хtkm�c;\P���v^�~���)�w��HZ�b6/J��E�1��2��cЇ��	�ɳ3cݙ��}̢]��+㻮r�[lG�Q��h����*�<G2�0l��b��p�:Z�{��x���vu%|������r��Tc��п�n����}�o�r�L��D���R����u���7�yk�ßu��r�]vz��g�NvŒ"�G�V�>x9�L	�ª�O"�o�����7�aA|��u�qžv<E�z_� �V ��䓰��-p(�k3ꀾ��kހ|��s=ʧ_W��d� "�1�&H��R��)=.~)�Z�Y�{���ս��j��	����Q�d����O���5���lW�z�3�95��7�B�;�����N��t��#I�X
��������1��[9{?��z��h�k9�&��Ђ��S�Ӳ�%�ؚ�gK㨏��=gHb��Ѿ9�)촿��"T
�S��a@�S�_��`/��S�T�����̜9c�ŝ�y����[���j�¿�2��g����$�;�9�;�W)���)����L�a2J�Z�ވ�E��S�8��D"��lAGWԿ|,�x�D����������1�O�����</"�"��H,���#>(Ɯ���֌=���f�6�4c�K{�
ù�&l٤��z�,���(�FY��(-(-�L�:S;5c����p�\2�� �w .h�[!�&R<k�@�|?%L�st����͖���W�^���s�m{P�ty�w)�Դ�W�4!�p��V|�"q�7d:NO����K�Fu�ŷk����n�Bz?�￤������o���YtJ
N�6,��4����(Ԭ�a�"�\m�*����BBw��{~̤�ɏ���P��I�]en�עQ��F�F[.7F�C�xw4�Ӽ�qǷSz�K�J�:��""":�A�N��i�B�ѥJ�dZ�P�S��Ku9�3��E�0*Z2�d��#���5"OǄVp����K���2���7�;��g�l*�\ ��W�؃����١75"����R���0�>7�v�۠�d"��x��`�����n��f9��PxFy�cZƉ�el���<QE��%u�R��n��|3v�,���qb̈́�$��I�/�猴�ZH1x��c��
e�݅���&})�aOC��1:�� >��Y]\�cV����:)�,c LNT2ߧ�u�lW����k����nt�,}��V9XL���r.���) �zl�������@F�E��pb`킡����D���\�UB?�)H�4"W�il�i[�b��(�ܖu�|�MPr,����@�JDʟ�G��<^$ɶ��JE|].�Q�� ,�ka��G��	O��~�;��j-q�<㦷��ҜNk�?���۽�J��9���.�K;�~��B��O򎆾c�
��w��h��ͦ���fҶ���F4���7�p�(�ס��"�7��M7��^cq��!�g'�� ����Dթ��ĝ,�):�^������Q������`	 ���׆ۡ�u��@�X�c	o�oJ����uU�a��s��M��t\�����ţ��� �]��c��UB�֣�*%�*���ӲX��7�N=* �S���o��dʭ���o|Vt����Y��a�1�v�-�[~���N������x�܆�����!�t�@�3��솪L~�2��l&��?B��@����`+���z?G9��hq��C��1�0iK�X�.��;�G#i�N�b�Q^��g�3o�n����DHc}S���ח+�5<���X��.D���<1Np����:L���lyum�\~��)F��0� ���a���}o>� �z�ѝ<�˴O�xXVP~p����gPZn6r_R�-ǀ���Z�Kp�;=&VYv��ܱq������H�h��������p!"��T�	HQ�j�2T6o�UbkI�#���!u���4K�땵��}��T�����Q�7W�
\MT%����t�f`���RnL1���oL���g�R�]��\�m�bIO�z�M�S���W g�B�e�%�ҕa�Sc��LW�uk4y�s�P@tv�ݯ�ѢR����g����J��q�Yd�բO���)�I�mI���D
��sVls`��\�m�gG�\hx�����`Y�)��&0f��k�l�@]��~�^W�"��R�~z�sF)�yuƟ��hiFdj���- )Y�u/���?<S�0�2�`%��P�#�(�@��=���H(�����{��&2�صg�L�T.V�=�i�̪�l���fD�ޥT͞};IGTʘFB2s�h�p�(YjX���W��� �$��� �n�0�Y����N�����1�v�=�Ta?�u��*ȘX�C��-�6�4�W}c��n[�ut��a|_�����Ť̩�4Ԫf-G��-����Hy�v!�J[Lu����9�ظ�"6j���A�4*����cܡ���y�M���tԺ�'�����u��ˍ|be6xG�'�12�&l]�ڶ=E�wa���4�����wׂ�^xIq\����A�v�Re���y��}�i��Yڞ��6���\%}0 ��-�C�_�#��� YZ� X����a[ŭK�;*	�$b)�4c4��oV�v�����Cÿ͵���:����&���d>)�e���,���|�Ɛ���<�^�q;�ֲ��8����fS����XE\������	�ӱ{C3Of5�mq��2W���~� h���#��d�_�����*�S?)f�Mm
� �e?:�'E�q���v1�7�(6�i���91a�1;Ғ���%�)*eF�`��W��ፃ�Q�;Sq�V!�9R�y���s�ᵿ^��dB4�?cp ���:C�n~?�)�L���n��6��jEi���
�y��f����$�	- Oj��$��@�OC��R�/sB3��v��54H��񥛔-�+��x�G-~��z�����6�Utȗ(�"�j��eEpi���Dg��Y�$[zÅ��XJ ��b�SY��X��7L[��п�_>�#�����|��\��������Zǀ	|��)��i�[�8a�I^)���6���Z���eL��w$}��âY�Y�x�A�!c���2#��m�X�vX?{�:nnݻЖ,�]b-��,7v���aAX:��ںi�"�m�ڼ�=�i��u°F� r ���7��KY�a�*A'��샙�]$�+=C��{k`A������>��7�?���SmW)����� 'Æ���8��3����cd��V�)����1������Hir^B���� �� ��mDr��cS}�Sr\KX�*��cq�?�$R󀺖W 9+�G?�g��"�g߻��m^�d)Ov�Ux:�ϝC+��)oJΎ���B%�53L�rM}��_3�r����Yt��d�߇FJV�$e�LA]Eq�^�9;⺊���qxH�q���, �P����j,�Y�l�5�{��lߡ��e5@��'� �6�u}��2�Fq�=W��e�p%-l{=@�+H��O��^4"K����K�_0۔��"��C�:D���ll��s_�Q�AR���hTk�У��Sܨ�� ��.|!�^q7�t�<2\��#3uIm����A��:����ؠ��W�/Zh�	i��
('9��:$���3P�7͖M�U2��N�sW�z�Cq�a�Z����Tu����˲ų�=X��ܢ���E�7V\��#c���'��}�I�_�:�� �_�yڷ բK�v� C�eՉ�B}~I��Qb9�)sO���{���ٕ���3��WW�X���ē�� K���i
���6TM#�T�E�2�=���jp���w�]���&���G�l���"����	d�vw��D>�<��p��o���N�I]�Au)h���� �;4�Vٰ�i]��6���u3{��o�4�o���=��&�fS7�+�O�SX� WZ�,�w�Z?`�c&���%$l��H}4%��qŴ���SD�<4�T.��c/:�]�2�CMw�$+��O��5�g����ˉ��yp6d���thP,������Z����su�(�v�T]�b6�o��i+�6%<���6l�?�#(!��\�h��qǐ����&�l�.��|c\���Rm8��:�����#�ګ�$p���ֽ��+٫b���0'�tv���/�꽙D�ӯ�AO�|(l������
�l'ݒd��x¦z��%|�~Nl;3\o�3Xg� �!���y/q��´�Ğ�0���x�Y�۶?
��D��]qϴ�+���]��%�4C��9YzH����As��B1l�B�S�W���
��t�[��t�a�*�ٹ)؝0&ȕUI�Z��m�����[���-"�D�^��ѵ`��7�J&�3�W��ږ�z�cY��з��<�4��P$/.Lݫ>���gX�'�Ml��+R�	FL�~|8�s�l�n	Re���gW>bT�.a�d���T#�zˇB��=��eG *�K�����$�W7>N� f�B	�L8�2����Z�Ԙ�a/����yx{��V?,o>����F�~��eœl��q��$4!��.C�����[V@�Kz^�`����yuIT��+�/LGR���!����R�]W����ӂ���5B0�������ȥ���Ov�[`�N��v�[�J(ᶆ/��d�a��rɴ3��qm�����|�e��n)��Ī��e�+:u�]5��%��ͽ�)����x�-�mS;Fe5C�H�0 �����M�E�V�=��ro�8������⿹�I���M�X��F>����$�(���� �R���sq�8�a�q��@o�J�&<i�|���cg���3��x��x������w�%�WZ3���� �S�����avF���ߨ�re�D�-@Q� (u�i�o�|z��<�����$�u30�[��G3Fϻ��/ޝ�kJ9g���)�\G"�D`���8wo{)��wH7J���� ^� Lvz⾆�(���	o���5�A~X�]�!Q�Jܻ��q��2Z��y�}s.�>*SbkdrG�a�`al�����Qa~~� "O�K��?.�?^�'綆VSx�B\f�B�њ?����7
~���~�;�%��M.4 6�=�&j���4E�̷^}�M苗48v���5b�(ސ���KLv@�q5�ᶴݢjIB�r�����ގ?F��x'�#��Aud��\<���Ok�HC�UD����K�P�bsI4hd���
��ٯU����L��3#B&�Ж�z���VϨ<Aױ_\�rZV�,C+�}���r�z�����N��
����7W�&5�����A��N��~,xur��A�5���sv;/k)�M��T�[�oz�:p7>OJ�>��1L�lI
���S����Пpm2Z�����T���ӾbK�8_Ώ���Ч��w���(���I�@�d@.`�R蕠��5��vvG��T��x÷�N/���ԑb-��|nJ>�3nE�򦵒?�� �>(�D,��栞J)Q�w׍e�ʧ+)?�^��6��a�eo�}ŌB{rDw���DZ��0���l�L#�Ş����o�g�kr�A��{�w�?�`.�&4o�qlʻß�Z HDz�#�`c%��\�DE;����R���C-E{�d�D���
�������������"mxĿ#'����D���!EQ� ����n4_��G�Z�C,&�����]�.P�oFM�#A�@H��lC�)|D�^
�_����j_	z� ٞa�������ae� ZV5��Q�C׫U"~�)�G�Q#�_F8�-���"�W�5��@�؍�%�S��v��	����}\���e
z<-��'W��.ќX]Ҵ8v�={	^<}Z(��yլ
�7.�:d�h�/��Z������+jߍ�G^C85@�S��Qh9b�N G��I񱱧p�HU$[��F+�F�0��P�	��z�\�R���v]��뮾r�t�^=��aۛL0�J5���
T�͵��7�SD^��Y�)9�H���e��<�u�P|��Һ)�߿��]����[c�^/��.�����H��u)��H�c{];u�%*H��h��އ2��Rb�
P��/AF�j����]� d����'������GJQk"����Щ������33.�-�a�cROc}��b}��^���C �	"J0Q�xB��7�@>%���L
X�2
��k�Л)��[�}�O;M?�x؍����S�P���9
�t��ҍ�1�q|_�h��\[���
r�$�ԮS���3�#�������F� Y�tW����!��ރu����v$�e�w��6�H��>���;��z����4S��P.��"E�m���\vu��Wbr�5@f�D���~M"^UyB�r4��zY`?��z0� s�l�i��Qk|Qʄ�ZEeV*�Q�5��o��1�C�dI������Lr~T��e��f8ԉD�q�!8��ug
�h$*f:�T���!�ڗt����g��%��"�'q��C]�m�ڃ��:�?+%�Ǡ��m�Y���8���W��=��]g�:�s)~!v:�p�ũ>`�� �9�U���]Oo�>ᇡy#.4�yo��bH2.>�� $�'`;�q��;$b������; �	��\
_hMW��i��rl�TW��w|j�J�/c��b���T\����E� Ę�
�{��c��. �.�Iz�M/�0yJ�>_���b�O@��������*qh�v��]e�{-����i��x~h
��>���P+�f>�5�17���|���.��M�*`]�6�f�N>=r`lJ�
F
��&�a��M�SJ����ѹ����Nqh�g������_	;h���<v�=�Id��f��0x/�6�^j9ӹ=��/�����}�,q���G�i���ߐ62k����/�uL:���^�R�V����w�S��YbD��<�2j /��8w˓j���傍��O��a�7k$ꑡ�_i�H��8&,�\�vFm�� ��soӸK'����/���)[�����e/
SԲ@�MR��x�:��$@"'��,���H$HߦrZ+�mο�-�iR=���䠫i=�`�U~`쨾�R�Κ��`�U�����UW<gD�dq|N]��<�c��6?��,`R�e��C��R�y�jל{�ݦ��do~0z��m.�v��jF �VID ? ʟ�>24:}��V��[6���[�'C���b�uǪ"U�D�Q�<qFv���6餅<=j}�O�D�2���q>z��d�1����	.�\��Ui^D�������'��")�����{p7�b��H�*%���, V�7��Ս�=�I���<��M[����y�� �&�\��}�Ue<P��Wd&��UH�����vY����ߚ�Y�҉��ˌ�K�\l�=��5u9�/�)0ln
s�6�IR���ώ�d���3��L�.�[�6��K�y�S`���e���������� ��;��L��1_ji"�z�r9�A*�׭��d�od��-�u(���(Z1-:�Q'\�1b��S��Ai�M��	��8q_]d]5�.&1H`"�{U�TX�(����c
���`o�"���u=&x�I�nń�B1������~�ŷ�&�t�	����sl���b���%�5�MI���C5�����!!��5����]�r�#�A~o�.��jD�f&l���״A�*`sXeP)ػ\
d �����K��"����Q3/��U�7M|
 /��~Fe6�=f(Wv-�8�[�e'l5���ͩ��r���^����ѿ���hAR'E��fh]��\EC<(�����d��8��Ҙ���$8�!^h*_�#��F���O_>1��E����ȑEמ�Qԥ�.$	<��Y��>~O �W�N�T6���ֿw��2�a��*���)O�*�Is%��Q�JO����
��i��4� ���#5���_|�ft�����$2t ���4F>�P��ҭ�긑�6џ��.��2�J�Y�2��ODU��	����jg�޸3���_�3�d�5u���������+U��n�$�Z�Ւ���C�>���f�S�A9�ݸ���2L/�w�=��������P�VNB��_���@�fP¸�`R�US�a��$���=����e'@��L���À�u�o.GE4�	���d|����֓�5��OJ���`��m�_ήQ����Np�_7��ٟ*SւD�`-���R��p�9�ef��}^e*l����o7~H��I����� ш� �i��P>�O����Z��E|�Y����bQb�d:�;;���q?KP4�|uF��r�&tT%�m�!̟L�8{����b��P���fvfVb��
�X�w�s7:�>����۞E2Ǜw;��?M�H��b3��3W�-3��\lf�~܇Q��0�Q9Ξ��w��G�b2����/D�hV��Y���-V���-�!���K��>��W�E3Q�q�<�ِE��X9�/��ˁ�D�D�Y0dC\�~b���;�F�.�ص�mvƍ�<]�s�ۻ�����ʘWІ�%�T���;'H,"�[<�+���E\�6CI�f[����%I�	�*,!�	m!3�A�4�#��,��"���M5����٣��b�T��MK�=p��z�TQ�Z����f����><-�{@ߟ)-\��f��j�F��烵e�����	D�&�kVH�O���:?\PȒ]�w�(ޠ],$�Mz��P*�W�(y.��k2������P�.G%�ͣ�.��Z�T%����X4�/���\x�\#lIg&h���MK�{�*
��\��D%�y��Uc��b���))�7W�]>��_8�ܒ�te%��[�����2�SĒ ���O���Z�Ŕ�r�i�����|�Jgf��-n�t.S`</z��Ŕ�B�}��lr�a�K���*��Z�SJm"�&��AʈE��_���"-�4l�( ;���X���QGy�yE�	>m{+@g�H�A:w㴨i3�8��h.���;^��8:���A�G8��	/�����ov��:F7�+��5��ۉ���@~�%_^���(G+�WO��S��Y@�߳����oӐQ"�0�+��3%�*�������[�n�TZ���P�ѕ��OY"�_Ƣ�/>anI��;sA}��U��W���n,�s���^Rv�����f�ǀEE����a�x�K�1|oj��y����T��L��Ζ�e���G�~�!г�#%^l2�&6D�����s]������S�����Y:���zգ�/�_���ò�[�S�fu8�2#����_�|`��6�{�9ޥ�/��!V~42!�>���hD��y�`)M	J�#m+J;������2~}��yv��}H>�6�������̓6`J�7L�����;1�;uݦm�v��\��C��H�ƧWb�6��T6�4{���ͳ�o���Ļ�D�C�bCo�e�J���[-*���4�Ʉ�v��b�B�B&��3g��9bL���d&�� ߕ�к�ݑk�X4�|Ʈ�e\�;�l�R&���!�v�Q����l=��k��y��Ҳ��qP��0����4�A�n�69��^��O���i#<2��`�%;c1:�V�.:� �6H�ݙҴ�;'���X��䕗'�<f�����E�/	?G�� ��c#��&
��k�`����I�R`(�; �ExN40p�����D%=\�f�o눡���0��LM}	�s%4�����W�L��!G���R}����w�\�ٹ�j8N`���A�����;�HRN?'9�Y���˒�u�w��P�{�+�N���,��cr8�8������8��J�&���`BX*�>�T���}f[~ep�O������O�y�9��&��v.!��^���3�\)H�)�3�Q��-[Ǉ8i�f1��'����\���,^�q�0�,ʼ�֋�v/-�!"�CwA�K��ޖ,�	��ey�I5��yV�ue]0�lt��B��2[�<�I���޺r����<M,�}�
�؏��T�H$ &�c�q8u��7����� �_&��]c�Q��Q<�){���=�w7}�G ^��8IO;8A!����Q_�B*�'������P�h���-�MS���|�z˭(4O��o��JS��s��ۓv1��5�3����&��.iE?V/Y�z�	�%;6�)�cG�w{��s�����7.&�him81�d��t��Q�g+��J�t��0��ާ	l�Ӗ��x�Vn���<5�h��9��lŋ,Kp��TQE�<O��\��j��@t�썞?krO|'�,`O ���H�?�;%�]��r:�uW˕�f����E�M X_�,��H��]�N`b�_��y
z���+;��Js�^��.�P�x�)Jo�>�n2^��R�h��h&̲������Fcu0v��C���g�R���G�6V��s�5e�@�pŁ`kx�u����Rv��4}� �z��Ĩ�~?ghc_:�	�ܽ~�~1@�Y�|ސ�+OK#a;;~�R��ɮ�2���d��1�rn��x.y��g���R�Fi���s��-0O*�^�i`ԝ�-�5aa�;��5r�e�%��[t;�7���9��NGW}�����y��6��n�X�4�9�kz
��*B�Y�"]��1��;�A�B���ꤕ�����)�����5g�0ؤ�2�3ڧM�p1��ݱ!�c�V�"<�I�T$�O����s�Ty�
���dT���G	|�6ЊE(:�,���V|}ϵ�2� ��X^n>�O��A�2LIӬ�� f��٘�
L#�F�� m���3����M����Iz" �hkA18"���H�|��,=�R��N����۱/ìFj)�P�fO:�{1p.i�Q1v�{^Y邱ސl��23A��ׂ�����4��2\���Ȣ�z<!����� 8Tq'y�{��R۲C�Y_��>�^e����@dC�	�{K�5����1���'���r�Y�_S���D�n8��VT�����@��%�Z�q+J'��5ci��=E�����ʊ͒�'5?�>��^��J���nh���`a\+����ȿ�m('��3��?H��}�������	ˁC��� ̜���o��]M�R��,!����`#3�����z�^'8J�A!A�z�F�3Q�wt1�y�T�]´��o0�bW�aJ�� `7 �އ�/b��#�F�m�H��A�ۦ�7�hc�ג?*OzI�E��:)1��G94�@We��i��@m��cq�K�$C3�����$-��Ԡo'v� �72MF�B$���qWN�?�ÂՉ��a����-�;T@q��s�5�qUC�U��F�O,oez�1���V ^����������j��#�#6�ؚ��+hOַ�d���D5�{�/4j��j��E[��T|���l�謮�y%_���"�3�S\A���	P�.�LE��x���� �����y���T��aI1��K��b�K�G�_#\?��ZS�(���o�.�"`>S>��$!�~���������q�nކx'*�`�Q�8���]��������V���!.P��.���G��7*E�p���0���b��T�!v���z�d�T����ΰ���y��Bn�o�IOj�T2��n{}J��Ł�v=��'ɀX�NKM�=B�f�Zҷ`y�rq�c�����&�9M���/�m2��2�b�i��3AR���.���0c�:#��[� V\`*��
3��^Y��:"�xш�g�;�>\�]�7*ȑZY,�ss6�/���(��g7�"%�ַ<!J�\�@q�[�80��Յ������wj	�Of��*�2����0�Qȉ�1J��X���էOH��lt�i9�>�ڜ�Ad�����
��G���S��NI&�"T5/��(ب�F��WJl]ɖ�B;�������>��Ԋ�'+����|�\-�;�yΜ����b9!p�b��yT,�<���l���T�˓��a�?���0���^j�<8�`�wٷ~����#
�W�uZ1��
%�lU��U�a�����H�@v���Ǟc�z�yOiྮ�m����+�ڠk�k^(,�_�=P��&����=m��$��naS��[�L�'? i"���v�b����x�W�w>K�� _MH;J���̋ZU�&�*�f�᳊x���q�/��A�.�kjm����b0�4D!�%���E�i=��V���p�&��^[0a�W�tf�B�EՎ.�8p��6(:\��q��a���Ъw�O���h_9v��u��S&`�Wϒ�eA���g� �(')d�@��<��+��gl�҇�/�[z���it%,bR��Y�-��<c<��F�����&����+���"��4�`e}4C(K�u�@�KL�G�4�z��[��v��=`���n%bЁ6���ts��-����pGN19g���5��*������M�ϛ:t�E;�Tņ-�TG=M�i��@�y�1�<a�"Vǁ�j.�!O%�bn9�U��ܴ�Ww��M���XX����0�G.�wн� �Eh��͡Cx�0w��q��)�ٕ�)Q/̣�3��W����#�'"��gV�XBW�e��0<��!5��_�jz}�?k^2���F�2%�I�Jݡ���x�Ht|RsA�Ɖ䡽18�OSͬ<����>�[9��H$rƮ��b�f��|D���