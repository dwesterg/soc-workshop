��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��T���q�Q���ڷ�~-��ShwI%��ikt�F�M7��'�V��]��w�QY.�|�~�Q�CfE�a�Lu�c���㜶ߪ�")	q�b�y�B��\v2�����5i�Z���A�?;J�h���vLwT���+��W( �S3�
)�-���G�*�
E����drP`g��j��ˏ����c���)�_	t/C`����C�3��-ʚ�X���ʟ]x5|��uZ#0�����B��*1�m�W��LpK,^��ܷ��5�����®���gv�� �M���k�ܽH�E2������*�'H=z�x���Қ��GO0QRI[�1疷5��˒��5�G&��q���5}T��[��--��W��]����(M"|���S���G,��wӃ��\$|���h� ��Q���w�Wx �Y���5$̩Σ�f���#Y���#|0�d�5��\�C��πm ]v ��h�Õ�ͦö]��ke@q5Z�m�Z8����/�'�7ȏ�����;�F�p<)�q�F�~*t$��c�/��	�� ;44c-.�1�罥�� 5mǰ�Q���s�!I�A�3S{�u����S���J�� ���{���Jw�aR�A�l>�.f��;�u����խr{F���D�#/)�i\���)����70�E��dڪ7�SJ�RVF+��xt`ٹ��[Ԩ��c�Ы�,9C�� Z�ή���e]>�m��(w@��O�Q�`*e�8��Ш)�����!�^�k*�m�TBD�W��v4��^��K�}iA`?֑n:�3���������&;�5�Ny0<n��	��n��!��N�a��5�P���њ��d�*0��D\/T�`K}�
�k��M�!s=;�g�Vo=R�����)2�⟓j���Y�n�x9jWA��=j��N�.�"u��i%M�9.�A͂x�ӎ������ɛ�m�Z��g�^
k�E/�:��|����gM7/�Wb�D��͆�圓��u������!L����f�j�K�v��3T2_�F��i�`2
Cn:�u���{�!�p����Vx�z��R��0b�}♡��q���3�	���	�N���@�A/����W��˙�˯	<ıU>����=��� 1Y�ֻ��oΩ��/��y_:7���= i�2�L���+S}(�T+�oS]<����v45T�Y[���\y������� ������ل:�J������Wl������ 5�Ce��ck���z��C��k�Lp���k������ĳ�3�b@XZ�8��g�o��K���"��s�$ŏ����!�G��Ս���R�n�c�(
��Z�Nʤgq��c\��j��[�]sOB�bu��y�@�11ba.2!ް>D36S����5�w��Xi˶6�Jx��+�U��0�.������&E7R CϖLÂ���_�Kٌb�uN�	���"p�4��	�e˵�i����pE�B���םd�ʠ��ѿ"#0
ܼ	��u�A閆�qa[t"G]�2���Wv� 1L3��F�p�^1lM�z���h'��ճ��-�N���Z�o�)��α��v��Q
��j�=+za�,� �X��D��s+�W����u�Lzn�@p�A�P��(ޡ���	�=Gw��Y���k��u��!L\S�)]��M!a����y��]�@Z �dLO�̨�,�]+���GJ�H���-�O������@:�1]���������Wm%��3�b��hc��%1>��͎��E/4FLI�ƩHu"^t�~)�	v@>�[��4�Y��5�n<q]��=�p���֯ȩ�G�w��A���A�~�?��O�|	�e��J(u,ji�~�f[Rb���@�'/��0�,Y��t�K!��B�"��$G���H��GX[��s!�KV��0�#��������)G�ްS��D�}S�8$��h�h[����jb��k�����O���AV����_�0_�{�kׄs��σGԊ�s����m���|��U&HW��e�~�)�D�.����2�#�zق�D�6�K5�	Aڜ�2�}qe~�5��V��L5�eL) ������Kc��6+�'�J�!g����Rz�ݔ|��Za�5A,�9�X5�	�*��^ja�{��X�U ��q]�7��b}�͹�ܺ�|��JBP��	{0����X�ܸR���P\�Wq��*� i��G�������:�+�nYtȜ'4���;�R�VZW��%���=\������aA�q�뮰��&�}!\���ֲ�����*V�|��tׂx�Ho�v�0�&����逮��^��8��D��XZ
@�y��Ď�۪��gr�$�[�������?
VS�v6��}��i��d<�H>I^'TJ�^�~zD	��]P�L� '�efu��M>�r�x��m;���s�iE�<O�B�.B�,��q~���H�D�&=��.�3��&9�\3i'��t�旾BR@m����NN2�=��<ZAO�$��/,��B�P�4�ItL�D����Mδdm�S���Z�0���Bw.Wꨰ���5����uǝt����v|�9U���� �a���&���
L-��,.�>��>�޲h���hS���lĆW�١��"��8f�P+�S�|��6��l8]�Ƞ�T1(�h�>4ǆ�9e�c�����<Y(A���=3�W$,[E���3���E��e{�}��B�4Z,
��/ůy�}�2��)	�Ev��cQ�	�д.�F\�5�.I�Q��I��eq@��S�uLY����8i[��S��^����!�;C+O�.KNZ�E���cm�	;<G������,`��]-}��ۭZ�����8%�7%_3;��ay`W96��
��?i��2r\��*��L��������iG�K�N�+A�/{��@���t054?쯏�uqQSrÜ\F�V�hK�����xH�~B"�T4�AE-/
�/,��8ED�!����~ܾ[xC[ߋDLj�����O0	 �͎e�!�M��-C`A��?�7"��[x���Xߚl��4��0�;Ƒ�A�J��2F�W�*l���U�ٽ�X�>�KXlɺp
���p�|���R�LZO^O�m�8��"N!Ľ║F�������O��G;D��B��6T(˵0������Ig9.�v�^q�"^ϫ�Ɉ�/��gs맖��w��&���߉�"�q�4@� m�!���6�EI��|�q�8�a^z��¼52S҇��^U>�����lE�K��}$	A*�D�>i��8�B�Q�Gm��x�T}i�ұ�`�f�R�ْ�RVp�5k��[��$�)���k�L?�����q�|���qh�7W� �'�ʬ����$�葔����V�wV�* T��F���y"ڟʑ����s
QZɿ��0�����&?üjGE���j�N�B5*K'�y)A�*��iG%����	��+�o�!q��rajl�r����?=���@V0��Ĩ��a��R6(˩Y	7����o>�(]"8�c�\����	�JH&��Ix�����Zæ�>.�[�4Q2�\?&���i; �K]9�s�a�Z����>ܘK	��o<�	��9� ��q+/�Y]�+? ���$�!4E��y�{:�;o�H\և �	�P7I$+I����`�Pf�+D\��?Lx'J�t�n�;�u��+�=DH�F�W�p�|�R+�{b��E���h�ǢU��U]j��I_��7�G\t[p�2=-1�O�h���b5��^����d�`T�P���R�ނA�S�#F��&)_!g^�3NR�	a�(�^�R�,4	�>�g�������1$?Ng(].%c JA���r!n���y�������P�Y�"�l�8�z9�_�'2Өډj�4{���\(y�hUC�*��59.g�`�@������<wQ?"ρ��Q�X�ʐ�������h\�0��L�.F����S�ܾ,r�7���<~r3� ��]vNn�����#P��e�,w�;'��#W+kմ�1�-�WM_P��@*{��h.ỻʦ�<�K�`ғJ�Q��3y���c�����唹�|�,4-+��}_��?y�%����V�~ ����?���>�W%�܌x e��)���T&�����Ľ'`M���]��U�qF��Fߺ[$嵮���n���3�X~bo�΢�+�9��Xг��$����u;�a�k�I���!��S|��5�fXW"��A/̆{\K�Y=�-=��P^a#����8���i4x�"��I�����ӓA����و�J�~Z�O�ߍj
sf�`��׭c�4]ǈ�� {�B#zXІ! ����ᗬ%��K�ZIO�Q���$J�*��a�%��C��7��]�E��k����4�N;�^
W��v=/����hQ�*1�l����5�>�,ގ�c��)�@��i�h���Pؔ�|X�p�%��h�9� ��b��x�u`�VGfK����HJ�?��hǁY8�:��]�<�!�ŉ4ik����H���˯[m7��D4r�������Iƚ���q��Cs֭8��l���)(�fn����
�<�jxt0%�,,�qޜ��)���eSп~B�-����@*>�V�kg
��PO�A�b\lDX�lm�S��s��B̗M��F�%���E:ٖ��aT
ʈ��Y9�tҗ}9ߔ����U��Z��Ĝ����R�H��5l�S�*x� ��(s>�9A���M�>)-�����_�b�?��_䋭t|� t�U[�������s;����(��/�G�j��Y�/S�0o�CG�?S=QxI�<-���K���n��հ�}<���e��$�m�=��s��K Ҵ�mF0�|�V��yp��{b�Al�F$+�X�������60������&�Na����S*�l�Q�.2�ν
�s�g�7|�O��*������FiX��6r��Y�>���ξ^�e,���(ڀ��7��ps���r��C�Vn%G�,�9�2|BA-���jG�Z~���ݯ�_��<�i��@�bUV�&�p���_�5M$��ֻ���6���ؑ` �z;c8�I/E;A&��1����cKpj�.4���1R-$���`ʢ��R�������.���8��������aV����98�?P� ̬�i���0

��0�PH ��q,��cP�p�{g�9�,��u�����}6
��ġ�����+�K	]�>.�3���`�q;�Rnj�1^����bH5��N_!L>AC7����[&�g?������a�0��2�
'��n-��.��g�6@�{2�pH���r��?z;�8��?ۆ�녶�l�v�����۩ɔ�Nqa}�z�$2�bh���0l�A\�J�%�{���ɢ"�'��>�j�X�T��|�����Ɖ��Nl��oR�s�/���F%���8��P�㇖��I���T�`���=f���y.G!gj8���p�2t`�ڒ�}����X_���Ȉ�YW��7tr�E�xK쨠2�=�[�x�1���ܓ+�7h�����2���:�^t?p�oզ�-��w�"�o�������]�"�lWs����u��H�H�1 ze��o6����b��џ�*��D��xɚ99t?p\�j����F��GmS)R���]�?���k/�o����u�I0����
��!|Ŭ��ET��-YV��6����<�j�W2��|zuK��[TF�ɎP#���`&4�L����Q-�8�7�M�0mt���t�(<�z�yY�L�"n� yECD�HN
���󞲸����*��C��
򉧖T/�J�Yŗ^��F.��R6�P�p��t��d���9�_FavW�}*=�Dc�j6�J�O9Qw?Y+�L̲w��l?�ͦ�\;���}:-t:��=Ux�K�����oC��ũ-��U͟�@�I?�?P�_�O/�p�l��vS��n�2�>�8���۪���?�ʐ�p>���F���$�xQ��������tj��>q�5?�8��bx��	c��G	��v� N�P=`j졇ɣ&N�TĞ@�_*�ea�����V���YsLx��p(���<#��|ʇ�_���8��&�^���5LZк�|J�bb�Av)̔-b��z#[���y6�j���Ԅޤ����P���K�G��d7�ld�etÔzt����ۥ�:�2_%Ԗ�/x����m�%(�d+��x�"B$����:�|Ǖ�}�	/ؤi�|�q��a:�#Y�CD�e�����]���p�O�:DOM�`���S" v��I��pi�<�4M_a-�&�zz��4M���-u�N֫�E�-����=o�y�K���L7���0ϯ �C$��N�/����s�f�@��w�6�}{�����wH�F*=��ȣ4r��E&$N�@�\ë0B�,��!��B3��{�����Q��Z�p��=�7�Kv����bʇ�|�������GJm�	��C���U��߹����a������oϴ�ĵ�!�[ ��H$��.ǽ������u=� '(dxR�O7�_fv>���Ͷ:��;cd�z���Y�P���pr�Hs�=lYH᮲��a3�2(v�!�K��<���g���ʖҖ����0�������u���� 9Ui���?k|��1(]�>c['K1B��k������٧�:<���݃��֜�����Z0�.j��}-
.����m�`[s��K2�8�t����'�" j�n�D�pC�oJ��p�WR6���AϽ C� O�9�~�&McG��6R�?���6=�5L=>9��Np���V']�KP@ԈO��}৵�)�k/V�2�.��_�8�ys]��?���j���Z��`蚦�:t��.�b#�����Bܓ%�/"D#� >����`�3�	+Sk�{/�֝^q�!���߃�%�--t��Q�5u�/��¬�g�o�M��c ݝl�ԯ"�(A�ӣ{���RL!��c(ZE�Y��hrc1�L�f�#��=v ��ԕ����)3B�2�.��8���CS��	�2z�t ཀ����+̿i�����dt�!#�dL��C�e�?��^�3���jӚ6������޸V�y'�e;a�N���Aq�ZSu��rx�ޑJg�~�WJ�Tuc��O��
)�æ���
m��������	�SMJ"]���U�m���Cͻ���: RC ��f��ܪaʾ��.����9�������w.���V#L7y^�"4]� S�M�wX�q(�����'	�N���P�/��]�8�~��m�e�l ��E�腴R
�OY5�j��u��Pz�]Nr�VS��gNX޾��a�w�U��9�f�E�F�Tj���*M�g)T�ޤ�2�!��xnZ:�����Y�K	��x���Q���?��霩�7|<�E�C�৫)�S�y�H���gL/��N��[>h��R��O�t�m�:g��2W=�(�����45�9TP�~�g����4ɖ{�������"�uG��JX!�fOAj��Vz�P�Ș�q>tA���5�wu�3R�`֒�&�l�����h.�/qh��+;�4��nj��N�j] �E�h�dZl��l�1�'��M�-�'꟒��%Z�
A6)�u<���N��S�o��.�A�?��s�&1v��~U�����7q3�κ2�B&u��5�T��yX��)���$�C�7F������(�`��{�<��Wþ�y�S��by�*�����1�7�y�x�Ӛ�9���E4��1��!f�J���Y�ڥ��6�WN5�Ӄ�F�F�,y����W\�ta��	}�u�R�� ��k��Y�C�[���V�c^���v�y�>�h�L����!p��P%�G=�=�9*� 0&U�aI�����	擛2��NP�հ3��kxS'�)��HȇUn������)�Y�$�� n!`a�	���U2n�;#?����s��^�k=[��w�i;ƌ,1�������:�qQ�9d��m��:mb�EV^K�3dTC�33����
Y�Xn��]J��C�9e$�˃�l�dݞ��+��� HSD���e R��X�M`�s��s��,�>+n�48��S���8�ٮg��h!!"p�Œ	8�^�K�h�90�:8TQIsg�`,��L�5]����X�	x�d8�4��qԳ�GBC��V"�'��5D�ۻ���@-x?�&pSo{kw`ؗp(J����A���ӲQ��_䙄��o����w�U4���c;�c�8�7�YR�S����{;-����O��+e�n�����>	5�$Ҁ^�l�@����|����`&��z��npd�S�<g�C�+�S�x����Ƨ�A�z�W�bb�	�����A�h���H�Q��^�8���*�ov;s��z���F��Wb�#=�.O�;��0)�2}{w��{�H!���ϲ���ǅ���	-c��b���4HY�~i�胳4~GݔF�)���`�ey��*,��:'��!��\>c��fG�ӛ������'~b�Ck����J�63�3"�=��4W�r�i��p�K��!��8n�Y��*�13�=�F���0<>�����B�^�����#Y��������]D���a<�7k��ș�T�� Խ�hŵ�p.9Z'}A2�<����L(��L��n�U��/<xh=��i��5�B�����G�z���4�H �2˾�ޕe2�<iiL��s�N�T����o"2Y���Q�^j+Ó�V��y����j��������?��ڸ#]�I�ͺ��yC�~�H�Ϛ��.����� ��RV��NA@�bMC�!s'��p(P�de��Zu�\�t�KY�X7մ���Lh���5
��J��p��W�zG��=��gԭD�=���#\v�r�T�-�ТxȰ��/�I(�����Z��֗eH�7� U�RM]Wl�)�v�Z�(3[G�������?#���*M*XP=�9e��|�vO��^=��^������|5����^���-�.XJ�s�#1'�oA�i�9qeL7W������HP�f{ey���\W^�^��Ǧ> �J���7�8$�'�Cc!��2	UGG�Bw����6[k�+.��y
;�_��ǥ�˸b���Z��ț��j�Y�7�o��^G��h����֋�6jpq ���������F��x�'�����޻���
�.'$����q~�M�����zR�������<{G@�YH���a<��E��W,�| �#��4��R��\*���ǅ����)�;�,�u?=:b ��,�����7���A�o=��Ϗ;��">B��]Q��س��,�ADgj���u��1�p��wA6Q-�,P��l_���t�Sdﴲ�Q�p>i�#4#���4��'���<~�3����4k�@�3�c�S&`37��&�&ğ���|h�= Td��Ʒ>ĵ�E���g��kD�P_I����f��"<l����6���,U�K`�L�"u�:P�ɐ#��H�P�pK���"�$�h�M��%�^52���1�����B���8<��**���>"��;ɫ�m������~�Ώ�]�x2D� м́{#�	c
g��5��a�
*��� ��n#C��`�n`�3z�r���-曇ja'��D ��ƕ��*�KM( ���
ܜ��a�uli��4(��G9\ ��M��/��e� �c��$	]�G힚�C�򳏤��+0`m�|L��g[�zC\���F�uOᙷXg����0�:S-�w�R��Y���K_����E��2�"��=��+��;�������vȗ�>GBg�ƴ�af-� W�ï��ʗ>ʕ۔��=���>yt�>V-m}{J%?��S#˒*�$����-��7������Գz������GJ�:����"�����*���Q�@QEZ�e>�@1����޴������)��$=�܂ߚ��A�+�^�ŕ&��AL�3��۝O�=%o~�mLͰf�1n��``���x݆# j�'چ9.�l�{�]���A�Z��i/�08�w�$ұ_�XEI��bװ�a�������R����!MRpI����Ц�?x�Q#	J=���v"xU���%�6��&�ڤ�Ա8�=3M#�QdVf�!���fM3e�F�H�G0L���s���!|ʖt3_ 0��|��~�M��z�O$rA���QJ���tw0�U aX�W�S���dJ� \Q��ûW��|N1��.��M}���9l�)�휪�/AƹVy'�(o���$�3�!�|Ļ n(�4Ɗ$F׋����@�XW_nR3T�Ŷ�n���W��V��e��'�xX��FƇ`�n��Č������0D(����}�Z^(
��Y%��tR�i�#��#�Љ~��>;?�'G���'"+vj�ꆾ��֐�!�����c�(�@Y�~"NA��8��̸w ��I���4oE�˹��� ����0�,�: