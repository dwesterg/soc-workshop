��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���KN�𢽟1k/�@8���Ec�����S]�Q{E�J�nc�?/</��?J�5���{��$�7�m��+}F%��yE�5���!�K�G>�tE�\�q��]bG��:JV	�-D��Cz��,��l�1�2���0�(h���t����Cv�r�h�S4X)%��2����(=b#D%�D:�W;�x���;u��-���k9�C�l��\g�1(CG��7p�)n�a-mZ�U1�����fmyy�>�	Ys�s����(�ʉ.ä\jP^pX^5��G��n[j�f]
�n[�=�C��ߘ���Ҋ	��)s�����n�ح~cR���:�7��|Vw&�op�p�%����JI��V�m ��uT��|/�ii�u����$9�wz)�W��3ϯ��/ȁc��kcuI���eGS<�u��C��3��ګY_NFQ��.~�֧�O%dɀtp�`1�Ŷ6^$�nI�@d����-�
�֓߼w_,�"�œ1�ԛU��/nK�/��L����Fn��biu��8�\J��a.ȵ�p-\I0�O�Y�o��ץ��]HN�s��-�e��I�TR����]�-�����A^�,F;q�� ��NtE|�����$�,c���f��d3Tc$OT�F�=NЮc���#��5�RSN^��z\I��W��s����,b��APǈ� ��QvӪˉH��-�t�k�6Jb�@ΑF^����Q�c�a�ب�Imā�1o��>͇n�[�4����	�#�S��àJb�	ny��fX��LNH�u��hZ��E��Ǿ2qHW���6�k�((�c��ˇ4䵘ض���;�3��mB��̅�xN�~s��v����n«�8x �Ǽc1}��-�/�7��q��ȓ��ab�Ҹ!<�K��>m��s�]��ɞ�cjDcʹ#S��5 *Z0�3�ܠ]p�ms)P�z�ڑi
��$nx�Z�6���Oq��Z5Z�il���Ϋ�[��Z���	��s=Y��+�eBP>��n��߳�Vj��3�pb�؅��p}q��nX"�]�g+�#u������>ߤj�E�+s�)'��W���gi�ؾ�IRd+�k��x�#�Hߣ�S�+�v��;�+*ڜ@I�r����E.���{��$�n|-��$�*b�$S��J�����ݶV��E���$��%7��B>����I�ݔ��'��S2�OS��ҫ���8��'�O1�H��9�Y~,�|g"���W�Y�8�r���
���g!n����0�ǏG$���{��xF�RÏ���P1���D�Oy�h~L��9�'��,��Z
�/Ba+ma�U�t�<���*�;�C	�\Z�b�����D�pܬFu2~ABU�Z�P)1��̳��\��'�)�n��p��X'wh7 ���i� G6u]`�$;�:I������,�ƳzwF5��Ղ�zZ�d���������u�2����CFӡ�c��M�#�U5fH�Z��dACg
�e@�X���!�
ߑ�$�����z� �<�
k�S>��!=��c�j�B>�+��� k��+���R����R� ���|ɦ������tS� :h|��Zc$kT=�<nP%������˟l_��1����B��+O.P�a3���LV>�>, .���X '�Mh1�3�����<(>�eֺ<0�H�#v^��;����%c��$��'���n��gh�?��j??�W~O���n�z9�N12��q�&�dxc�����F&��tbr^&ۄ���s?�a��@�6'�؁�"qO�(��sUy���\4۫�B��o3޸K��BsXښ��/���n��D��e�y�)
9ގ�p���o?5�{��ZNk�i�#mq�7|bp.:�`k��?�vC�j����!.�ÒB��{Ͼ&�ev�u�	����ͽ��Io�U��G;�$�v\s�!�s�s������[S�����3ηv2dj'�tJ��kĺ?h	w6͋pg6���IP��#�ԅ`�b^��Gz����%�Y�G8�jD#�9y��(K]�������'T���3C �3QYP��Y؛���r'��|FZ�G��+�[/P{�6�i2��r>-��;��
% 	F�o<��� W �c�O�/�N~T�t唘�t���� �)���sIr�qY偉[ڸ�� Qt���`8ef>�r��2�ۑ��U�����"@��*��^aӋTC�����7B���$��"fl�|���H�h�>��Z+t�1��Q�0��f�CS���6��S�;��f����-B�o�`��������SZ���%,5\���;�̝M&Fp� ;�+@b�u�)X�v�[E&*� ��|M�`�&�߼}��'�E�N#��z9��}���A�sh�gXg\��!�ڽ�1�)ϓ�Y3Z#����t��H���f�u�����p���<�3*��bK)|�.*���^n�M�B!|]	� щ�c �d.�H��_~q��~�����FA�𔀄_��$MϠ�~8Q���첦����k�p�[��g]��}�����Q�Yl�@(S��/}2 �CU;� �6��a�ѹ�{H�Tn��Hg���6S���H�-F�;Cj�Z[x�������S5��=�HI��O��M�l��;i���-ɫ�(�K�uvx&��c��.�ʦp�H�%�a��w+b�O�
��G3��R9�x�)%�4Rt����#���i����!�s���� m2��E��C�Z"),�L5Y"�U�J�(l8s'����s��i�݅��I�|����A| �Q�:`�R�Y���V4�h�:	�%P+����l�����ʯ��3��E������;SQ ^%�����.����T�$�Ȫ9�j�'}M�Hā��Vtis�!Jl����$���LbuB m�X^^��ח�H�@�Q�WK<���ܗ��(JJ�m��m	dV!-~O����w^y�i��uP�31�H?5qR}jz���w=1]D�t�\�2�p����o.��/�� �������D} ����p#��U�"�j�uqd_'lR���'tqeU(8z.yg�I!U��*�IO�*�GL{os��څ�y� Ӌ$��������C��B�V�ϑ���-���4�������l���b� � W�j�րM���5&��5{S��ib�y�X�$��#��ũ��#%��^E�讳�~ð��-��9 7ͬ�:��E����3?$v��B3��#m(����C�����yh �i���l�Ψ��x�)V ��� ��d  :g�1H��r��K��6�I��᡻27Z���2F��j+H[h}Y�Xŭ��9)/g�|u��8#LT�H{r��^�j�!ꨇ�
��w1q�#/��C�t��O�<�$�,֎�/M]j�I�������'���x ��(Gi:{�k�Q��	�By`w��� B�@�p�]`T�o��E�̗��2Um��I�&0�����҅�6E 1���DW���EѮ���d Ab@�Z<�*�?JP�W�j�Hs�����D�_��f8+i��9��beMi,����9M 7�o;�!�zf_�x��������Zl<��x��)��$���E��N@kDO�	�hX�0î9�O�)��KH*þ�1}�,F��7K�27]o[C��QO9Wy8�G�&���d��$T����D��(����*��4�8\�����B�XH������D� y�0V��'���B;-����sU��nM�>��OYn�dZ_Aɿ:���2tS Zۊ㇡y'?��'�Á�[���',5��.[ "Ga]��d�'CĦb��)�&��\�$�JZ<S`�d��5^y�$�G��2��K�;:�� ���=�����p��tu��̜I>}h�P�����-4Pz��|�����5ێ���V�db?.�?s�'��:��_����t��N�ă��yt����q�i�E��l�s@�P�V��h��k˓o��'��HQ1�N�a��'NͼPƺ�Be�iLDz�|:��T]w�M�H�֖K�ypy����{�U��ו�M��0|��f���ڻg�B��9OI\'��D����u*w��~�P�~:�����L�;< ���7��]baMC��z^��Ϙ�{MÄ����ژ8�&S��đ�o�/���F��&ow��4lS�?�=�x0�s"t��,s�'*}P�}����C2SP�?��pz;�En���{+��ȎV��|d��E3�~"?����H=���:��	ޒm��+�k%`p5;���z�은~���g�y^�I�B��&P��۽zb��BسD�j~�(���xz�\E�&r���խ$��S�$�[r�V�M��D����)���}�G'S^�V�.VX�X�d��O���>\���X�O����,j�-(���}b�����&���5�z��qL�R�,%L��.���Y&��x>F�w��͚�K�j�e�tS;7����H��:i�I��_怒K�d`g'�C#�����G<�ɓ�g��j�2b��zqV���R��2op�I�b/�9o��lgN���,������E�`v3Yd�~'���^hZ��@H;��&�"�Z{�Y�BgR5�bV��w��BbT�i���||�Z'�/�a��Qd$�