��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�BdC���ޖ���'��aDEt3��a,�ى��!1 �d:{A�D��=�CPb��E��ق�o�ֳ�}��=��aӮvS�� j���힨t^4*�P �VPc�0��̤UV�P��aK�2�k�6.r��[t ������[c�\�k���H��!T�3�᷽�^� L���b]?���%�JbM��-_�M�g��r�`��̏�>r⢊�ܜ*.�v�Qn �^#��b6u޺������&a�J3Kp��5�G2ߘ�]\�se�A݄g�yU�ԝ���&�NXe�ǧ �T8a_K�e_f�݊�w�/����6Dl�����Bx{��?T����	AI(Qh�;y�c�d�]��.��&�	�ђ}�[{Z�$��e�C�yJˁ��|�$��u
y�	�sm[�d8�%�
Rj�r]�P���L�a�7w�ذ�A�$I?��b!�0���i\&⟜�ȔU�Vr�ϣ07l�(w!�ڛIs�5>���9?� �?�,h�ə^�W���g���`	�Xo��%M�׏�Ez����m!�nVv޲��6<��>6�E j��PsY^��-)��|�9��\16�Kwj��y|O7L����ͽ���T�@ro�;������?	G���\8[����K=�T:Ḧ�P\r���ugݧw���<>�x@�3`PeZBTf��
ݜ���<�F�"��7< ƴ(e��E[�vG�4�E ��7$v6E�u5����v�E��*Rm�F�O�[��=q���%�?s e8/������Wύ���$7M��0���z���O��}%�	wN̊	/������#r3<���ߠ�ޠf�_&&9�� ��:FCW�~/�k;��Cl��-4�7x��!��(�ɭ���l�%`� ��Y����7������^G����Q��Zd��O��pO�?��z�(�R'�a��L7#� �x �20\_[4c��$I��_Ӓ�'	~8C޺����5{Rn�Ǽ6*��mx��zhZ���"֒ض,�/�(^,������!��T�D�(>�Ʊ�zl����r���d������[�l���a"��y"X�
X�EE�mE���HYv�%?�ȮsGD�R�a��~�C���/��ޖW�@vĒj��lI����L:�|���Nj�~�8`G��V2��B~�j�-\�}Ս�i3���~����ԋ/�XY�9�q���쾋@�B(c_����K�;+���Q�\��24��#d��\�#�Bc����3�HMsF+~G�"ov�^8u��W�1��u�ے:���w@nk�W%)�X��G��>Ģ:�M�Y]��E���mTп3�}�_8��D�i0D}�"�?|�D�a�r�{��Qg������\}�����>�P��� �j�f�����pq� ���(�Z7�d<>}�܇7�&2���9tR��4RZ���_��I�o�n� �w^q�'Q`��ݤP�[�������L�*'�y|�Z��6��Y)��RA..l�&c�Ty�����L��(|%B�!?��-mE�f	|:4��a�\�_{�Ck��{��FyD~ϡx�t�T�j^"�t�{���C⎓�<��{h�:���Q6PE�ېf�����ne��Oν�c61v��r�.�������?�a����Њ�����Ù�Zq�a����*�E���1m�bWa];�Z��e@�9�����K4\�� 7��q���bAN�k'�'ƕ�P�2<��h_f�6S��W$$�[��
��>����}�緻�6���.8�=�Vm�Kd�O�I�^��$����K���sn�w ő�mK
�Ǉ���$����:�n�FF�I/��z%���\O{3J����ťG���^��S]`sc/��2Q�P� �Q=ulw�a�Uټ���9�+�,_���&\�@� ��,����%H�G�>7���Ӆ�5�z:k OC�������61B�8�&�e��,�g��H��q-W�j�`��@d	LXqST�h�5�ŉ3x��^����?;7���@Mj-�y��Jģ��Ě�X����g�	S����,��Hv��,�jLu)�U�W ���o��3������l�i
#�e�X�5Ù���@y�~�֘sF����ճA�K�|��7-���q��%����%�����#J��j�y:$OAII�m��O*1W��`}�]����[$�q�k<5���v��&�Y�m�$�i����*K�@w�D�(@����&�K�R@�U �-���$�7�:��D/Z����|��ցX�AFLf?�G7?���ǰ�I�T56��J7�h�V��n�J�m�tzr5*��n/{�x�8H5+�����6 �i=z\�x6�m���9�5��"�c�6EOA|0������|��0�/���[��[����`w?|���"��p
=���j�aeW�ö����l�&L��/b�o�J�z�y<��Pt�I���<Ha�RW�2(��M�2)�Q�s�ǹC�8��h�C�~��A��:�U�>{�RCz�|=�42�b���J�9l�=�}�F!���xg�����FZǍ���3h{�C�.j�{�7���g��HR�qt��T��_`E���K���̀) ����/��O�yƬw��s�m�m���
Y�NqDĥ��L���3�Z���vc�it�S�Ш]cR��	�)QP��u|��Sa(�b��Z=����ғ����T]^\����6$��/�,hЙ�6vP�ߡ�>�籄9�:	�5�"@��`�:�[�>�
>�b��հ��99�,iDFu驏΋G2���ߒ�Z4h�Z��jsv�J�eo��5�Au���� �7��ǁ�<�^�t��2h�`ꆂ���F��%3B����c
u1پ��k��C��5?^�����F�#�`kw-o����Ao��Ǟ@����Ъ�*��H�8�k)��kSCء[�k��=t�q����\?�t�1_����B���#�E)5:��Was�����j�S�O�����3�{�kS�b,�F�J�J��S�(r��c�~p�=Qu�.] ��v�C�i�hH�ϊ���!{lu�h���4�L�aK/�� ���\(\LeĹVS�E��ாB����b����JK4��8):$SQ��OFv5xz��Ļ�Huk��	�\L��t��Y���s�˸��D���D�;���W��a�IԞʣ��I��ఐc�H�9�ܓ2��+��w�B���g�z���=������'��]�_(��:�<��j�[ͱ|��	��XyXNܬq�¨�Z�JǽS�e�,�����	��.��.��V��`�*���T�c��k�g� Q����n�N��RI� � D�#hd�Z* ���Y[L�J�%�ą��
��DY�8Ӯ@@����"ɒ��d>?�ZS$����z�yFD�����}�XWBn6��O]`�!<��?X��٘����klg˓k��Z[g�.��������:$����Ti��ث{G����/�7=��b�n�Tȫ�B� �9gy#����fIZ��	�0<^`��AZiݭ Z�Y�sJ���ؓ�V/�0� ��T�/���}`�oe��T��x*4R:X�*o�.0�Bn���E��I^�\�h�V�>�W��t�d��\���Yꪦ����0�{�������]p����G�9�8��8'��68�5�a����w�w��_w�'�S�����v��A ��)��+�Xs�8�<��\�V��t0�u��bܗ[o�ղC����-RU}%D(P���U��w�B�����NR�^H�mE�<24���id�I�[�D��Y ���0�۝��,�A�w(�hk7��7V?�h�}���Mo����X.#��v���+F0�_�p���ۉ�FЅ���jq�^��|J)PI�	Q�/K2a#
�5#���xD�V��Mī]�k�����Q]��`!�}���
��%K�h�ic�88��L��EO&r�<+"u��⺁F�42�),��M3��[��В��Ҵi�7@���2��
�#��7W��]KJ���@˼ΐ��7ֽWq38�����Q+u��8���
@H��ᜥ�="P��|9)[�΋-I.�O)�h_Y�7�Eu��@�j��/J!�&��,YB���\<gS:<���A��s�in����e��66�ֈV|��*MgaW��������� ��A�[AU^yP��� `��o��B�;0�#1A4H{�����{�`T	H�.�eTT�;1!k4m����lǶ#����7n��=éT�O�S�-��v�Ê}x<7^�a���X�	'���W�����B���?��J?i\8����-e�˴$S�Wl�!�[C;��v1`���<���k �<��H�"ƍ�<3e���O_ٹ��X�O�S�F��~�󩤨���s�^)�a�MY��S`��#?>�]ÿ�oR�c�kn���v�'�e�M<�|/l�ѧ���S��E�3nO�7Ҩ������Hj8_W��z>�*����k�."plmz�o�8���~=�Wd�K�w��J��%�Z�Y�㒾BS�x�� 3۪5[b�����]Si�U���	j�O��ӥ@�:���s	�<�,��y@H���n��n_��}ߨe��8�Ve��!{긛u���68��4�������q���5���KX��aJ�@���O���]tX�3?��>tV��
-��Jr�(��,$�I`��I�B<��h�W����3	�M��߉R�H�n��|�O1��-F�����փ��d�8�y��W��\�T��nU:F�� ��[��B�7��
��>�2ek��4z�5�K�U���Y�qCm(�SȔu��^�	]-=���Q��X�s[n_])`��d�װ#,�v�2W�|�Ѓ�M��!���:5St������	#�j�Q.�o�� �:�5t�/���=��{����a����&'�,� 3�&�E���+�fW�-��ި���|Xu�����2J#E"L�.��LPzg�:�<�#.ȁ�Di|q��q��$M��dT��c$3��l�t�T��c�:EO`gn^�f̎��,�.K�5��g�X�R�p����/�\؊Z+��7�)���k��{m�?������C_�<a�Ռ�-�-)�C��w�v剪���um��~�/_Li� ������:�C=�X|ys��I�pO-K�ɹX�|���x�ZN���*���F���7'7�dn2�#H�V|H��Tߗ%Nj���vp��S�s�h�k�{j�f�V��k�J 2
������
���xA�oL�DY& ^�[��> �}\=yX�/��W7�-�L��4��.�8��Qe�='���֏�4ȋ31+��t	�������$�f���!�v�;T��:���b)������-.4��eHA7mEl̩��E�"|zZ�J� �%e'+�q���I��s��YaH����s�%����xݒ�)L�/�<}�z�|��mH��~n��D@���g����؄�u�J)�S��u�.|w��2=��3zNƁ �[����{PC���Cŉ`�kݲ�L�L���/��.&.)�L6������p#��>��p��i���w��|��.*{b�Ƙ��"�E7ı��gg�ND3"�W����.g�p�,���1;_ig�_�μ�d����'���\�����v3/��v��#|
<�}<
ӓ�^4�D��R�fg�H��_��A��GB����G4,+x�vq����tڏT���%9D����
U���ƊJ��>�	��c�����x�'�;ia���O�/H���ʧ�H���v�N�q֕��`&Ko$E��fQLO�+\j�F�p4&�&+��_��A+�����s��$�ԦK��&�>��<m���"�JzG�c��Xb�-V�3O����W�=�M��e	���a|���kc��wo��W����k�>�q���Ḵ3�%�wǻwnbݣ�)��R�(��\)͙�-�t�Q\3�O�8����(��3d�fL�r�J{�:�������ƶď͋@�4��5�R��0@ձOl�����W��A�������C�����m&�>�vv(Ж]ݒ�Y�ہ������b�2#t�d��ս���w�*r�s:�ױ{�K@%�aV��yf�Jg��>� �qw���R;�sc�Y4� ��E��d3�:1���'�3�"�&|���#�'�c�Y4wCq�~���_�0�Q��i�.Tq�RAΩ��U �ޫ>C��Q���!w���_���t*)��[�S3:#>��-q�m���w�P�z������z�p�n,0��:��&2V�7o�@
L�vK�ٟ��b�;(Ya�P��ɴw*��=6�;-3���j��u	���@��+���Jv��$zJ�WG-+3Q �!
2|�>n7� �R��)I≊̞�=q���2j��?q<��w�ӘÅ�)�����+���0�����
j�ny�f�\���zve
G?�y�r�;�7�@H���D}}Z�#��5QXy"�u"����q���Vo4�9�eበۢ��;����>E,ܔ[&a&c��K��̮bC���q�^b��]�-ҢO�KQo�km潜
9Q����~����QI�Ƀ��+�Ir�XK��;ҥ5ѩߒ?\�B��� �[Z^pM%���!L���-�s�"Z���V��]��Na1���ȵ�D���Zେli��<FM�LҰ��O�����ŲZsq�!�����8�%�iNI�!�z4 +^��}�}�7�y=���p�����'�~Z�� ���kh%����_}
0{�1���G!c�YD?XY�nC�Y�W�Ųg�s�R)v^����r�z��h���ʃ�¬�����id!�����:��2�#�g&O�^��ePuZ+U�g��q�:3z2Zn���D��$�X������4���
vm��KZ�<&�٩��l��d��#�y��%��W���Q^�
�`�Gf����t0��cЕ����u;��L/�Kl�Rں�Zv���̨�������W9;y`4�\}�*��Z��g�ʾ�I<�
8ﯓHG�g�e������f��Y8V/��_����g�W��.J�QzX��=�ݘ2�w���j����g����\�[*C�eʿ%,{�]�#0(w�%���^:�����4�����G�=��Ӕ�TNp��������4�@�$x��ťsh�z�{��h&��Y+���x9�u9%9d~ ��S7��5�� oܬ����`�J�=�*�:�ċ�va����~Ӳ��8��q%�ꉹyiY^3���X�5�x)�s)�w�-���m\�m,J-`hK��f��)�s3d(�\��m�:9�_���YFI�C���o�� �şI�a�R�]�X��d�g':?�AJ{0��P��	.:�W88���W8����?��R��JA��0~��?�^����Y����t��t��7���� ��0�I��y�q�"�j�#��Z5��eb�0��6�u�c��=V�r�h?Cx�=H��!�(��x�5MD�If![�l��V�\�ȴ�@��%�:E�]�YZ��#�bO_Д.GR��N������'4w�&d�����K����ru�q�tϝ'����}O��bq��5���ٕz��,�7�I�~k�/ZK���"�.�8�m]ݲ��7.�y�V"�P�h��<�s�zD������b �wd�z:�'����r2n���P)�[PJU*6��B;�3u O�k��������y���{f��<F.�ҵ^������ S��x�p�M�!��uVpM-ÿ�)��8�r׃��B�����2-i�)�g���ߴ�6ȝ�*14����3���wy�&���f��+q����ʅ�����u�Xk�Y4⨪�O�L�K�%��}����}���N��G*��?F�����4y�c�e�`��.� Բ�'�6�K��n�|��/ݖk��� �I�H��5�Ee.R��h����O�@a ������5����Q/lh��c�K�4���m1��@	�/]�+X�(��&ӄy��`/.���k�oLg/����S��;p�'Qg�I���ӠPA�7���^��:�U��U$�H�Dg��ˁ�@L�tH�V{�怚Q�>?8��'fn�k�
���A/�JbN)���6�Rv"I��-�)��H�f}>5��w��K.��1�J3|5؁���r��߇j�V92�"�g`�n�Уn߀�v�v�s����Q��oƠ�ܡ���ØS��w���2�^a�s������L�({�xfN�&0��F��l;��*���"%d}V��OhdK|���a��S�����q���@�W6�����b0���h�e�ƓӅ�Xz�HfO�O���Y#Gm�kG!�Y֪�!b=��x@ҍ�iH�G�j�M��/��/7:�0�ڵ��Y�(�޸��g]W�b溸�[�:an>��P��C�+ �މ/�
��ȥ~0a+��� ������k�;�$�����Ug��z�B�#|	Q_.��l��Pc�����-�%���������:T8|���n��X63H�)��.1�H�ЦS�i��4�r���(��`ߊn��(Ws~E(}ʋS .�rI]Q9(b���Z�y�4v�mΉ�K���h���Ec��%kA��O��_�(��4��@O���_�:2($�Y�'Cw>U{�ݦ�$�,P��h��������vN((-24��Ɔ7�E���E��L��2�ؗ|#C�c�y���Խ��lMH܃��U���o�7�Y=����%��?� 3L��M�@����#f�>yu!3�ɼu?��+���?O<�S�	܅��ȳ����g��{��]�R�H�d�F�d�p���R�F��H�`�,ݍ�U�k��Œ���F�*C���b��1$�VZnW�(I�/
񤶛�^i�r����pZ;����\{Q���ͼ�lLҏu����zS�(�G���8��B$����R��s1��ܬ7z�j��r�2�򛵺��KN�(�V���>�� ��#��c[��?>շt&4�l�%�E ��׃2�kf<�@y�&�EdR^z����� 98x��#�B��G4m�+�KZ+�Y!06��I@�6p�S��[����u�:"ܭK,JǸ�B�p������֢�B�b���^K�Gs�?��:���s7�}~���PN����޻v�B}w`��~q��J����/�e)̨i������r[(���Ìc39��t���_ߋӌϾ}e��$WN�be��U�E��"<�O���l��$�<gPw&�G��juD�"
rܔ�u�u��|X�����@�[?B1�6Hf&���]ֻ3�ءj�d��ї-��A��"���%U�	�3�«U�c�F�d{�P�y=_�#Nk*�[F�����q7��*��z����U�*��]4z|��q���P?��E<�S�is�`/��ԡB�-JG�U�f!���c`3(�]���*Q���d�<x}jW9@���?Ɵ�'��B�L7�7�#�/��,u��� v� � �T��nm�>��u��� 1�Z�RÒ��cn"D��/N�&�g{�A<�P<�Qד���'�*=ɽ�	��W�{S��Ǚ{K�O5�8v�fzN^@�*��ذ��Ȉ^�R\P8�^Z,���|K	�&R�����S6�|Ţ]]ʽ��߆�{9
3�c=擏Ό�9��mϝ��òң���atvs����I�:�{gg�Q/�H��=�B�]�V�jQ�q�p�< �eS���cM4�d��]5�kc�)��
�G6��� Ӕp��f^N��}����K���U����ݭ���{{J�]����J(��l�jʘ3uz��Wx��S�R����P�|!g|<�
�	<����4��t����uv�#��&Ыs��Y����/����,�RHΰ�������4�L��R�V��!���X'�7l�(|��l��v�1* �Ϸ���Fm��=y�c)9��y��%��,J��-i�%G�V� ��ꔈF�|%B������h��)$�Sz�ao5�.hӅ5��?HQf(�Z��Eٗ�R���_m$�U����s﯏%���F�s���?��
m�ԙZg��K��j*��ߧ��l븞�o�j�	�ʌΑq9�
�!�y�7i���aC����@�\��[�9?/�9N��P#�9g�Ͽ�k���m�Ԑ�o�POٜ�Hs,W>Q�|o�,���c�3D���IbQPdg��D�\��Ya����:���S���&�:`��&��\L�c���ʃW Q�5M���=����v�7�4��Z��{�y�g������dXZH�ف�4=L^vs�uE�.��˫�-�O�V"���f��>�B�XI�d���o8ؾԴ)��su]}���mtܡ@+|t�Ŵ4���w]�]#�� >b�P��g"]%a<z���̉�]K!������B�e)�#+ 5����s@��e�`��O��ǚb|��\�W}BS�������D; EzV"�o"��>b�Ӻ�UF�Qݳ�1�( �����tln¬�1�|�X�ޚFIfS6�Z!ZUɓ�l��j�.��J��mW���BrA[LQ'X�:#C>�WV����\��ǡv��}T��b��aQ�O
��>Vp;B��1�)�q�Iݾkp*^<�AJ}����^�|U��ci�]�Jf/�:��.GQW�x�Ne<����jpp�f��CK�<�	o�i����l�;ꉼ	f����7���}^.�X����#�����U�# �$�3#	��N@P��!j�A��m^C� 2�;���7�+Zn�����&���;�0�R��2u�[k���xW�-Pw��c�i*;]V���P����a��3����^<�D��D
F�$ʛ�a�z#'4�~\ud{@�r���Ѭ�\�zh�?0�7Z>��d���m�����-�Rs� ��%���F��%��U3X�3���� �
.�/�g�-1Ӹ�MV۽��-X��CQn�3���C���&"�w��dQ-A	���+N*�3���B0��N(VS子d��pPA��fEk��p���I�X%|W��d���VI����5K�1�`�Q�yg�'�̢��&���XrͿL?3��>`m�(�j����Lg!|@�����z�!h���;����v8�������&�p���j+�ydlY��&�����	�����C�9���N������r*�!<-\w �X��k��^��4N3h��B��LW�>����+g�Ao�̖� Q\3����/�\�M��hɠ����	�w��7�g�+�8IvO���@��#�#s@�#_�~�@%�'��%�g��m�V��t9�Aw��5���e`���E�!�-dT&���q�S.���?��G�qAȰ(�"�r�5�u����9}�n��d�����9� 5���x�`�t#>)�L�e�<<G ��vS�IV�A�+��Xp�/��GZ�"Fs6c؃,z^��)����-#���?wfȭ�^�&�:tY=6�x�