��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�>�u��?�H�z-I�w��kTCi4�c���	>Ж�A85���
jԽO�1n�����8��.8�q�h�d�w��Eg��������q>��R@�G�e ��5㵞OͶ��6�UpDw�s�T"�%A��~���}�/y�q@�@�	y6��g�
j���
��Ë�%��J�'����M���.�S��8Q^z؉�r��_9��F51xל��k�s^������	�a�%sx[�bF��.���
2m�6_��"Ҋ��_�F���՜�+i�Y�DCP��A���7��dq85M���;K3Z�����מe�\��2�Bڞ[��9�$/?"��v��L�C~n�?��7�F�w�e�/�svߵC��
j
��m.eM����~�ͮv�56��Y�I�c�Pf���T˙�n�5g�����;��6MƯ��%q��Xe��j�?d�+qO�4�9�b�4�4?�{��ύ�������|�Ec>�:�+ZA��GԌ	�������"���r�v/s쀭|�0|l��$����]�����eͭ݉T��X��}ɚ��6�R0�'��s��!��~���S��z�A�xI����$�m�����~�j� ���f��1���f�!��_��2Ǿ�b���G ӉGRTa	���yv�F���թ�vP��^"й�<�-N!�(�e��EwOyA
��!��1�D�a���;�%�*Ҥ&؈x�������0�T���s�P��Wc�jDǥ�,e0���&��p<�Bvd�٪j�BH��q�V��/�~��A��l�-]GI�hSC%�}�0�0�a�T����p��ɇ��:d�HM�LX���Apn�H0�V\Z(���1���7<+]���,'���$�!��ѯ^z�zoQl��0��]��7�A��0k�����z�S��j^�a/0px-.�P��WI���8<���P䲱�0�ư��]5��m�@�!2އX2�i�y��1��L�꥟V�_-U�U"�F��~���I�(a�Q����(�zS~�aU������S�:I�~��5&d����_�x���o�#�6"j�A|,s�%����]�����#�KkD+Lq��1�m�
qk���!q�l�����p?�z�9q��\)=��+���*U�h/#v��%D��;,�A'�~�`���ʶ>ã6�%6*HA���W�����^FWc%+Ś8���v�a����{W��J�B�'�5<���[,s����C"�	+��N`B��-���_��
?E�\<�ɣ�{��E~��m�ѱ�}�ubH�_�A��6���~��E���|�����g��������I���K[|�4������#<Cq���i�+�kL-�kL������K����D�I$���&���j�@`g�JZ֤u!���d�� e�ߥls��S�(�F0G͏>�$�9�х�������{)��Q{�*�b}�Nǻ=����xF�Bg���ҡ�Y˰�D�1O+����c@t�k�~W�(z��
rl ��9,\sV��� p�ג%T�v��oJ��͜R���8��A�%��=fK#�=M<�Lf�����4-��I��/U�$@�\���H4�E�|I���=�.��FaWE��$.���sQ
�OQ�\���Q�R��Ĳ�x���0˟F�WV�`I�t�ȵ�[������Ռh=����}��`��燻5���+��ų�V��X�mZKL�
��(��k�z�8m ���S*e�W@�!r��(H�U�P�F�bP7�3��ԦzX���|K��{�37=v��$�,��,IGn���g�"��V��Z"�Ҝс����ݷH)�� �)�w`a���"1���rPų���a�~:���F���\�?�ǘ"uǪ�+�O�N3��0|>���Z��	�y#�?�d�j+���Jf{̩�0��Yc!7����x����r"g;Pπ�;.	E�w_f,M���Jޫ@aί�޻)�Ŏݍmqh<�G50ӏ��k�q�����b/d�2�';c>�k?C�f�N��[�BI���j�sȜj��2�G}��$�.6�"�J��m�I9X׵�{+�E1���۹�Y9���s]AD��P��r�(�l�����cdq��_�����nT�Ro���Y,�:����w�AbY,��
��xoZ��������񰰪�K~p�|*�w���OE��喠��^iEC��4nǅ)����^`��P/5��-3k���Whoo�>����|st..�.�9����9�*�g�pa*�A��lql�x�#XҚ���dM��
��:��\���0���?���/�
��@,��r�N�Lm��F�4צ{�I�}�[�0�J�	M�B�|8��t��֯�z�W>N�[����L��y��/z��Aj�̷F�|�#Fx�k��f�� �?}��y;%-�M�^GM��	W7s����,�b�r���4�����p������M��Ǫ�����*�SF��t����ͼ�ּP�R�c'�ļ�r����(�J�K����&�%%��ߗ�� M�8�s�5TDw�@��w0��!.%��^��>����^K�Vy�qfC.4k�'h��/�{�+=o�iV����n))j\�QN�B���V��s2�]M*��'v��}�m��
��`<�%Q@��\� ��Zf��\(_��^m�[u<���V1x��^�^�~��~�=u��O�=z��,���h���6�RY>拘��ӔW�Ȱ=��m>jR��jw(=M��|Լ�;��_��gi�]��,|�?:��b7��[�Iv����D?k"�4Csy���S����B�, �l-wkӊ���B�Q�Ե������uv��u!'5�k)��3�)�u:�@����h�)�Pq��=�z�^��Y�%>{��|������9y_��W�+��@ղݐK�(�~P�b�l�渄�g]=^���#
�h�O,C�z�#^pF�YKux��~�V�b��]���K������� �(
�N�����q[�V�����D�@�,Ɋ܈��n@�^��(#h�-*�6�\"�[���2K{�ɹ�m��>�J��!�^?g�f���R˰I�#ȱe�a��xO��)׺7"�'nE��p }���c���q�Zū��C1���G�@�������rK���WW9�����7�v2�K�Z��tO}��:k�s��B�t�G�Lr�>씟�U�g�@��˽&��h҇�:Wu�7r9���׳��T�ڂYūC{�n���P�<�X^l(�md'J�xy_ ?��\{�^��>I��I0PAjYO���c�D�_���9R��- O?t�9f�d����P��i�Dit*��=s�ʦ���]�)
�� ;5��uE˘jo{$O4ó�-7�a ̡��D�^����~޾A�������s���M�<��W	b�h�
v��y3�l/�\��s�AM��$J�w�7΀�����bY�WžPjX�����faH�Ɇ9�������t���z��2
�����C��0<ɶ�(������c'wpV*�P� &?\���%��QQ�[�+�}[F�/O��� �4[�0a�c(ƥ%9Ԭo���������a�BI!��ͳ�2��jx2� �.�1�������	��Y��7F�`���G���ֺ�aYn��=�bXi^��Fȧ��D�N,���-$T�M�l�Ds�<ie2��z��gv�m�{��0�b�oS��0�Ȇq�ߩxm-�����x4(�J7;�ۓZr���k88N�iե�"R�J����	�g�;]��*~@��?�ބ�����Oρ��o�kT�h���_�)�2�?�L���P�;/�~.ĦԼ�S�!n�b�(�����I^�"(fa��~�(<
�D�<��*3�(a5EGw�I��bRO�io�5xu��?��-t�������$���jSx���!|ƤY(�L��=H���SU܎Ǻ# ��<���4�ܴ�;�D�}2z�b�䆔��u��ч*�t;:R� �q���`�I������(�d���v�-Fhs	����k9����z�q3#*�8���/�K�7�0����]D����'�K��m�+ީe�i2\ÔbX��s0��h��Bn�l��P�ի��qg�y�46)���+�j-z��a.�X�!M7��c���a���l�0y�S�$D\��DVDtF,i� �=3�L��v��wX<���-xp�� �vK�&���b��k �������tJ�����}�W"Q�hS�Yɪ8#MD��\��N��+�:R�D�G���mƧ>� ^�r�R�*��Ր�Hc�p�uW�?�SR��o�bt�����*}�V�F�{��5g���5Yܲ�E�!0�1hH[��-���]���ʹ��"�Z�B��"��s�սp�|�B�ԑ�Jh��I�x��I�^m!?���˂/�K�h]ڋ�]A�J�G@y���m�z���lg�P푳�m�O�\�04|�=>�:[{�����*��������������2�#ӑ 4��ze~ v��qݲ�kI6h�+��g+������ u� SVone��F-��[�#5��`?*�(��x���TSի�MqYy�����!�j���Y�l��L�3D���u�Y��@vH��o���4�w}�n�!���$�<�j���.SlB�K�'�~.ó�*EgR��_�?x<\�5��]W�.tˎ���#�W5+P�Fp�^cI*��+؋~/5�?��"a\'���}Qt�q`[��E�^I�g}���oret�����0�Jo�=���X�R�K����#V��_������,E\��A������1��u��dn�yQ`�(���"�C�%�/2�(F6M����{A�y/3P}�P5�]�88(e�>fe��\!N�^Bx [B}�de�����׈�P�&�|d� y�2x���&�ϭ�V+ C�W����wa1'H�	��	D�����r��2Pu+�7L�kFGƭ8|�Pq҂A��BP�Ǧ�/)yΟ\.��`�y&�K7�2[7�[���I��	�Խ��ں���`W*ف�U����P�	�s�d"�F��K5�:`΃m)�G"�>��Q���W�e��@U"�8mˮ�n���Z��R<�c�(9D��Z��{�^�/FP�E��5$|a�aٿ/�`[� ��[G��Ю,�������'��Vn�W�[�ôu���MoP���}VY6�{������'�WԺ�%1��!����_�Zû��ګ�s_ඝ�၏z�i�2΂�֐���	Fr�����
��ƹM."VП�h���2AW��l(����̙�Bf��Z�	I]Y�cG�#?�Ψ�N��oDU�]� z�<��ڮF�XԐM?n�����亡j� `ue�~�j��M(x簯���F���@����kei�+��R��j'�)` k�Z�ܲ�Vax�$QK+����A�@�N��c���?��@������q��/�u�����kf5]5����"Ο)�T��n�bϜ��{	KIϚ��9U1u��{:����JN�>��ާY�gy��������H���9�n��0&��Ƕ�0�Ξl��L.�'����	�R�� ˹��Ƌ�~��G���
i,� G���t���-J��.�~`7NT��J5�m�>����F������~5T��Ė/��Ƿ�o��,�f3&]��{ss�f�>�w�M�l4��X��HX���rS�3����E�KV-�	����5�T�L��U��gj�id��	�W�};?������AN�QXC����B=^X�)d8��,�߻���"��I���A�Ճ�|�b�ɐx��>�5O9/-D�wM�ջ�$�e��n��'k����	���2ҧ��Yj7��eu7Z!��]G��f_F��@��DZ,u�4��Po�.�C�Y��-�*��E%��������(�M$=��KX��<֛��T���y�D�j{K��!�T��(�>4��Y�3c9쯗��6�<�/�4�i�>�����w:TV��8{�$:��dv}�t�~��s�v}(Z'�ս�����/5�����_��jpP�x���)�����~�6ѹ�y������ذd�jl��J���N��!���	-�`��kF���F)_�VA�@��mz�G�z�U6lcT���=j)g�̪"�fAs�Z3�����o�$*��֘Z.$<pl�o�65��U��B�Y��آ����DTX���S�6�Z���P��k�����B���7A��p��(� �^V�|?Hp�9�)�����<���nnP~����2H�׫͍�s���p�ͷ�G��O�6q%K�Weg��Ѡ�S����pV,���4i��nK/��ϫNj2a���_I"4���U���0-?) �r�}d*a�%��{ѻV{�>����pћӷ;�q�!�4�L�v��e��&L�|�fgTSˮ�]��Q�9	��ڇ��k��z�p�}�ÿ��f�8��P�Ǽ��9d��:(�Mp����ۨ�a�X�	&�0����A�ǡ�ܵձ��>�V�fRHD�=�-E�u���Ʋ�9͔�	��^�kG��O����0�h9,?J��Kl6�@�j�<lԆ�5�Ϩ=��p�Ykc����yc��x���s�X���[:�a��t̏�:'Tn �D_����̴��o�>m������@�3��d�)�hϜ��f����٦F�[�=GKpaJ����[DƠq���\�sJo�8�S������`k|�lE�%��D�wP�yb�0m�����-0�+hU��%G�A����h0��*��>��d4�^��B�0(�</�3�����A@�0��~#3�}?����0�̚�K�O�jCs�ۦQ�8%_�J�w�@�
������}�Ґj�|ۿ���j�4$B����u����	%~�]��3$����oӈ��n3�h}F��~J`}П���Q�Ő���gp���&�.[U�J ��S%} ��j����t �7��*�3㼩����&������>��^ס]3.�^�VT���БWB�rÖ~�ƿ�F�xa���8trp]�A��xoKz���U��1z�
G��5��Ao���Bf���f5J�M��n���Zb���Ze=�,��d2��r��%)��/o��)	���@
�V�}j�u�����̦�
��8m�΄s���o�;
{�'}���9��q��Q\}�ʼ�v�mqw���'1>�A��e� �n�G��t��pk~�?׌"-lv�}+Ik��5�R���9���2Dԟ��>�m+t����_��M[,L�6��E�'E�UP\v|�p��R��9��X�:�XB�[��S13Mb�]]��������>=yx�F=ʮ�X�C���K,w��O�$��ߖOo����-8�m��.�P���>����Ɨ��	�l	xe�=	�D�<�9M����8F3�Q>i|b�bQ �.�R��Z9��t��Q�{LYaZ2 �����pc��iq��yY���y�1"����}A�Ǚ3�	�jw�#���F�F�v����EK��Ԟ�I��}
SBC�Y����iB�E���K���=�3W%��H7�E߾c'׫s���i>� ��dc�`Wl+��ӝ�I~�~��*�ΠIP�P:��@}�CZ��G=/>�64!��j�+�Sʣ�2\��\����6�m�k�����7w����p�/)4N72�Q�v�J�%�U���[~��Kto��=�O���v�R9$T�R�Y1�C&]?q�j|�#'~~ΐ\�v�2�oRBR;�%�.��eB�,%��N�k�-yd
[��P�-�PJ�kG+pNh椲��s�Iz������'<��Zg+�������-!��8NT���"dz�c=G��-3f	��o��E��W��U�/ϙZ@��V�"�.������%�H��^hs̟�BJ����j�iô�S�pKb%3��&���",<�ؿ���d}CQ���A���	�?�� ���$���a�q�s����b����.�HHQH�o����*��%~I�\unF{��AM#swBh?w�|����˵א��"ƳA���w�^�J0LA,�|}��-6Y%��ң��FGtw3��9e���.r���GM�}V̀�y8ŏ��v�{0:�<G�NY��R͹��!�9c�kb�qA��X g�d&�i��Sg��u��B�UcT���S��BY�e�	
xL:�iqNU�,Bv	~�r�Ւz��ƭu4���_:�Qo��vR|9;���ܣ��X�E�ػ�^ �/��:I��'B�.����h~y[8{���@0�,X��4�1���|F_�D� Y)LWuQ2��L!�����O��E/ڃr-u�A��y+3%H���r�R�/ ��}yM~�p�w%�c�ύG��*�F�,�^9^�D~	Q{F$l[���UȲ-����~G��Y!�X���Z��oa�c��qA�X��}���{�#��1�I�A�a��o�o�I��ԉ���;�1�n~��(.�P#BPN1D��֙&��"�Y�zL��HD����2s�EG�6��8�F'�Q����6��*W������2��@�Ȯ��Tr���b����r��'�kp6�UG�q�{8��L�zJ�V�u�G���b�j�caړI+<��B"�J�<0k;)G�������7��hMx�o�r�����v�{Loy6�F;�ɓK�Y���D-��������?�x)b�ƒ��6S��ަ���~�'�;_i3Y�D6E��pȷ�T&����Ad����!0��^���7F�S��L�)����Br3W�]A����8��X7�o/��*&���m���1���l��H�<�.�q��_�NYքD��*Wأ�sh����!F�l�f֕��V�Z�V=���V��;�ms��X����7��q �	�Y��������	rO=�Wz�[Y�?t�-X�7�Io��3�5!�0�w[�G��"�c��c�7;֏p�j,���s?�Tr�o⛤����ls#���Qb�:��Ҏ.������[< �-J����(x0��Drx-�[�L�� ������($���!��&�|����vP8��>�ї��E7n�O#��e�:�Y�tguj_9bh��;���N/V�]*}R��!��?�1�׋o8�:Fk���
�;_ʶ�]P�I7�s�a��h�#3��#L�G�3O���Z0�7`�]�g�t��0z���F^�ߏTpQ�lk�T����T�Ӹ����y3�ϫG4��k�O�I�
��{R��9Z��򚭧�b����P�(g݀��gv.F⟜��/��y�n��d��u��v�{aY�H� f��
��i9Gn����E_â��R�h��^6�r���0����9��YY&��>�d��o�Jz�pa;>���G�T����>�%�R�R4 ��k�<�"&4C� ������EO��������v�N����t�I&�yQ���QtL�:��s؜l���t�]~��}A��am�9�� ����C!�ScCR>��*��su�p�l65k�K�P�:`����̽�=�-?�K�����(:�hh��<�qA���)�;:n"Qſ�w�9f���X�B�8V�E�d4�mXz���&�U�'e�A���g9���!䍙�	-
Two��R^��s��'�Y�(B�an�FB�}7o�;i���y<�y� W��Pߌ&W���bmtAq;11��%NG�Y�Ω�?��n��A��v󳠂m��f������|�)��N9��L>�0��,lX?�yu�j[?E� 9�21	��/�\��� �!aR�t1;h��S�w�h�Ϩ(�N�Vl$F�?�gjTSZ-̽�ح7�ӥ��j�	+PM�)l(��� V`�2'��Hy
�A�����~!�U��kl�ۖ����*-ţC`mk� � ����ޠǖUb}-����V#���dŷ��--P6��,mx�.���̏�K���	��	���+6���dI� Q)�AZ ���y2�.u� +?��=�տuF�l�����b��
l��t�A���H�WC���M
�xkmC�#/ҕ<U+w����7�.H��h����4�.*� G�[����A���^I�B@E�����T�#M�+Q�u��t.T[������'��ɰ?�q@�E�?� �'�bUԬ�H�
�_���p&41��؞��J��s=���~~V�9�m���VW?9�`bCd���-��^l�z{����	a9������0=:�co�x斟�(�X�]�3�0Ω��K52��e?~��l���ƋS��]}k,�k�$��}*U�`� �AU��f><Xa��~u!���6_�Je�_턥���H|����9�E���2a����3U�d�@�����+�.D�� *h�5Kb�[��)�*���y,%8��3n���1�ų��W+��s��J�|��-1��@u�k�p����_6��Lmܕo5�ўO��e�\zgx<��3dc.�5�\w�� �ٓ���J�*Pl>)��	<�@aD
���k�.����Elϱ����A���T��F*Z���E$aM��`Eb<� ���vQ�ЄV��Կ��gõn�����у�Y)���;��8D�Z�ZG�����T���=*��\��9��I��yy�8�����a{ ҿ9��j^4��;�}+3�LgɼG}���Tr0��[*���`� �a�F�C���t� �2�c��gn=s����L�}ȁ�6oP���r���x��>*���Z��C�鑣�~>7��=� j��E���;中�^�z��}T�:����n��.(4��Vg�j��kҙ��މ��S-�DRP��`���V����@q,����l�.ܬ�o�� ��_����k{I+��Z	&vK�&~���D	�3�@�\W]۲	3����9� ׈���w���$x�J�~�$`����ṞV
���{��}�Uԗ�0�m��i�s���B,�%	����Ld�W��td� �j�]���|��7?m~mx�rKl>�='�y}���G�i�C�ѓ�H��O�/�U�C@O�����q���S�*��NV��B�����oүr�P�Y Py�ܼ@�.�Hۚ�VAQ����|Ð�it7l+�XR����f�7�\Ţ�.A�p�,��a�%��@F�C�9��~���b)�ګ�[ H��@��.�H�6Ֆ]����55�t��6��A�`�]�4y���7J"c#zI<����Ļ���'�ɛu�P�tt̘��pa5�N%BS�d�����H1���W��˥�`{+*!����\������qĔ�����C�R>VP�{V��Y�]��h����&#�����������K��y�{��(��,�g��ܫ�V�3~1ݧ�H?�M���R��I��mH���EB��Fm�ɬg�><�i$B���3�C�}-��ϔ����/��"V����YL^3@���C�F":W�K��q�6h��) @sV�����yyk���[ɹE]H�0���h�tġ��	��%����(���)��0O�U�W'�E�[$�K��Z�?��E	tK�sL�	A�Z�)�V@!���g����w̒���,��eO������,����� �����F���b����R�$͐��Ʋ$��>Fs��14;WƧ�
D�8iG���a�K�M,����T7K��7k������'�I�t*��v�վ�R���	Ϩw���aܮ�vx��Sjɵl��72y��|��@ԭ+ѭZvl�lG�Ŵ��oG�]�w��V�y~�n�L4�k
[���j��ӦVN�=zk�\�m����,q���K������B1��n��u���i��.4B+7�iVʉ���|z��O<���1��&=��~�O�|0�O;$3��|i����Xf(8�A}�5��L�4�р�+u�뭆hy�e�_R4,M,--�¼�$GkQ������va� ����b�z��D�h��3����M�$�t����q7��V���4E�<�gB�G<� �Dj����*���|��[��.%�EC�o�Q�(��o0�3 {*��C�´�ő����~A�_"���WT�-���6��a�:����0��u�D�HH$�*�]�8M�k�7�����^��dN��Y;�����2[�:H5y�m\���\7Y%�T�斬��=���H��w�J?�u�(J��P)n�������&'��<(q���5ZՉH���x�����)~��"=o�6�fLm��E�ϱ۬�I9�}�9~j^EkZ�U
YL����zq�t��G�,�f\O�>22��	$��qF�m�f ������8=Hs�B�*���?G�����-��H�DU��v��@��N^X^��϶=�?�p̣Wc���7�)���(_�h���me9 Q�8��h�4��/y�c��3f��d���0�'���8B�X��cQ9EH���!њ)�{�4Jݖ��I	Ӕz��)��_����q�|Kxl��ȇ�7��룣�5f:��9�L�k1A��)��i��t�N*<ܸl���\�q��iHv���sa#X2P���y	R$��d���X8�8�K��N".��уH��ѻ��j����1}@�>�������z$�%i7�,g��V����C5HqMzC�π���?n5:���҅ي���{���N+A�rV'~����F���~甕b%�Ak�x�kX���H(�{��,l���>�G��,Vo�h�REV�{1��Т�(K�q;�9eR�7��F	�<��*}��x|qj��Z"��a�@.������G
^j��Dk���x�>fPI�}ˣ��ɦS=Og`�Vv�;܃'1��nC3ƍ��W|�f�޶�R7֒��=�&��O��QŊ7�J��^�?�JL���]��ޞW3PB�ϼ��I���.�W$�E�}�H�6�s��(�M�p�+��Y[��1Xf��:<\��e<9o�D�轿v��(Hf�_"ؤnS�s�� �֨	�/+ģ�v�c��׆�6�g;S\0$���@ ���g3�u�� �lbͩu�؋���$��׷r�shQ�ͧ� @�*S4&FJ�L���a��|��T��7�$!_�똯5܀���K�.��/�拘R,����A�I
R��/Cg�Y�3nz�MAL ["�,}a܃d2�3����W��b�^\$�V�щ�pG��{��E�hv����0^+��s �'��_l��ݴ���!Sfh*�Uc���{5���ai/E=&�7�ˏd����=�N_Ê��8�����O>a	pJQ'�C�,��ء_y��4ײ���gʟEP<k�G����/��sO��q�!�[��5tW�D�����O	C{_��~>!�I�S��8�Z�t��b���<9�����-y�j�h]:���:2�?��q��k~���EՎ(�pC/�ڶ���i��?9H*d\J������"����[ы35oQ��;e/��9s���ș�\V4�YH�<����wbFRc�j�m���@�]�8dL�)Q�y�d!�n7�SwV�b���WVJ����m|ؙ��}��������?Ú�>Kxw7V��Q|�:�}��z;�C-�ءm�P�5'��.�5�m��J�r�v��Y���1����Uj~�,sK�3������4�W26	����9�a������C���~\�Ӡ�:�?��{�s���ng�h7k�6�<�o��7Y�n�TS�~��?�}���`��Զկ��v����vtv����Rq���).�{�}1t�F0�3|%�A|IF��	��1i��^��{5��i�X=uvkh����,'�θ�����[�X3v�ka0)�!Eqeg1hH ^1f��>q�|z,�����H�rK�j��k �������n��%q��M�Es3�E�vۘ�־jz�8W_Xv�E�O�����=9�:)q�kD}�fW4j���E��ـ���Î��9MLL�b�Y�����b���Ԯ��>0P�N�S��9놞�9E�[���G���M����X��A�Aa�G�MR;�Qr]��8�.rN��@o9;t�D�5t=�n[���J ��-�C�y\�)�0�^��s���K�8��|����}��TC�F�$���O9�?6��hܾF��4ˑbdc+�ܮth"U7E�b\h�zD��7dY�q�8�u)�|}]�Dq�(��݌�%�����6�ː�#i�����&�.��E�+\~�8L����uR�����dUNA~�9E��K�_��mO��ԫ�]	U�J�Ǉ��J���J�Ŭ+����C�I�cԎ��:5��՗�M;V����kQ�w��/፹�R�&��W�8\VGN�?v����4�b���-p@@6	�ƺ�
�[�>��)���.�� :��0}�6��q�c��@�����^���h������"~�
�d6p(p���F�C�@o���fX"H��y��yZ?ւ��/�|���mIg�����h���g�sҳ7��l�k��gzo�;�`CH�C�i>��v��Z�,�ha'>z�H?L��ة��}=��U�?�~��VkG��IE9Rڍ��y�1Fƥ����)���}�a
�VO�ce,V#g~�K7�'*��F6A3k"*��Ky[r<�;����(�6��Ϭs��fv��7�,\Mv����܀��ʈk�>,�>`�� ����x���$�8F�jfM=rY%gh�-."��H6�$�q@/�7o��� ��cd�o�@�@`�o2�������5zx~ȡ�e=���A~�8˟Wc�ok��\����Ҹ8�ل7��T����AVCj �Ot������� ��.��=����d�V��vq
�Q����H#��S��ڪ7��@	���_��ˊ6�g�}'��0�]��W��Q܁P'��������J����4X ��3�`�\�d2d��V��<�G#�}�!���E��=���l�.�U�u�&�J�|��u�N�49��1��Q"Fl�Z=�dU�9T�t�;A�z��>g4K�������#�r}�����W;�G�����!Ep��=���G���KN�W��{�NW"�ɋx��̉���w�5����@�s-�A��3R�DJ$0g_%��s��Al����8
˷Kj��$N!%0�p�΁G��$gI�$�F�da���p��{��m1�%�� 1������f�V�,ӥ1�^b��ȴ����q\�*׋���n6+e`���n����o�N��C� ��(`�������J��z�Y �=z���_]n���C�o9綪�Wd�m���^����!��( �8-���\)K�%����d���p�ʼ&$���B���o�@V?`�U���S�J�Y��m[="�B%�_�j�;����K�R���$��UW�S�"!��� 0t>pd����f�_�µpDԞ���4�D{	��*z5\p��<-�]1�à��]�Hk׊iQ�i�5��c�B*��Mq�����t��|~��<Q�Ukt�sk��m�V��G�
��o� <x�G-q��U��l{1�[{�W���Uy�YDO��+$S��&���Ln[�BZ��P�9�4y��w�resm����*_^�k~��SL?����f�L�$h�bQhT�B[�(� �r��
Z�����k�#0z��U�p�ȟr �A�+���oV��N��B� ��+�0~���Y�nD����lG�)��޽܏���2���+e�cŭ=IB�_�T�cC|�9���S��`7]'Q��%^)���rjv0�x�>r�pӌ��$�5#k���|+k�֔.��-�&J�v�kn���|:A�����~�*Nu������D1ǋ��l�L�������@|hgВ�����ʷ'�%�}ފ�ǜ���� �
'ZXΘ/��b��˩N��`�'��Ҳ���^��1�ҟ�[vo�Q����D�uy�KdGvn(���aR����8U�	U�9�eig@�d"�k"�ȏn�ۂ�����f���ݢ�W�o��M
uﶌ	81��i��3|�t\��b��ʖ4�/mlV����7��DI`�u�]ܺ�<a���RE����� ������q��;����Z�sW=��<ӗ�e���\1�*���B���k���X����q�(���y+��2���y��ʚ��������-��Ī
|:���)*�NL?�bd�I�e��TDZ� Q|ڏq���W?�L�
��z[/4%YDp̞�Gy3a��E�^�2KL�Ϋ���:Ü�}uwpQ!N��P�Â��Y���ΔOj�L�'��r��E����>��u�1ϸ��uc?����m*�O2���dą�J���V����~Ha���=��ƴ
Y��n�M���[��1��Z"u���wv�-HLk��^uyaTz���/��E�(tgg���C+;�2�����7����������M�B��V��n�����7��q<�)L����h��f;��0��@��'LǪ6+,�^ ]t�^�6o�]�yf"
9�%��\M�X$�З5������{�+���薦�#|��xJ���*����*�^� �8Y��Ac����(2Şi�g!Ure�x�vyfǙ�ܗ�x�E=h �~\4�L��C�U0��"+��JLĖ��4��P��"�$��Sʧ��dl�2����&�">9/��OvK�����e�W�5z#�s7�������tw���9��mJ���O�1C�>��@�D���7��P�1���)�ؐ�m�e�\2�T�r@>�B�b�N�O �
�>F�f��snr�Ȅ�1q�mo(�>6g�c��uF$^�#:�
��d��b�����sB ��c��QM�B���b�((b��!*��y��k����P��""���k�?:��B��!38��"ꗛr�,���Ѡ	����ƥM՛h*�h�R���v�_?��m������I��O��(����7�y�w$i���Ǜԛ��'�a&���s=qǑ_@�o���1�Y|�yu�n:B���a�!EK��Q�N���엮4�\�,m��>>�I�sGi�áN̋:��:�ko��F�m�>���1l	J�R9�&	"��h{jo;Ez�ۢw�.,��"�ddf���j1�.i��on�����ϯjͫ�6ΝO	�D ׮(�_��y![N�'X5�����?Nr��ڻC%]Y�Y�+�P���oeTM%��f�$M7��`3��U�a�����"[B��U���Mګ��T��) �ˣ_���8R��M~٣�^n��6�6�ǿkC�Fb�p�!U�k{30�ݱ��Z��d�^ܚPٳ�0���G>���]X�Z��ß���Dߐ<Ci�����ȵC����%�I������(�Hv+5P�z�WS3e�\2�[}fc�)HJuE���b�6P�ӨQRe�/����ﺝN~�qZ��*�mzIP�2�β�c'r��l��g=h%�;�K���[Ä�c*- x7j���-O2Z��Zj,2����!�Uڑk�_Ň��10Tf��O��R��F�e��6���\P���#Bw�q�c�����F;�{̘}��eS�A�<JT}F�m����ߟ��9f��|߯ ���i�N�l�k�^�4�ɳ�Ѳj��X��<�(5�z��0˰|K�4�3��o�ή����^�W�m�E����6���+�y)�������2����n�ir���9���i[
���z�����[Q;�.K�Y�t� � �M8!��M����5� ���gF4o)�l�%"=}��2!�A��ʴ�s�J���y�����)Tw9�d��*t��ϗ��-�?�Vs�t\��&�����/Ѱ9��>?$��������!�a #_�ū�k9Gk
� u�X�G�T<��3���f�c<ףa�+��N8��"vc��O��g/�o��^��{�Τ�ëѮf�}OΡ�jXŕ�ڎ���L6ˉk���7Vl�;ė��ҥ�B�B.��Lĺ�x��ġ^a�Q����L��pC9�����Z lFO9��ߙ���[Ϭ�&p�;qzԧ0����W8�� �<5�����b��\A����B�[&��$�����r���,e\��q�;�yu-"����B���=ч)N���
NY�k|F��@���N��c�"�D�x���BX+0
�t��f"�f����m�]��"�>��#���-����T1�@���:���١�d���i�朖y�2�,[q���y�A��.<m��v��j
j�	�����\�+�H��{A� )n%�"�د�R�?7
��?t����_�
�9�f���s�@�x'�Uq�#�)S�^�l\l4��r��U
	E��:ċ�������<�6��!�����@�X��IА�;?�Fh�.q�(�Q"����D簙%f�2Q���c���k�'śzX�S�(q�_�S��іP�ނ��׆D�(�fc'��BLP����s_��I�@�.%U�5�ĵ��K�Z�~������Ã)2l�mQ�&�(�&��]�s����]~�&����=�i �P`����'⯌�v29�{-9y��?��G)�q�.U���	CV�S��C^B�W��A��pP&��+<m��&pt�[�qq�-��ⴙ�YX�.4'��o����Z��PhTu�}�&����*W���趃z� [2�"�r�}�$ƃ2F��E��4���R4�1Mʼ�Ik܆�':J8=1�-)�u�r�|����7���	_@g��K��F��?'���4�kLh�`��a�:��2\�H�ǂ��j�>����.�K�*W��^s`3bRY4p�'��[���۬Y�憹G�m�qE����p���G��Y��mۂJ1�����p���U��8��a�>�b���vz� B%��w���GU������'K�W��<�^���1?-r��&DQ0����~3:���C�;�"7to:�b-��]�U�E�a��%��J`u0���) �a"
h�=T���,�X0=��<
9�G�Nq.s��U�o���C�q|_@}�ʰ@]�d�i�>���z��k�4�K��Jv���KRu1����A��-2�		�N�rџ����_��#��3�/ �B)O�/

Y^��!��B6ܽO��������qdCԩ��\Zۧ���3��#3L�{F��տJ":��F.Ff�X����h�c^W�etV˷��,{<��$�3vV��Pţ����Z��мKDF��av�,e�J�'����i�G��f'��*`�#�=����Ve�6�����3W�{e�t�~������8Pۛ���G�:���d[�fF8���͐�8�J{��`�C	E-�
�Tl0bTU(uHݤ)��ۢh٣F���Z/n��΄G���v1��U�����Y�	�c.��Xy��7%����;�ѩЧ��\!��2�R̆�*կU&��s |�>j��� l=>��һn�����@��!��[r/�)z|I(��D��	$_ߑzO�}K�Z�R�m"R�.��n��`@�ǚ��-�o%�q�QX�z��K~�ܕ	<H�3���>�uUFI�s��a�� ���޻�a�D_M�n���+^�a���i����3�R�E�2ި?e��\�+�f��=5�WV����z��c�ⱸWB����D����Mp���;� ��w�Y��Ҁ�94�jkk*���C&�1v�,�l�QxL��d�DJ��T]�v�l���_�=՘����:���I����۵��̬�/��Q�@
��*ύ#�IW�_m��?�7�y����*� �Ѱ���!^��~{.���0Ĭo�@Z�`���H`ﯝ�H=���G
�Qu̩b�|���~�.���҈px=:�f��<O��M����q=�a|H��c����eE�d||���N��7�`i���+�BH�A7�n�I%b&W�~#�n���KT3�;֬���+��2�0U�P�]�����&������N��j�ҥ�^X\����A��=h��J�f�LɜO"�L<��v��$�ܲ�PF�W�y��x����L�ш��(|���/���x�
���*[|�B	[�v��,G���T-j�IJ�6�O!�U_wWyD^	!�����6��7���#؛�3�aա_h�S�[v�-Fo���5�{���{�9W�@�`B��3�թi���_�>�4�2��r�x����+ܞ��0�9�F&��A�\�"��|S�<�2x�O2� ��)���[ބ*y�B�AzC��IIOG/���+z�}�d�t�gYFL�ü��C͚�=�C9�
��[�~ϽT/U�o
�A��@
Q�z���fL;��A*�-�?d�]�*,����(f��m��2��ڣ��Kg��šoC�P44�L�{57t%$h�|H�v�]z�,q�.����b��s�2�C0%4&���+e=���0�&رń���L��hҫ{KV�?���!<���5�Q�0�z����5�z��2^Pg�r�)n�k���߅����rp6�rm�j��G� O��gG�фu�͒��w�~������^^D<z�n�^�)��/'�O��_�iBo��7G�_1R�����ϥ}�����<xq}���Eg�},\l�n=4�$|�_�cd������Z@cF3�H�>���-i��֊e��}�pb/e���'�7����.���;=�G�:�sy��� m6���e/�jE�ҡUQ:E��!^$�D}��l�ss	X�.h�欬��y�bI�Jo�;@YX����g��и�V��9�����Zb��A�ö�ղ�qA�9�!7��Q��~Q��#>d�\Q2LXvnz��#��tBB�@��U�V��ҥ��a���=3�l�j�$��0�87�u�>�KZ|�ٻ�*o�h�}f��Ig�Sa�;m��h2��0�1v��Yd��c{]�W�6S��A!���a*��b��2����:x�]�K�1���=MqvI�ng?Q�����P�|����&�4����	k�t#.ĊkPd�$`5k
������0	���W��&j�j0���m�4�X��ݳӛ�}��u.s�-$S:�L�m�j�!�����LD `w��q�	+u�Ո!�i�v���ob�M)^�b��=�o��k�7��b��F�������+$��P����Mn� � L*{^ξ; ޯ&��=kl�>���;�^� �������>��CT��OO��!rE�(z7�8�
b@��b�Mg�!Y`���oP\+`O+T��\�hZ��k[�/w-��i�hF��)�	���	W����C��_px�O�2���Ƒ���#Z|��G�i�h�F���4_�|��e��R6�R����6ه�j��X�e�\�����|� )�X���@��y����zN��n��5d#��@4p��o��O��twI�W�aՉ��>���FO �R9�JA��$b�Ç�1�h�*m��&@|m���W?\�+�������Jw"�����.O6WX b�+�p"�d��
�����M�������
ޔ�<i���A}W,Au��'�)e����]I�&�p�a�r�X�s?����1��j(A*5�â��y��j3qg#��6��<��Y�K�(v-!|���4��sv��wm,p���[Ło�V�K?�sfuh�/9�مm$c�8	p]Mv�ʘ��O���!c0
K�
\]Rv"g�Ϩ��hkE��mRd�9��U�I07�
��~���������O8��M�W�rw�q���H����h�c�h��G�f*w�<���!�<P5��1?�_
ӹ�(u�<�����	Oi�l��;�4(5�wI�e�i(?H�V1j�m���p��o�O��a�q���+��G��#��,�6	.d����?��E��(6Ć��󰌲�t��<
�����kcb]��x�Djot�C����;A&Y7�����M�V,2=i� �g����̴��`����C&���zU�e���~BR���ϻ	�B�CS�cʊ3�u���G4AAb�6��[Qʰ(�X֤�_�
r;���Y�Ŭ���~f)=;�΃����m�X�X�Ī��CL,@Sj�cޫ�!���& �
SN��&Xp���Jˋ�|:Xn�# ܞU}���QD�p������87༧����a��u�Ac��2ǅ�!.��Y�",u���F�k�U MP��qq�1�>�����/^��������>"߰D[�8V-��}�\�G���И�� YG�$�":m3����_03W<msP�{;�˸��^Ȍ�UO��G����b�g�"�f��i\�;d��:��1Cy�C�W��oȀAz�!�S7{X��1���[�¶�k����%S���t�7qv�� �6i�Ř�hd1(��k;�ol5����Z����86Z����[��-�&!:&1k�H�S�Ś��˃]0Ã�&�A�� �|�T� =F;o���f
ʺ='������p�",���!l rz 6�z�!O"<�"�Ch4�d?D6BO���d� 8��uA@�;c����*��`����"vi�ӎ��֐��q�3 =�`�J�v�- ��-/�M��y�������,��1���Zc���^,o[�xr����SM��y�9�qǷ�)���&p���H8صR�D�l9������,%~�(�'qĩι�@���o�����7�^�|0�"�˩�iu�7(c�i�Qv��9����p�@���ЌN�4�:.ղ�)D��)�Q��};�'J�=���O<l{W�*ʡ���K��/�upq��]�^����mGݠ
��Tch-�`�d7�;�ƽ��ܟ�!ےβD�c��}|�g�"[�G���ǈК�>��������=2�����Z�殉���%4�� �l$�$�-f�#���L�LV��@F�j۴�g�;���PL��f+|TC��cڭ�I�V_*��S�ؑXnmݰA��	u���pC}��#�r_�Li&\p�	���',���O-%Td�3�J$�cIe��t�����jJ�K��O�d�T�5��iUz��lZ�4;3�)�nN��i�Co6Q��V�Dyl��X+	�-����m���2/�CВ~����o4𦳗!�'�
O�����ԕ�K+���� �އ�)�\��@O<q\�ȥ���a�2֓����d�4��!"s��"�#.�"m�����9�nSg/2��sw��v���9����[���Z����I���8& |6�7lS�d�~w��*������Cu���3{������M��`��u�z�
�4L}i�D�Kdވ~�ƥ%��g�5���Ǣ%ֲ֮����od��K@�����,�,}+���1aas�$N�,�ng�3%HF,��f>�$���Q�"�X�@��w�e1�콇�ϻN�Yˏ�6b��R�^�X��(tc��ȭt�\�qS1o�$�	�JM`i�f��NH��V2�[����b3�R������9����MX�S��-��g��,�=қ�ub�"���,
��s�ğY�'��_�vNvK�^����>�)��_5FE���<�I�$,��%��$�\斎�RA�5~c��m~���S��4�`bM�h���9��{���D{����?[#z����)�i�1��c+�ͮf`�Y���**iG��9F�i#X�-�u<��Џj�h�`a�a]�ν
范���"� vYU�c�{Js���$*O�.��t�M�O��cF���� ޮ��o: �zҙ�|F��W���)���6��_�,l�/m=���*�k�zsRnT�_m�(y�Ò��Kb[wN��>�``� $[qՋT�}'6���hC�M��/�)�ŉ�~mјw^��IP�	�R��=�<�O�)�I��6vL3��P*̰=�!GI���3�L億����g�Z���2�n���/�1��*�Z� ���i��'�����f[��^�~�%���m�&o[�Pv�`�eMr���+NX s\�Urְ������`{�M�$<������Mո�U���������eW=���a�	����g�hn�--~�]�2�J�r�#3ų�I=�U�?��%���ʑ]?_�F�gw�{t~]I҃Y��@vIv��V�?~,Mf�j�|����I�t�В�3M3����Z�{�ra��_'R������s���p���S޾֮�����)��kc /�JQ�/�p��� ���|Z��f�~l`�9����=~�|e�>��x�*��Ǌ�륾x`{�U/,�����.�AH��.KNX�)���/����Ր�	UK1������b/%�P�����`z��P�P�w��]!u4��/�&_U�F��;����Y8R���wm��as�1Lʒ���Dg��!gk�Ym��f]��~9��C���׌���* �v˸]�T�{N`��}�P�^�$�/�]����N�!�����Kj/���B�.�"ßmAa #"Q@���}�#�ZHFp���`L-}���/l�]4Mn�Q\��dOT�d��!�⻔�$�3�Z�����2�=A¿���ղ�� �٪�U�HĖ+�;�{_LS\x�����ӊ�����H�c�}c&삈��U���B�v��"��[�T�@�{-�#��s5og�1��wj{��l��ŗ��p�KDIa��s�Z(t�Z�<�5����N��'���jB���<Bj�+�-�#@�N���Z�<Td	�4�C9N���+�6��'��p�7�?IM)�ӳqT�capԹR��j�Y/g܍�A�jZ�!��i{lr�6A���Fw�0��j�����>�d�E>�F6����M�P�Q;��Zʠ���^��`N��B�Jq���"VV���0�������@��X1�h���_���3�6������궕=��!��/u�&Y��V)�����҂O�ז������\xi��L�����E�����PB�uJ.��A>�H�fK��C17�Z��n��/�� ��c>���;���������n�I�m�՜2�Ͻl���'��rp��nZ(vv"N�(݀�n�uI��vRc��P�a��5���]�eF���.|`:�ayQF����F��}|�`Y�Xe�v�+�:4������o):��9�ν������nt�k�d�{tC����(F7�֞*m��	���5���	3�ž~W�e�ֲ/��}��?& ���<X�X�G3���8�n��Qe]�t���=x�*�3���Yh��������I�24�H�B+=��u�:��
��đ�	�b��g���43<���/>�>���!G&�����W���톥����u[�'(e�䳴��/X�n�N���_y��=^;GO��a�Y�Ie��]�iƼ���7/.:���H ׵K�zC�+�ID��d9�Җ����2NZ�l.��+ʽ�<�=�g�8q���{����@��?����%Mb<�I�-���4���r�d�굒����ͥ�ŵ�j֎�"�aY�冷ȓ{��	&U'س���o�֍P�μ(J�po?��<!���6뭩{���I�6�%�O$p��5����ď��5� -	��+s�OU	~U���������M�@��A��urP?�|���e�ى���{�3�1����$��p=yRˉ=o��x�'�*V��߱VQ�$^`�gK�+T�Pݡ�[ļ���\Bb៕D�__��2Z��8�3�k 'R0������C�a��۞�{�� S,�������p+�}����i+��<�W�z�ݜ���>@e	�_�]/��Җ��¥��X�Bs��TvO�� u+�m^��AT�<&�D���bU�-E��>�&�\N�\_ٽ�����b�E�$眂����L#pxS�#0���\�.��9_R��E㻌����^���:����G�v\U��#����T���\S��]P��*����% F/�y�}okw���|Ǌ�����j�mo�o�:�4i�\.�e�k��m9Mbf�#��Lf��Jݕ������͕����IF�nua�3Ci�X�z�3��C�I��8
�&U��-p=q����NE���vQ�y�YzD\�>G�b����Ι�f���!j�%����(�
W�p�=��R�=�I���O�x���)"lVa�3�#b��]�̗�0�m��qӓ(�k�ͮ���6a'^���j��֧�l�f�4vN�X)t3�UD�mO�E!���@����,4�sp�8;\�܍*rOzm��;���b��<QM�<�W8���V'W��Z��@���`x2� 7�R7�s���R�n���':�p��@E�u��@�����P>\k[Z�C����\N����͋ɦ�1�%>��z�����-�p�&��xBbN�~q��j�^����:���K�X�vr��|xP�y�u���Y`�E1gL�#��agItP�k���\2��>Í�b��_љ7��P���(���w-Fa�^�������B9�}g�S� {}��G����{C��Bl��1L���1㎳��G�8q��;@~y�_R�~��T��A}}v�����/d��tg���֩e�o�G�B�9�"O"!*��7� PBK���F�*-�ƾ(f�N�l8C�Wp'V!��h������bN�	�v�{'�4C=��U�2{b��j"ʸ��v"o�AW���˻b�����[m{��}�M�Le/u%k�d�娶H��~��b�2R}@+
U��0?2
-��h����-�F[t���T!i&r�4��G|��TH�7��l�yb@�`��2�r��Ҟ8����U!������Z�y6� 0k#jZޔ~?!q\�i5�;�N��j�D&��(��oJ���V��t��Tj�1�.	��w^�n���I�X����ܰ���Z�p�ȧ.Kx]"Xw๩2�S��oKԽ�$0~����Fbƒ���> ��c���o��y�z����ˬ��3��[�d�X�����)#\}'6K6����Jqm+����ޖ𫞋
�������+��&���:�mv��yυ�ÿ�U z�4�Slѓ���cN=����\g��mQ<��	�/Bp4�^u���:�Ҵ���N��حw���?R�;'x������,�M#�*ޚ{�~�{��F�~�S�[�+���X�����xd�-
���Y9İ��G?f���Y��咙�2t�^���$����Kk[U�l��U�t���$z܌��$F��H~�T=�$�9�
,��.d2DN�s;�8�ƈ���1d�p����~��Q�X��\W$�"J�4sUc�/�,C:,O![19+.��_	�pM~}	ɯ�Aތ��c��S�Iu����q���Q_yV���M��)f�*&��������U�X��0zZ2��uM���E����?fA"�i�k��$�Dh�kF�[�`�5W��m߅sp���O�Y��J�`�,��#���>pP6�L�;�RB��T��zQ*�H\�����g@Te���������-���s�G����x�N��� �ر~��i'�V��7�%�0�rc����=l��P������r�;'��ȏ����d��$:�
6$�N3��#SVjɢ�B�{����n�}Sis�Z}�vr.����dϔ���Z�n��0c;*�hZ���w2�(�k��+@t�`ЫW'�@����p��{>������?�/����2�+ⓙ��$!���c��1A����m{��x�X���V�0[o�$ޒ��ԱIOl[�M�_�w�}��o���s�Zj�I��%���'C��ݐ$�7��A���(�`C2�H���?9)
��Ã��G��+���Y�&	\�T
�e�D*i!��Ra���zM�1��ܺTQ�iK��eׯ�WN�E�<W\D��[�ֵ�_t���"�;꘎�1��	笌w)��i�@=氎#��u��U>*�V$ep��,X�=�\;�E�[�vWH�A�-��ì�g
+���@W�
��v�h.w�C^���G�:�Z1s�"M�ܨ�>��nqd��]O=��ʝ<a���oy��_">���V#���a䫎^M�#�f��.lL�P�n��k5��݄0L�)�b��y]0V
ziN���:��j�c��8��ӖʓǟyO$+�v��?���^ӚU}��I����!�����ϵ|�r,�ts�E��	dg"�i�M�9O�:�¯�6#�E�-��h�=��)�[��4k��`$���#"�]X�bS��d�d
�heG�'��6����?9:!�����g�m�$?�M�z�~��"���(ڝq���C��Q\�c�	9P�*���|�Fq�y��g�wB��`~����85��א� *�P�bY���xq��]V,Gh�q�Lz8�obU|�{��7��� ��~�K� �F@�� b�L��Rh�56F�C�P��\�0�=��CB�� >Il��X�`�b4g:���9:!fh���r/��p�#�?v��n�Օi��(6�HO���ԍ�%o��z?o�D�1�A�a�ͅ�a+˛��v�]����k0l��gmښ������;1ֳ�m�}8���V��<��<�k!%�)���;͡��H%�%��a�#HoM;��#�&��[I���S-��p�8��y��/2��Е^S~��5ƚy��7�A� �xӁ.�RY�#V�'՟}��b�Y!�P����R���L���:�6�fK5Ejo2+R[�h��='Ś8�l�2��1��u�uZ��f�P4c!ޑ]�x������[%��ڬb��oK�4d�p�� 3�z�6�m����9�=�ق}���=:LeG�?��-�����0�g4֕�����s��;���*�gI�5�C�Bn��~Þ�{4��s�p͕��|d���huJ`:{ҭ}���QI������zӤ`�� נiL�Q0�>7(���gSJ�["�!�x��%��c�RIc�f+έy��q��)8���1Qz�%��?4���Ȟ;�\h�[�  ����w�и�͖�9�$��Jk8`N�yDY� ��L�gDB���	���E�wWge��}O�Z\��n�y˰�\	�� �]�A�t
d��V�r�T��eǫź�	��B�x�x涤�qC�b��y�]�JPZ������6WJ�R\�X����Widv�}�o�����Nwǅ  ��d���O+�%VFt�ǔT��D>QQ�ǖ�֓����"	���X��Q��i��؛R���,A�ew�{�ě+��
|�ث_³����.���DI�':<�����u"qD4.���]�"�_�P1Ә+ v'd�b��ٔ��*�����l�E�wnQ��U��0|t�p�S0��i���#�;i��-!��o/Y�@;��bΣ��Mp.�S)���M�\e�3O���]���<7��>jģ
�QZ}E�ͤ(�B1�[G��!9	������Z�ז&�[G<�a�
���ԯV;�`�LJY�EE���z���������BV[V�j	�tH�JcB��V�_�8�d3���8] ��aS�������,íB�:�o��T�j�-�* >6d�����w�ˋ;!�ͯ=�N(�'����� ݑ�jxxh�hW��|��0ޤ�a���U�.�$-���*��>,9��-j�k�����}�5[�$����>��./���ٰyR&�F�H��=�Q�W�T
�Z��8��q�ߒź*��[l�=�%JH�@���[��1R4�o֡�zN�!��N	�x���{��t�C8�q��l{�;�iTS+۫��d<��F�У�I2YqaxWñ��ߗ�=7~o{��\���6H67���m��T���\�#��&���ȏE�꨸���:@��n�n��\^���_���G·]���x���E
!Y]� ~�pv�MA[�@B�r2��sB��A0j؃�g�a{�q���XbCz����}`���]�l!��UD������7��ĕ���k���c�`@�/5��|����0��y�*V��um+�DkyI��r�h�R_��R�6o ���|�����:F��T�߰;�����:�����M��\�����`1z�����'�T�V�j�6��g��z��T�S7�NZ��o-A,�l5`�!��Zs�7��(�#��{���^8��O�0+/{z�I�y&����������񩼪$�K��[DF_h���8Ns� �~;��}�7\�kU�!@΂�w�m���~��(�c�<0�q�]	ߪ��0!����y'��fɔ'���ί`VE $%�����Z�{��2��w~��%��$e�I�b!�- �m�9���(u%ՇXv;�o��w�;ʄ;U��є	8����q��w�6�~Lo~�|����<�Jk~t���PoP��$0릕��S;#�d���l)���*a�_�_F�PD�SҎ�ZN�ؗ�=ߜ!��ľrFQ\��_���7x�/�%�<Te��,�O5�~b�}��N#攑�["����I���C��f^qs�.�=U|q��`�J/,�����Z�?|Q����QMc8r:�I�e�����Y��.����]�B�v�,���R�Q"�Fݗ-�}�׭O�����3�)iK���abP��bg$�7e�n�$�����Q�K ��a�DrQz���>	��o�D�04���c5��F��q�q��Deo�3�8��O.�[���5\�����m	�?"y��:�Jɶ%L��q楴���b�4Dݾq.>X��7~w�bf��֖�t��C;Ǎ��������S{׍S E��dз�Yϕf~qdI8_,ǅ�J1��$�X�{�aY����b\�A��Oiss�T�i���[^���Q���8�4����|9e-�
Y�	����Z������8��+�$����ǟR�s��}j�?�K��,(�
�ϴwI�7��'�%>�s�x	%x���P�t����7bQ x��6o�^l��c�^��3G7�ܣ��2��Ȝa�����"�aR^�^ZƯ���������x�V;��*zF�YBN4b@i�ZD?1��_b���r��!w��6���V�N5�ɹ��UTO^@~�8ѶV$*&�(H=���}	�=Mi�)j�B��1�!��+OK�2U�JG,�[��E���w�ۆכXRQI P��XDnOOk�B�GΉ%CC�V��7�!f��ը��Y���p��j��d`ESM�5��>��Oԛ@�mB�<u���Z�I(�Gk5�t3�t��h�eW˾������cP�`�����KK�`�S�uSe} ���m�
��U`Gh�b��H��}���&��$��՞�bi8�J7��r��}_�F~����$�G�*Vb����`�Y�Q� �P�j`�ixl%���*L�R$}Bn%�G't�"��]��g8H`�+���i������?��N�̉�Q�e�l�ik:�7�K�W��Q�>���T�P�����k���kj]�ܘ6B�挋�y�o#�-��k�ż���Wܪ|�Mdƕ�����ӈ^�L� 4.%1������dx�Ӫ�2	�]%8�LJ�\N��pQ�a�P=���,<�i�`��W���GLO1�&�j�B_�	,'���w:�,�g��a� z!��c39�u#NA��6I$�47q�lGj��W��K�-�[�r�$2�"ك��c$��K�9i'������\���f���h�a�|{Eb��������5�/t[�����:��=?��ϝz��\s�\��f�ͽ��)m�'���/o�/ch!y�ެ�
.#^hb6��.E��)P!0����1��=�}��|*��OCE��8's��})0�Y�KI���`3nkի2���Aפ�=��73�����>D�&U7G���P�"�V�����d~E���C��g/;S�n{$����r��n��f���,Z�ZE�fe��u�b�G�G�SHg��
r��&�A}q]��Ѹf��?7�#x���C ֚�bQ�~H�C�S�T���.l��Y�L,=4ƚ���D��/Qr��_LyQ�����N�N������ۯ�*�H��{ti���Ә�� -���ntb�s�@��t��=�'�<ޅ%�z�����vP��� ɨu�H��4�t�f��zG'@�����}G���+�0e)�۝�������Y�o-L=R��$a��i��x܈4C��w�&��@���{@�����r�CX�H�^�=�x�O3�؃8���{+�(���'@�,.���;����M�v��9ۭ�J���D�0;�����H"0�gA�v�{4uvI����A�l2m�'�c|� 0D>�S4w%�m���Z:��"���*k�o�s(����yx��*R�!�zy��l�bG#��v�������K�O�2��*Zɕ8e��� ��
.x��*_5a<r�b�$�.�;���G�8�G!$�<3�*F)E�&i�4k!v_����v�6��9b����}�dQ�0��������D���ʹ�L�-$�\ ���X�CJ��x�]����$�s2�����[��#@���@���9��ȇ�z�)�C�1\���L>(@���/S\Ɖ Pֈ��]$�RǷ������]M�#�nj7F۽ ��f�\)@:z��P�,w��Β&�o�	�������b��
���mőS��z���P��V���:��.S�2�����
���X�E���;��'�ތ�Q������BI�nH��C��N�����s��G^w5շ����/����L�ڇ�~x�De>���J.��ZH�N��=�0U�)�%-�)|�A��}���Jj����D��[ q h��3�C3�a�6��tG��'�T�;�h���bi�nP!u*��?�E*�a⮦_�wЧ?����>�f�,�T�6P�l)G��ILw>��}���-�TZzɆ�s�ք��˅u%�UK���7�*}[��L�y����2����xSD��@br�]��\���eK��4u�y�Uâ8J�=si#y$'I i��˖#�-8�r�����t��m��) ���+�M��i��n�l�g��;�j^~
ˋ ��pk��A��m�W�·�O��&d�7�
:�`�|4�F�e�@z���d�`v���9��oi�wa,h�w���`Q�<�O�5�Q�,���D?�+�LU�Ä���&6�:���c�a*R�,�ac8�3Gy���+�N����(I<0c	����.��P2�ru6B�u5^�ku��7�F����d����j����8���9vI-V�.���Q��s��UiF 
�اe;îy��[,CF�HC����
�U�7��������	�X�F��1w7_�@ʑ1��x>��j��@c��bI�*��\���cFB���=�9o�5���BOM-o�b�'��[B��K�7��yQ�IѮܭ�C���#� ���/�k$�1#�|>�x�ITX��U0��:���d ����`�/��H;BaЬ��0�Y�2�� i�|��3�J��D����}]�+���"����d�q���2���&�/�#<�"�#�v[��;
^XɆ�&�)
։Ml@6�+�7�����3����a1�9���O�;V�?ܺI�4��u�s�7�<�f�"Ry�ܔ��{�$�^��ܖr�Ze6�Q��TҞ����b�T�]����8ɘ�s]G��l3�FNh�N\ �w���3��Ãݹ�&Yϝ�z�Y,MBwa���ȳg�<���x�m���%��޷ցw��s$U�E�w�MG�-�ӊ�cK���cV^�j�N�Ɇ9�@EN+��r��)�Dt����Y[$��(�pHH����i��/���B�/a*�ց `�j��S����Y�e/�q�;gm��c�Py	���=&���5E�G����bW3�%.��<P��c��ȋp�
hI��}�O������}پ��
��*�G���l���j �xx0p5J0���� n���XsjA>��ep��z��2�'��+�_K����>2Ȩ��W3�_Ac��T�D���P�Qvz!�Lu�/����O�G$��㖥�g���� �P�Z�&�ck��M՛}����kO�~1|��`�~7� ykq�$�M��썲őd
��9�S�f�@�L���
F>�Ipb,���-��C��^����6�+���؃���'��>��a���2X�>�q�J��ԑ=���.�� ��侨'��HY2�Rct��yO6�6e�̇R3u@w�����5<���֡}�V2oC�E�����(ߪ�+�-����Q���%�a4�`U���S�g��N� R5�OS�W�42��t��t��}�	)P��E�aZ�c��@�%���ʜw�(Ňc�T�py"�pH�ݞB����ӭ�f�5�D�>IY���1="3�{�r���p�;�`�{�.�vne�w}>Ƹ�y�oM�e�ϝ�4�<R�2�c"�@�C�����Y���]���Fۤ��.�cU���� �>?j-H��)�>�*	#@� ��ʾD�"�H����E�[*���k�Q�ŋ��N�`9��9�Z�Sw"b�3�,zJ�>���8�$�y,sʌ�.�d�5jz�� x���iٯ���U�a6�
 �$2��##�0�#�M�W��՜h� ���S%mD{3z��6蓜J��L!L��]g�eE�ڨ�-Wr�s�Gt�ކ��7��>{��?ʾT9w��3o|��k�R�P/[�� 4"������ǩ*ᬼ���,��-t��U�p�E��������}�o�D���{Z�c��|�}��#EP!3�9ȥC��GH�{���~���ŜV{P��X�Ck'9y>� �����]޴�a�k����v+ʿ���:(4�R(3�]��e�ȶQ���e�[	ym�u�u�c;�徚��W�U�;�`���L�W̷�6�P�z��Nm9�E�m�:�[��"da���qOJI7�'�bÝ�L�A��X�cZ��
P�'>#� ��d���2����f����J4����g:�rᲜ�;����f���"�>�gw�����>�h��E��"@�V���ّ.�ʘ^l��3�쁯�1x�����a#^�le~��3��ˋǾ�;i
ot�-u� �-��y|��j�Qe�.J �u �!ܸ����9�(�Q��:N�N�x|�A�A��N/
��6\��xΕ�д_�q���h��~^�+c(�,k|���eT��r�濿��V��	��|���n��W���/��{i".)O��X��^���b&3�V
��>��`�E}��WY!i�<ڵ �t�rS�܈�~`Y��]���H�!��&��+��t����9b��4[)��s�*�����>�; ;'D��؊4`k�$�w[Lv~��C;��D���ӝ��ᄜdH�n%[z�#F�|�v��[�"��S\�&ˀ;4�Y��;ނat��[��g���z�N�艸8�x9��[�<U�����1���Ƽ��0�c>I������V���p�<TܐCu��7���=�(�	/'?�=8��h�c�s&
/�i�Awsǌ�﵁�:�!Q��d�X+�۪Y���i��vn���w#93��3�V�/�>a���Vh�!J�a�f�h��\	��)ft*�Q�H�9j�L��`̖^�/'����M���$�S2f]Xb&�d����� ?jo�A�<�yL�$뜒n��!�s�����1�	�`��"�o�M�˫/%.��޺&	�b��qߣ�A2ٴ>�H��R����o[@+3S�1�^�g�#AMJfl#�$�3�D��PQ� �:i���ff�>�-���'=������H@�B�A��q얉����n_1�JCܓ�غ)��-�o�:A*ڈ��в�N֙�Fs��ډwN1!�26-4�R�%�,����'�J ���i�e{��b�*D@�����>�!p=%��T��:��8�u�d7X���J-�ڡ.X=�d�����%�c��|��4�F��n�QtA��3��	u���֯�r�-��/D���y��J�/3 �r�Va*�^f����U�����e�-i��q�u��{�#�����m?���B��f
ދ��^��������X��Y��h��^2�̀b)8��x�g�|�|��ږ��Z�g�+jc���yJ^28�#T�t+x�N\sg+%�=��#YUPoX�u_�b��Vy2٨F�̔y� �И�Ha��n�9ƪ�A���x.��` ~( PfP����gl����Rڧ��j�Y϶@�n�wAi��'6B�L���8��k��.������e��F�~NE%a�&��fF>��aX�]�R���"���$�p����I���>V����ӟ��X�o�y)� � 1�~��(d��ywP�B.�J��_���6�WeLZZJ��9W��A����ȰD��,�)�`^W�D��~h��4.�%Bݤ�Qk_�>zHg�$O����'�:�A���?*-ˬ��G�H6ɯo$���r���Y��U:F$5T�{���b�)[�|u�O�=7<-��+�,h���X`�>N�K�Pꓲ|�O���.�7�`��G~qTk����"@脯MPs�WV���h�6)�b�'!Dޑ������Pw���bj6m�f�	:���KQ��>5R�����H|]+gO��1f�~�i�O�,��k=B��鼽�Kp7ة@�M]m��q}/�
y=��7$�4�,.~AmH_ �S��ϿZ7+c�-�h�Tc�E�>qB����1Y�������e���5WH��0i�/`����{�r*� ����y�J�}����)��杈�~�оǨ�����ʃe��ë�c���$������D�����������@�3X-���z�;d���x �G��49~�Ӭ��g"g�D��L,�J��!��'l(�e�g�K��:�E
ϲ �j09��N�W����M�:G�+j�����}�n�ws��5�,Z�
�n4�=��������b�t�@-��&�:H��Ay��ёZv�P=���-@q�\��8�fGp�E0��gi~�q�����\5��T`�:6vK�Q/Q�g�q���h�5Υ���95@r�5g倍:�;x�K�&dp&[��cB���!�������Ǫ/x�.n���H�\^eғ�D��q�X��,(f*��� ����a���YRZ�A4^ň�a��D�D�\��H������Õ�L 	�(5>'�c�c�ɨh�mz��k��@���Θ���y�<g��(��_��V`�����1X��w�����ְ�F��_h`]dya
�]������}��d��/�m��hj��YzLɎE�;�QsgT��BA^�ΞX��0�����N�ŧ4{�����}���gSH%(���|ʾ�)�-Z�(9����Е�C��q'�з���e-M��Ҋ�J��n��\����B�`����VGa�{��;���,dt�$L�D�G��	B�V�ẖ��)��,W�o
p���e�Ae���GV�%Q��g���w��6�,r8�Kq1L�ϧ�:���ӥl�R3�� ��hA�O��8��D����^�-h�]'��ˏ�(�T)J�h�:�[{4*K�ċ���ބ�"���򪏘e"����=�/O�$%JK�G�1/F)O��9i	v!X�=����Iq�"�`1�H�_�/`͂��ع�̚#�#�c%��&�>+��+�W~ �ߧ�2���E*uf�N�ex ��;a4����kc�`�|=�.�!0qQ��+�8跕��K?��	L؀dA�}Ё�LK��d_��UT5���?�Ш��¤��A�Mv"�u5��%9���l�����^s��M�tHIq?�gZ���zXbK�k�f jͮr�gw��Q�E�C��PR0��Nju�������P�8.؀�
��6.U��RV�}�3����Ҹ'q%Nϛ�|�)^��O��nU4�*Sm0�z����tĦ�&��f�,��b�픕y(�*�
���i���QI2r��C�C�������="���BZ���ԓ��	Kh�k4R�3�p_�U�-��>�i�;`�9��?�����J��QFe� 9B� ����(}&��7%�,�m]-�6�|�x�K}�P�{0)K?����O~D]w������,�щķT��ַU$~���JD����m�ل��,�C��O�|���������n9�?V��zYlߋ�d�I��vX��R����#n.���4̸ ��]����E�#�,�r���Ӷ��f��A�αP�V�����al��p�,q;�X���e�SvQ��{��)��j��|����P[uG��-D�� ���I�N���L�^j��;�?�����~���3����rt��8�B���!E%�1Q����{�"����b�̮VIA	�B�Wm֗�e5 !��3+���S�T;(��m��>w�g�U�,����"�b�A����r����04��kH+O���.j�h�i;�n�S���E�m�&�T����oN����l�Ǒr��m������8��!�~Ze�|sR���1�y8�?�B��Sn��cq�᜻�\���K�@�$�Kz_�B����3������;'I���ژ�;b��}މ�u�}y�d ���^��:7^�v4u�c���O	�M�<�'�#���]2K6����A�����&�'�@���,��#8�_ھ�GPWed�h�C�
Vvv���U�pA|a�[�.2��v-Z{��Ub�CE��p�􏠙��s`�K�[cܕ)��篁)G3-R��ъ�1�>Wy�l5V�U��:��Z�WL!��y�b��әd�w07����3���@+s-�]��
 ��Q(#�V�q����$6��c����擻V�P�g7��7��ߴ���=L&<�؏V�/!xDԁ^I�E���)��"~!�85-���|�)����[s��/Ys@悥�-۲��S�App���1[ M�R��l�7��!B}"3�R�|a�!�s�1pG>�ev}��:t�
O㥵��cۓ�܎wHt�K{�ve�|fʽ �s6!�ی�Q.�O����VdV�I���<��VU]����<Ȅ-�[���tv\����	�ZWS���t]�W�� � ����e��׎z)�Z2Ă>e)ܹθ�rV)R�z�z�8�o�=Br�7$ø{9Ц��M۞�Td��wŶT��A��r�J.��QJ�� c�H���S�2��Mz�6qX�Rt��(RW�� _���-�;5���p���Ә���?���� ����"2��J������+��l��)p=U`������,���4����7��+�O��w6X���	�������L�'�x*AزY%�/�iږ�8f�:)��h�j��LW��b����mQ��p`%�u��*�0�&�f��w��K�g�WxƦ����qs1ɧDdRG@;��K<8<<���^TYy���I[p�XJ��z�4>#qT���QGq,���x��a#^�Nc��6�9 J.���̯}2�Vұ�J�o�=�i6���0�@b2%��"�$���>�<�m�ԁ���ۇ��|��-~�>�պ�j!b��H��2��O�y�oP�g�7�T���{7EP��Z��<a�o�\���n���?d|� ��+y�E����R]�X]�K�-�`����ϩ�%�YH��4r���������G�*Q�d^�䜚��꺤=
�����fKOi�[H?������m7��Lh�3�K�7/h�5�6\\���^sxĆO�V��� �Dm�DV� �a˞:Z��Gts�E.^�R��]φ��W��*���d߀@i�|�BƢ�T�q��.��Ҋc�	����Ue)�@�p�;rQks�*(hՄ��d]�B?��R����z >HLV�G�R�f�w/�鎾�&�4hF�w[���b�-�dX�:��煖/X�����}�4c��&=��]̪�lX_cO�8�Lг�6�_ �%�8�I�$��á�C .�IL��`!]�f��P�2E�&�f��cO�7���[�Y�'�#n��(=�^�%��y�lhD+:�b�hl�Cx`e�Y����}]�TI"�O����Z�ψ�H}́X�B��T�9�h	����7�B�<EB�.�;m�gV`��oy���A�����&*���E�>�p�S׈j�p�r�����Me�B��l�i�Y�A����6_g�q���XA��G^{D\]��]��k=IE�W���Zf9mإ�$u'�c�1ԡ*�����Jҳ,(9��=�1��u��0��;�:�#�sf�4��W���d_�v�Jr�q��=2NƩOEiV�F{g�*H+�IVz��0���#�b8�4�!��XՀl^H���L��ZU��7���p�_T��#�#[��]������Ӳ���d��Q��M�S�7��[�nuk������s5T�3h�O�3�M�D��Sl�:`�AS��v2��)bg��H��νv�5gE�b�G����p)�R�{�A���B9�g�3�-��oq������D�}�n<�@��eE]�ʑ�}��YX�Z �U���3b/llfpLG�R�2r��ޑ"��B3�K��/
��Q��5vq� ���������KQ:��kB	���&��L��6v��/}.ڧ���i�I��n�v�z���D�}E����W��R!��%������bl>4K����3����=04[ƻ؟p������9,������"6].}F(U38�.Q�{��P4�-=���c8��9�P?q	De08��#��|���U2Gމ-��)�Lq^������I�_ɖ`��l��`�ź��,�mܐcB,��D���kf0V���Q�3Jh*tC�_�N�ِSqP�?2�����j��A|,��;}X�C1�h�������эb�(�_�z�)��v����6B�:�V�]O�E#�1t� �Nq.z��E�V��ԂB3����VW�$rq<�t����onO���7:�r���.�lӣj�Sl�7h�њ����ikn�~k3D�zѽ�v�HZ�A&Q�/ƓH��@���pl����D���,b/,-���8эnN��3��J����EЪ�F��2Q�PP�{������ѶF��r�oݹ:kp����(ɪ%S169_>y�ϫ���m�[g�S0��<�B�莪\��9o��-*Ll���p�($̑��-����Yo��8��8^��HQ���(f&���� �^^_����U� �	���̯@���}S�S���)�F���U�P�$�rf�U`J6�n�ʜ呆��+�*�{| 0B���F��4�9��9�+�2o�7�:��k���d��SȄIe��@W�e�Y��y������+�XU/y�����}�k?.EE�&-��˸%,��+o��E�YTk��eןO'�9<��]����%�w���{/���q6���	�����F���\�ŕ�T;�,��&��y䕜�/� �0S�
�ę3i��������wӒ(��k�����uoI���!�5��lk�Q����3�V[=طk���sOfb�qȶ6��l�^˙�m ���~��%LJ뚦۴�Չ�qz������0�R����O���Y�F�D�Ź@q��l����Buᵩ��7v0��w]Z��ʼ�0�f��4�B"`t3�$�y�68����2��H��-4y��0��4��6��K�C��0HL��h%m`WxIJO)J�¨c�"��U��}����[�A�Gǫn�k�kX�=�Z�D�������L��J#U(��n��_
�ا8b�B��=�
ɱmH8\5��!�c� ��%�%���9dLE��pt}+ޠ�z����+����ngH/^_&���L�}��𵁽-q���"��j�#��y�.���d�N\��g���%M-��ٶHke(��o��.CRL�k]��6�/�G'�GL�HD���v �;wF�@�O���&L��Fy�x��m�[4�b�䢨�Ы��������vo�*���L�>���2�$HeJ�m[`,D#n7�L�'V������d+ǉyi\�C8W�]!�\.<�x~(B�׆�9u�?n#�T�ړ��sO<z�_1agn�����o�CҚ���v�A'e��ø�����e�l���R(M��I&��z�MP���fl��
y{�^��}�0=w�AHU�,+� *HZ��9!��*wx��$��7ej�	K��X�*T)
(����l�M�.��y4[�]��*	c����� �}��B�C�w��`�7Bh۷�2�:�=Ne�Hk
��1-��y64�9D_�@�92j��2hy�߷O4o���6V�U��F{m���;�������B>�@��?w��#_���O�N �Nl�УA��6��8�8C���4ԧ��s�@���F#:u�tP~$��[*�u�#:ͤh���c�K��>�V�~M��*?�!���Eñi������~�G��{D�'�.�!�<�fn�N�6�h�n�>�Li��@���-��Ϣ�2��D>9թ��ά�(e�q��X�6�L!��7$� *�{�1�x�0WL�U��"��^*�P��8rv,����<��[UWO�����-JUu����A<m�MH�!n��3���߇w���q���l�����lw������cSS@�m{�uLQ��<n�ln}��������[%<>E �v�k��~�5CYMր�>)���Q+_�T�b���E}
Ai&��I����%d�JcX��QG�Ta�����<ŭ���Z�����2uQ�k�z?4ݤ,F���)�tno*��/�}��{L��|�}�T�І�0[Ǯ�d�	W��z�n6��x�%�bl=!����{�}{�v�NX1�F}0F�Ƞ��|?��U�PkF͗�U+�J?h��8��W����|�����Gɮ���.�ӈ��� ��_l ���m.�$��]�-a�_�#��*+Q�4���>�d��sp�Kq�K�^����{Yel�b��c�Q��ʿ_�#`���T]��ɲPS`��]���f�yi�r.(�։�b�5��jT�U��˶�	y�Lw4{Bl���R1���8I&�c���'�������m��<W��R���B��C�������hn�I<����f����y*T8��+KA�CV|T�W���sA�LY��a+KuJ[��
F���m��ª��4Q�[�h9�0��V�qI��[7;n�k=�P���0,4��^�6;;8݃����Wl1|��h峤-2�?Qa��dX�&�7�,�p�P'�H��;b��S�?�T-/i�������^}��s����B{2"}�Q��~ՠ;�)e�%�]X��(�v���� b��
y�:wW-f�=��V ��#�#;mpm^���˃�B�3���D���Y����uz�����Ib���cN��Rf5�#�pf̧�s�6�����\�
���Ō�#�n��еK+�]Z�9I��z�zW|ո01��˟ L��}]���70;]b�xf��F�JU�1�D�i�U�g�)�_���~��-d�=����L�̼�t�o�}v���).�� �ܠ�4�N'mi�)�ڮ~[=��3lq�B��L_.Z��'j�d�\K��Q�Ll�|zM�"�X�a��ڍŨ�V�Ɗ���p�õ���;�Mݏ���r�/��=Å*R+�J\v�I�7������;�䐁 �zY8�r��.�(�����J���D��?j�L�`���Y)[c[�����=j������9�O�E������y��y1Ø��8��Wc�� O������@�lsQa&� X��� ���f���r�����NӶ�te�p_�g�� �K��<1?$�q�x��xK���e�%��Q,D���*�̏�w���ыJ��ge\k�c6��(�uh=Q���D� I�L؁��:t�<,�`��!*UA����`�HMA��飶� ����V�68�%���?/���D�n��n�_�kg�>�
�(��̤%ؤ6�[�#Ʀ�A��N�'�r�k�D�ڝ����y���n�j`T,�>/8��MH�@dJD��C)�|��`�~8��]�Byl�}�4��/H�݇TKyi1|�|�ǖ|�}5�J��X�*�$����w���QB�\	��IQ�i� J@�Ŵ�/'r��#�xUYk!3õ�\|W��x6"N\F!Q���C�0�`�RE�S.Q6����}�$p�7�n�ĞJӡ@b{�k6���[�K��$�̽.��e�?H�?�:G�e���5�/������T<�u[x��O�2mjv�����Lߚ(����#��n�0���Gxl�� Mc�#H8�?�>�F�yt�n�����D�Ǖ2�7/vxcn�cv�]'@����i��+��^9��]�=O���A�6�56IK�lsHH{梶a\�+��6�X���Oh����Άa����y���|�䧱�b�,s�1��4�Tt�W[�4��-�U��+P0�����p�$�g�M�8��痷�Ŕn8�q�>�O)́7yb3�a�S��M^�!Ŝ����h�k�X|��1��x"7�ȕjZ�*�����j��l���ػ�;�`�P��g����b����t��8�$ӳW��EeR�����$�u��?�uP㾍o����z�F]U�� ��|��k�Zx�ҩ�r��nK,~sI��T�X�
^�@H�@:
U3lpR�\|If����e�]\��V�b$�D`Jz:��g7,��^]��)'xh�]"Ҝ�9!���-HiJ���K��l���~i����\h��&kUa�6|b�T�{�q1ؼ�Ħ����%�z�	t+N���L�����3��O��H0~�Z޳RڍD��څK��e�^`�غ��y�p(9gz��e�~	\��в��_F�e���U� .5b�� �h`��?k��iv�8��:�h�*��z9A�[2��x y3�S�V�$V�Ͳ�z)�����*�9$���t���E�:�k�O,u�B�=��?�=h��)��U����q,����.6C���5�Cm��BNW+��#T�U�ѱV=އ=1�>���q#�<�Փ��v�9�ӏ'��t�8����ܝ,pw�'<0�(F=%��"�����-La	\�d��9��;
�{؋�R�5��J��� `��H���|��/#u6#d��V�6�D��$G��B���ֲ�hԍvީ�G�9o*��b��4���B���n�ڳE�Y ~-M��� m޻�Ea�6߃} }�|.��N����Z:��g��Yu��nCN��~����/��Rg����� ������G��	������wW,��(e^HY��d�P<hG��`���@S=�@9uk��v���^����
��G����8���"����y(V��
]��x�2n��QB!�e�]�/[�I�(�U)�Ay�8��ы��7U�,�ݎ�cM�����g�@���'��ڏ	x�!e��d{�t�XضC�����T��@A�ߨz�ʿ�Ҭ���֮�{�3%؏�%ǻ��.�P4J�����c@�p(o h䥋��ڶ*i����9SS��^L��d�C�M���;Ԟ!�
���'�B�%����|���GƩ�=V^�Pzx́��\`�A�^h~2�]�]�]�]u�(P�I��j<w$2;��ө�[t${��L��i�c+
oP���\�1�~����Y~�ɫpZ��[V�W܌p��B�lX9�3k������2������4{ϝ��&�t��T�)��d���^N��Қf����r�a�/��;a���O��o�é%hV[�@0�ܭ)�㒒����%8���+��;����7��������߇ M\=�����AN��) %�Xs9+=�i���\K�Y\�~���Al#�+�n��#I ],a�L��قc���C��~U�^.S��:�k/R1�����|�	zS��\����l`�(�A��ۜԀÁ ��Q-��j2�7&ϹS�a�M�R\��)Z�<U�w��&ۜϻ��b6[�;��ƙϺA�F(�UR�&"uH �A,p���B�sq:�hX����Xm�>Z�F��'Ns+�B�sy�L�f����!����l��ە�3?���a�j��جL�c�-Gu��#+����p�>��[s`��E�kBG�{=d�-�?�����j�?�ox�q���|�t�s��dU+�8�I�of?_Ab���x��` ]&�*��Dz���&����_��C���G{ж)��@\垬]X�h1]�L��#r��ɰ������U���O7�v�9�ţ��*��n:9�X�B���LAzR4A�6���,�N8ı�=��d�#p
Y3�q��g�&>�v���{�u˦3��4�A[Y��9؃5v��|���S,�v^a��G-
�]�_�Cc��R4���!��Ҙ懀� ��)Jj�3����$��R 
��\�d�X?��5�9�3�Ԝ(̼2��K'q�+�8������f�G��1t��\2:t9X��yc��k-2�W\��_�zPtC�<��@$%�4�������?���!�P�����Ԧ����Y��'�7��Et����j<̩��y�=��*̼��3�g��e2RZ��q�ˌ��%��m��#�׎˜�Y��H�&�Wm�w&�+����iW���1vZ��v�'��ּŊ���N���|�ID������ ��ڑP��D��M���o�!_�2dA��L�)��[R����M��x��9N����F׆�/U���"7g�c���9��U�����J �lR� .�d[;�Z?Η�n
�iΆ� ?g�l�KczEPx�u͓	�G�k�Q}On�aV����ݛK�O�ce�ӯ�{�<F�6|os[%��o���1��I*���1D�c�� -%�o�Mb^���شi����̘�5�U� K*����� |��B�)3�9d�q��!\e˨/����KN����Ez��>���yg�f_�Do&=+Tzؒp���?���ȆK�C%�#y�,��Q 8�����̇��������}s����N��л$7%�oNt?ev��M˖)Sv�,��#�z��{y�ѨR�?=y����|�ʷW����.�*��?�e�
WuCl"gw���3�~H�v�~N2�:�R%m�4��ʡ\���g�$�Rk^�&1��?P�����������M�({�x���_�qݔ{���5�|.}�R�I5�_���hی���K�ube��>�t���e�?"���,L��
.`..O+R�x�f����(I!��J1x�0�6��`�P�-1���=����� >yz�X
��E�Ĝ���6O�q�i�q���7f�[��h��p����c)Nӆ\�!�/�*X��b~��f���#�׏*	FS)�v���a��?�*�p�ڂP'�g�v^T�(��I'�؉i��%u-��$Sޅ/�% R]-HV� E���ʟtzҶ>���>���X�.)�|�a���νz�rv ���}Bs�C�¾�r����#Gd���0,�t�u��_IJ�������/Xv��[���zv6C�&�Cf�+8�G�]��#�^��
�e�>$�$5 � &�<�N�-b�Nt�8Oz0M	p5��Ǣ�� �6��="+�x7+� D�_ѱz;����xF��yM�����-$���,涛�<���چp���e�iW����M�#@!Pn������gg��T�&�y��J�an���]�*l��D��� �.G8F}{2��V���ar�h
�kD���{;3}��0b36ҮAd��}n��$ro����S9 %���")o>Q/p�ﺸ���\'4�Xd�����Uh9{��&�K����&І҈>�k�*����t��&��A�]�ѿ��S�S�^t�I%�|�]:Ǝ�1V�\`��9��k%�+�Ȏ�i9֤�0���4?o �/�3u�
ȺQ6%z��ÿ+�w2�¶��5��#P�㏵
�����^^e�3EKc�\��d{L�:Y�����dl��O?R�?FUr�$���S���Y%"t!��91��u?���3?�&[�B��ɢ�Ԧ�	͡��a|7�����+��ܮA����o\(d�25�r�(��+��'�4:��H}v�c��j�N�8?s�;�4�>^���g%l����E����$V�#�r���Lx<������]:v��j���峸M�\���;;-�������m�id���PG�&_�M!6�Bѕ����JlHG��������o�ƴn��P���xy���0�t�+Z��kti�ћɒr�l�ɏ�±G�=��>���K?|7�C�IȌ�����v(������ �H���jhPv��C'�x���
(Mn`�,����f^M�����Y\?�����	��8C�`�VwA�3�
qP] �iV() ��^�A�E	�U�U�Yo՞(���X���G�'v\��oe�F�C϶p��QF�[��5�=�YP��aE�Մ$Ѕ��"�P����993��V����e��-j�ﺈս�y�vj͇� �V�&"a�<�
6�� ��~��I��1�kd%������v
�� |ዖB��7�
��<(6	G,"����	�O�Ϋ��9x�I"�٦�Z	o��$�g�e�Mz��B�G��M�k@���}����|L$I*���eK�������Pj"����R���KB���	w���s$H'l4��5�|������T��9W���[�C�9��%��:+��.�D��=��:��xm�Ǵ�!ލc��<V�a캄Mg}@�f�`�����]J��Iۿnb��̤�I�lI��[Fν��&bJ�pb~i�چm.9`W�-�����5ƘR��%Ϡ�����6e��n�u��	�X71Y�f�)�0�V�N�����y�w�	�}a[���4���.����>ԕj���o�� Z�����+n��ě�o�9����B1G ?9�g��`� ��9r�p�/�����	�*:&7�ۜ>��sD$��r��h��a����[6TT�ѫ�C�h�	�����
�4w!>8Xc'��:i��	�_q��~��k�Zr7����r-l���сՁwV��?���>|o�4}�ZT��%���N�R���'82Ti3�̊2���HT�sFR���V�TZv�7�v�i(˿��mI:�����X�������DlE�q����}�u����D�%��'�.��� 2�X6�= ���CQPe甞5ѢQyZ�>��6���&�fJ���E�sU�I&��,�M��X�e�<
���W�wF4�N�{�Jp!HY�����	Ȑ�ǣx�p$�w��a��G�Qu���5��5E��q>b��v�XRd��XGPqU�ta@�4o�������r-�}?���RQ�ԙ[�ҖE�c!��^��ˆ���-Oe�4 ��xl��>���a��>��#����E����4�E����Q/9r�bI�}���L��-2�`X����,�oб���S�*~`��.����MW�����\��dDg]ov���2a�D�<��C0�l�͓5� �آ�W�<�B��xb`����:�8���t�y��ܞ�����Z�}��g�����U�AL���nf�)�#�
��^���I#W��7�I?M�������Y���ڥ� ����N�>i?���K������5%c�p=��0F0n�0��%D0��TX�|��ꗮZ
/t���~:���g��B������n����`�5\8T��Lhw� �(ov��Ib�Q���~ɮ4��}�sxz�H�~`���W3-Ly}�tG�w˽O���������Ԟ���9i��u�bD6<I�G�@���\�*��l��՝L4����A�<�:���+������m����mUt��Nr�ˏь��� Y��#����yā���`u��D7́u�$vW69�m�D���%�f���-Ͻ,W!@`J����^�^R<p5���w����z�K�#6��
E��Qԝ�����LE�7�8��˳O�%�+���P�%��~\�,�>����E��	bE�ч�Q��+k-�[>�(�Cpt�g���=?�U����u3�ʗ��ǅ�($�qM��EV �<���=C�o��:��%g+�>�Q�\۠��$���r�%K{6&�ιM�A����o?�{.��=�z����?�h@��I��9�����E���:P��&G�nO���Y�n����������t)V99N�s!���}=�f�mWaS�"�����SLNTٽy����]�Y�ҥS�9���q�tI�k�r�Q��UJs����3vxy����)���'OʄB��l�;_��' 1�׉Et�<Ɲ��2�P|�c�C���e�K�b)Re�� ���R�\�Q�*�?����������J���>��{�^CHYY7f��2j?lі��v�N�������ŷ�0q�}�(Ɲ�oUbn�G��;�m�?n��
��%���ԣ� <X���u`���q���n]�P\�;������i`��o0㮎ŏ�Lg�jHt�,Ԃj��U�*���$�V��6�-� Y�϶��K�]_��4��y�U=����iR	3�ſnL��6��p�uZ(������W
7x��|�����d��9�#0~�s�O��ߓ*e���[r�����nH�'t��O�t��%�w�̳C&�f���]fN2s!� ���^i�J��!�x���9����+�:Wa�ޠk��`�N���>��d�*�1���+�ߨH�XO��N~p��� �0��{��0~�N%R�ƺ1�\���
�f��'������Á�]�e٤(E�^O��������.�ܔ�V���&j����>ǀ~�s�:p��/��/EF���9I�K1;��[*��#[�A��R�`yR�2��w�����E�˾�aY"�/z���2�T����:X7�h��-
>��r�G�	�g��$s�o,�՜t�̎u�g��<�W��il��<s�*-��`좻��H����h�����Ȫ	!l���V�u��(,J�k��������J��Eɦ�_nZ��&3���}�o$4��/q]��cP�����,�q$�����AQ�jc!��N���o["��2���࢏����e*��㛨|��/&���b~��0�S�G��;��X]�-EXϦ}�Y�� ��5f~9}]\��W����tV��o�������ۏں����u&���ԙ������&�`�����Q��~�e�����B�/Oe��Gc
�:��a�QT��i�Ν-�K1�<���]������?�'y��"b�,� �6z���F3�����`����nn�X�ӷKrG��w���ܳϵ�OE��ϻ�����A� N#�ASW��UviЇ>Qr��L�Vz,�8�#Dfλ���$P�G��YCq����۸����{$�Tvz���m��&��
��p�<�A��<P�,����VGt!r3�q��xy���}��G5k�j_`7�䅿K�O+��}M��f�<������YR���ƴ൙+��Q����|(ƺ>]HGQ�e��)��������^��,���>�v��"���;cq�Eg�}��,?��Sj���֢�AK��Mh���4���&ON,X(2x,��T&V�i��^EԳmf�D�w5�w�e8N>gba-���	6�[�+�B��(�5�׬���xj�m����f7���5¨a(a�"�UBz��˱�֜��%�J��'_2L���V��=�z6���Z��V#)��=�j_�?Փ��!`���?Y��ă��#�b<��\S��T�j	�!�ց
�ߘ�l���œ?<BYE�A(���-1�*����#��<g��mcm<!���V]�,��Fll	p ��,,m,?�N/_�\<]muO}$�4}\��E�И�����)�I9�5�ՏZZG�]�;�8%m���/�K���5u�� �@�}����eE�$#|UJWy�v�`丧M6	?VD���T6b��/L`���'`��bҎ`Q�c���I\/�£y�x7��%m�$#�hs�5�W��LF7q�������Y�J���0��b�?]ۧ��W�-S�\����[�4"\����i�����?p���U,�u�>����(/]��Ao&V�է��J�{� �e����f/��"��X�%��b�����maE.�����4�?��~���B.���fI1��h�oWz�=�:�1uRn��p[թ����z�X��<О'Ȱ�T��P�]D��N��V�+�j��ck;��e�"s=R���]'�

ja27�)%�>$�~�l3i�U�4�n��1��'"�CvJ���׀�����se���R�Y�z�1��^�O0�똱�xK��Qs~J��Wj	�6EX��00v���o@�d�L�
ǐ�U�M�<�
�y�2�x=�-�r}TQ��e�	�k#O5�&߱��q�v���n7@Oqx�����S`ף�,���5m��	`!:�Q���wބn�a���b���!L6�����dN�D	N�^�4;j
AچV����'�t� >����{1]�����B	`�S��(2K�h������֊�x���̫EF�t�j��	���vd���@�W 6�EJ^۫�PHy��2*M�鈬��?�[Ca�1A*�3eL�
4[=�4ں�7����/�ǰ���䷁t�Ƨ�L�����T���&�FeP]j��4!}:��"��h�H�mpr?�E�L+]e�J@��5��C�#�ز�ᡮ'u3D"�Z������YU�c~����sv&S��ߐ��mbl�D�1��-��﫽�[��JK2�"�X;@���~�5�ݺCӟ��/��7���K�cZ�^2ri�v5>{Yu�C�"���W��A>Ky��fp)�4b��͹3s�W=��4b�4���ڕ����9vU�M�*�\��W��RY1qUQ�r�o0��kP[(���j��B��Po?���ه��&�}:�-��`$D1�5���)�ݰ��4�+�hf ߳<�sw	Ց�6=i�0n��Q�Ʌ�4�>��h�A9�M[M�s`�m1��s���wa�FW(F �CF%^���3��*o ��/&r.��^ƈ(��C���gT!��72/W�a�g�UMD*��s�č2r�P��D������EPYA��t\s�K��	לi���/��+scD� yO{�ɥ_�p�^h���8�-�o&�e:����K=RT+,��2��ܯ���4�1��S����c��Jb`��_�T[`B��S? v�9¶���<�o�����F��P��?��:����f4]��h�.��|���%���"2:�c�������#�1Ц�#y���8�$iw�m��=s�l^�`�/D����ԓ��<h ��R �ȷ�9�}]t�&Nr�����_���[c�u�*p�R}'R�C�)��ak����tњxQ�r�f.��>+Z����𙣮������g��48)=Z�ۄ�(�)�)����x��9xȶK���a^
c~��S0)Wp>�\K'.䔠=_D^n�"���v.�o�4M��0H���,��KD����I�Tyj��N4�	i<?kN,�d���x�J��7q9@��	�0��XԠ��C����q�I]i�?5�X���Er�a�ދ��g,m����r"�0����Qa��/�ja��p��Z%%�m�Cbݚ\�9`!���<�'�z�\n:Z�1|��-V.G#���{-����o*: 3�\R�fK/cxu�+d���W�d�_#	��w�&_�{`�u7Qn�ku��@�[�A��8�pdD0���ȎK�B�c�IJ�%9>�w� &�<U�^��!�3��<�85>r�"�f��S�k��>	��]{�e�m�hY�ஞ�o��@��Ź��aa�ƒ��K�Zš�����CJ��ԭDhE�}*Ǭ�ѳF�b'{!i$]��"�(�����m](-�U��|�,������z�pc�m]Xc|��Iz
j�R�|�5 �m.���v�m�쥥�����K8i#R�dh m)����m�����c�zQN�X���g�ece��v�1�d�3��[��|0��͍,�ܙV(�f��a&ga`�O����NH��H4ֽ�DK=i������$d;Ӛq���@Q���[(��R�QK�qFk��W9�����f#�_�c%+��ݜ�]��(�6��Fa��\��>Z��P����~�*�(ǝ�B��Y�qG��� j+�_��شY)hu�ҚZ���@@o�0������t$�Ԍ#r�~��>-{�����<}�0X���
Q����*y�b�Vj�:&�\��dGvp�Ϣ=�Ji@�#�J���Y�dc{B1���0~�q��Q�S���k��\��P]�E?U��mh��X�>������WS��R^�Vڇ߉%'���_��NaM
��W{�1;�hWT����#��CDO1�f����D�N]u4�ӱ�,�� ~�b*j�3kf��Y8�?�nS�}��r�w������\�xO����O�/�	n�;?���o𝽂9�0q���{���Һ&>!a˺6rh����">�*�n�=ݰX��<[�B�"��ZyY�}ԥ��"״b���g����'!�5y�uw�!&p�+%�v����:d�eSWG3:�-\�RЖ�sE�!=qr��u��l�
��lؙ�k"�F���I�^~؆�X�.A��%e�3�?ǝD�	"C��k}���5厄��$}Ny?l\�4���ϝ1�����x�K�K{l�������g�'l��&�q�Jf3 �n�����)V���9o��g�b4���(��+�õ,�qKxLQh���	���J����e%�6f�\M�����?�а˶ Y�Ua��NL=] �Cn��ɺ�\�ɟ��o�Mɫ8���<��Z������`�o�G���}'a�����f�,�)��C�'6��������`��X�^����i�?�`�|g���kl7��ܣ97��Avk�Q���YU�Y�B{��wv25��^������_z�`�"���[`M_�19�ʓ05"��9�?R���z3�6�[I5�v~�9�mJ��=cC�F����QIxB�8?8R�A�kQ��xډ�yj?*nDG��� �a���srx@�xPw;N�cwT:��MY��[6�pw)B�>���i׿���OsgOf���YODG��A�8ak���Y�)��4A���>��,��f�y�xcB�Z��9�|���Ё\��!�'[�@o�`h-��N���o�� �k7��*�z�"ͱ/כ�ott�w��S&`>r${<=^G��?�~�����Ia\)E/��vw
�FV����2($}�Eq|7��A+~��<̗fٌ�:���U>RIf6%��#B��g�*�������v5}GslUq{���k���y6ĔM���%%A�lf��S7<(��k�_�����\Jc�7����?�؇ې)�G"[�d����b��(@��q��Q�*r+�I��R��2[gNZ��M�Sʢ���J\1�D���iZ/Ɵ�o
�f�p�2zAe���{_"��kSw�$ߋ9V�)k�v6 �hĀ�[g�:���Uްbx��ִ}v��8�eFX~[0�u�ї��O�:�r>�j�U�Gp�܌x
'j����ڒ����.���Rc;�q���l\m�e�7W5�e@��Գ*��H��-�q���&�Uz��,�G~��� �tp&x�f�k���o9-�qT8^D����Β�z���|T��Qש��>�Y��|bӻ�t^q\S�q�r����[D7�v/���.���<@P�Mu��_�x".� �E3�ؠ��S�sC��D�3̕p=17��8���vʷ�~2B<%[�n�KX�}�.`w3�⑂�>d��קN0�hۃ2���# ҋ�,O��0���]���-w� 
W��h���c�9{�����@xz`�06ɫ�\?��Wj���Rܣ9���[M�u&P�e���H��,�b�3�^-�*ak蹸��ٖ��Jq-0I]>��UOV~N���]q�|ʧlዎ7��X��"�%����Q�ަ9�A��P�#���ž�`�0����B8�f�ڞ;3{oQh�,�GSK��ۺ�~�b��Jx�Cd��)��F�tY�����c�{�A�g��8YL�,�3jh�
@�t6����͜{q]�1쿻�<!�@:�)�<��I�<q��Y�[A,7��8���u��Ҽ?vU�5���$%�t�����!�}YDcCWl<æ�1L��y=�c�=d�+U�W�;[1�Eg�\8¦_�D
���=m�N�-����0��sh�4�C��`І�����M��6=3n�o�!��Q~�ؑ���t���̍�of�9蕣�`'A��j?�q���DA����$�T�1�s�y�u�n�50��wT�W�m�D �$�5��\�[����^��A�w1�C�vR���ô��rL�S�a�K1�G�=Y�6�Upb�a����ý��Ovb����ܹ#�X��|��n��|#���]�
�܀�2ɅL��!��9x7C�]���oգl4�]|6Ӟ�h��],b�����|��!�1B3��*6�<�#��<'ě��1���w�s��īM�q��W|�����6═���G�����M{��-d��̮�,��]���CeA�~ph�c �Qͳ�X<�g��N}��_��4����4l \;2�K^������ݤ~S/~�Y ���ԑu���k۴΁6�/_���?��� �+�v��]���;]y�V�א���,���moS A��U1}`r���,1�.�������+F��1�������x�s_�#/б��Jh�Y�%����$Sn�����x�%�,�. Um�{߫�?����78���f��,a� t�9mC�Qӳ,7
��a&�WN�^�U����C�/�o��6λ�5��lM>X�b��������n��)�p�.�l��7�%�G~\�(\���?i��Y֐E���y�����#=�����8a����ᮌw6�t�ǣ�w�p� `�H�w':��$���Z&�PT�i'B\���quV(t���Ċ_�l�A���<	-Ġ�I�WM����^���t�����N�]2�JĞ��s�ɟ�<2['��� �G�
8,�ָ�k�-m/<�/55i���j3)��
�FꂈEH����m�} P[����{(����8z|L��~�^�EY6<l�D��&��X6�+��t`ir!V�AB�����	���h�ݞ�l��⚘�񻑢�^å��N�!\X�U�p~��rK�����TRf��5������= ���!�@�Hw�<&�_�S˩�[��ѷ�И��G�X��*b:�]�KKh�4K��r���┺ V� ��	zz6���4c:�C^�(Z�H��`��2���F�}@l��7�,���"e��JЦ�'�{Iv՛���d�J�S2��o׶�VF��y"�u��e��>^�S���v�#W��� ����ӝ�2]wh�O�q�G)
y��rVuPL�*&{�m+��dB�K�|�V-W��6����܊� Ð?��B���b�;J���fd��E8zZ̻�]lH1���]2�s�b32|�Y���Ӌ��t@�̨o,�8bKp�T�ձ6�5"�9.��
˿L�P�����m��ᜟ-�T��u�N|>K�t�T���9��uy����s�c��/W��%�w�TB��擩�찅�ʉTe��i�ɐ"��gTC�2c ���{̛v��=�Y ��9��L��q>�=J!�����<��f��Y�\0 pךY��E���ƠegEk�Z�W�i��slPO�w�+�2����� ����MC��.�6���P�,�N�CњC�8�\F���/�<B��2�q�w��<ĦIU�o[g�@��   Y�?+L��5�`�S<˖��0Ms�C#~�<�l���Qb�(��2A@�́.��5�OV�PY��h�It�S꾆�E�&�����%<�ń�yڞ:NxO�+�'w��
Y&������j�N�@��h�ʽB��0<ϛ�tMg�G}��]8f:x��3	I��
.�{��բ�aVx�79kР�acoi��5F7@&�qgK{j�
w�.Ѩb.������5�Fw��"�ˢ���Zu%���z슑�6�#%u8�Eh��Ynˊ2��U�n\��þ&�4..Q��-+�����~V!M~|�Y�����T��Y&��]��Ȗ�"Y4�/<΂"�N�5�xQ�L�v�)�a���������d���B	"%�2��lm��FUƽ�����d̮v#ݏ���ax����wYzf}5���@$�A��d�z��*;N��Ԁc~8�m7#^��["i�#��Q�(N.����P�#�:�X����:�-���(�e�_��r
�_��yG{�"K�g
y�>Q�M(�쵙�$��M҂�,�"��X�����o���k�/�r�1�o�>��!k�em�>��[Cu��-�A+��z/��}�
!~�n,��SGBB|�I�����{fu<%�P%2El�����E5�Z(��8�>2����AY����3[���عJv��/�0w�����W���ldN�7_�*9c)O�_�6��D|�	�v���s��`�Ѥ0F07,m6�1�|��@�����{�Vx�聫J����W���!����G��rv�{5�n��|�K���S!ڲ:+�!H�C��Ne-�5�
ZA&+�3
�M�}ܯi�ˇ�,�s�_dv|ؔ��7^�l���姱�S��g����4d����7��nS�[��l�S�h���!�L�H&�Ő�x���$Й\�LW�ef�ʁ1+�`7���n�B�'�O�>*\%�����g��~��[�8�Sp���_/�2"��z�R�P0� e����q��W=�tO����4����>� ]�'�Б;����~T>�j���8�W�z쩉���l~�2�i:�D���C�'i|�נ�[l�G�q<���н�uwNOh�F�2���pxG���ea�w�m$�0e��ڈd��fO�hd��Xk���xC|F��,��'��t����7���X�n��6��_�ЊY�%ZH��ϸ�-@��>+����R�4?6��*G� ���5&�����a�"_�QF3y� ����iOEpE2�m��r�z�&��C_��m��,#&]�SY����\�'���| l��,�x��Y'er��И���W�Ѧ�u��[��4ؠElѠ�{�}卸��Ыpz�l��s�4c��|[a���{��r]ާ�	�K0���!Qw�)1�����2�y!̂M�ƃ4Y⴦�5vJ����0D���?�|�����~���D�F��\#��\]��R��x1�ޅґ	� �� �0ܚm̲ѯ/�l���ыqx1�ygu9ζ9����i : ��~�g�;�����'��y�q�Pt�`tA{��7�D�?�X-�0�6+(�=�F�H��-DC�N�>_�FJ��C�#��:c�N�Y�1����K�-A�^��Qv��}�x�֘�eڍ�1���ho�o�I*f�a�Р��'���aw@�6h�Pٍ�T��_��LP���w��EΖ��﬛d��Ia�u�gU%L\(�	��	���|9\��R���o�l�v��#���Rr����e�9I6D=���*d��J_���2؛Q썦RPF ҸŰ�F}����3E�#=���N���Zf���mL��p�*�J�B����ԘC�r(f���~�[�i���~ƕ�V[˒�uti�דR��/��^2|�L��C�ʫ�c\͛mZ��VI��QjE�z�* �3�݃v@F���(x���8P2��s�>>g8�6|{�<�|ʪ��l�,�Ou��|ft \����p6J�B]'X��t�3#G�־��7m���>���5{�X��T���z��oNN�Z0%x��`y�M/���@hშ��6�vi���V�T==X�������>����@����N�q%��2�VEP���=B���=+��mHQla��]1!p[0��cC�{���Mi� ���Pי�k�����F�_Sb|�����H�h�0���٭WVR�m�d�3P٭�(�T���,�� L&`"��M����>#jgz2��ԏRێ���t`��%�?J�\��4��$@��Pt	�A1�F��0����u�#ʪ�	A�R��v�ъq�hUn�v^ϻ\G/�P��pPT�)a>f&�GPPZ��M������)�\����[��؍����UՒ��$�{2���T��6tE�Z�q	;���z�.���	����Z��{�1J�hC�|=m\�O. ��+
1�u���R�f���N}��_���F��zH #����V�K��K�9!��g�xݷ�f��4����	e�cN~\tlN�h�-/�{��g��S.⩔�rCp�}�L��y��Ss�W�p��U�61�MS�)����b���tҐ$�ܸi���j�_Z��2Y�Q��
�ZtO8��TG��GɁր���@]SԊC8).U$�[V<���*zd����X�+���-
XJW��R��j�u��3m_��G��iLfT_*JB��l#�x�ґi��0�)�+�Ϣ��o򕘟~���J�����q����,�z�<�-��k���=���.�*�\-�>�_)�@�CS�v˟X���	���ڽ9���Y�9&��n�>��O�g_yۤ�>�Gd��V5�N�ܵ�	34p�z,�&���6�5����Sü�I�сR�iա���"��k���HVH�<р��( 9�1qlY���C$_݅c�\��/m��f�F��+l'� �Px|ϼ$����j\c!*h��l��)0����Ni�L��Ts*�$�J�G2 xwVƒ���a��L���Iyʲ%�����j�4>M̸%M�Źs�ƹA�y�)���M��6�t(tv���P��>3�<��!F�^'7�<�f���Ñ]ʬ�+���+�˯��n��/]ڥī  ��G�9��#�_�m~�l����1�	���m�1<�F��FJ��'c��w;}D��:V����f����!���)k~��˂�P��(贈��VB��P�Z.Q��.����.�J�՟I�N�_��e�X�@40֫�DS���Rͷ�	�y��N�1ܒoc��`Ν����x�e@U�u;��s ��Z-��:�k�����&e\Vja1�}��Vu�H�E=$�az�Ԫ�;���~���3!�n�S��1��Х5rA��˝���Ʒw~7b$&a	�J~=�V4c)��j�=�-��,������|4��Yϗ�DympK��dr	!tW�t
�v�i}F�]ewD$�.�F�A���l�S�(���6E����\����uNƞ��j� Kx�|�����5�b4i����l_��6�t"��6�
���r�]e��͝r��0��ҎcI��B6�E��%�-�6�O+�]ȐJ7��S��U��c����FY��PT[�ʵ6�c�Y�q��s�O�\�u}2O׸"��=/6v�m���uD��s{*ʍlA��2��3�u��ny��C[>/���P�{�a�I3Q����|M3��f��J,WR]d�i�$"��&6�'e�w�C=��èo���3TG��=�̀���­��jy��wͳ�hd��{3"%zZBݎP?�ڂ�k�f��vdU�B����,�;������H�Pʭn	���㹋x���'y!m{��(��\y�����J�I��07u��^�F��<wD7�a�1S�C5z<i�I/���!׷,)K��٤TH��f���d\��7�?N������xAu�t���km��=R���C���
7�6c��u�;��d��!�'5�3�.EE�3��d�������^��X��f��*,_���0a��T&�^M��7�
��u�"L�{no#F��y��=Ė]ч���g޾]]w�ƒ}�)��$z���7OڃF�� {?�zъ�\c=��-�cQ��}x��R�0+����Mpe��´"kcX���U�{tSr��|��S��®�۶V��.u��s�DGYXɣ?��V�w@|���~���� �jo��=�n��I�w����J�<)�x\��k�',ku�0�T��x�o�	@V	����`XW�>�Q���]�R�
-#vXmz�VH���(T/e������yh�=�o�� }8|������)~����|>� ٝO�2?�����s��^t4^�q���M�̝8��yca�]�ϝJ,���g�C9�M�,f�͸�؏�Y2Ӛy�ʡ����[���9� �O�����5x����+�@�-}J�¨�ǂ�'t3�Dn��1��!�Do$N���1Nj�60��jc�r�`Y�[�}A��� �������n{�Tt˓50r�U2wr��뀲Bm����#����!HJ�wC<K�B�1���M�H���R���vjX�a��*(���6US��2����|�fuGI6:Y��a�=��/���Pc��Ɂ����Dd�������K���1�g���&u�!Dq����e*�f$Թ���LE*�^�3�97�&7�[������D� ��O3��N�;H��P,���/�N�KuaS��!Z�����N�~Y�02=�v��دc�%��um�I��n����(O�0tA�@9��R���:�H�e����TfN���ȍo_����s��ۗ�b�e�;eKlIp�L����'�	0�B�s�WFw����oh��)M�����~��pNT�;M�"!����^�w5��G�1�J��y���HO�P��߿��{��H����)�0q?Z7-w���*���W��/�9���C���6�'uJ+��ߊ�5�%[����O�,6�lh��շ�Us�m���H�c¼����tJ.��,8��i������哞�ڣg���P
��������>�<؏;�=IM�ѩM GT̹��	��-�y���lì'����.��9�&>L*�X�%A�ȁ[nFS��W9��ߓ�a�0���1��ؽ���� ��E��P����i���]���6�)��B;�=-aRqf�"�L�MOw�'�;�T���m<��xB\��J�M�ZW�K��\.G�m����s���k��=�T���r����H'�0)Q���f L�1����'_�+6��j?m�Sm������{�w�8�Q^s`.2|6�q�p�lH$�,҅����]�fCi�]����[b��[��'�04�Q����o#������曽�4IqeXpYb��$t��BO�=�����T����Նyl�X ���x��J-/��ΑKجc��g�@�6��mvs�/�@�n�~�o�^����+77�Q<���_QJ��tx�-DzV ��L��dגi�)H=�rB����ݔ��Qӌ������>�?���)}�2'UW��X��� �@7� YǺ~H݆Y��ϋC)�,L�cu����â�� ��f�`,;�ynӨ$o�;c�X��΍G���F����P'�����t�9�c�a@Wy�SǍ�����-���I�ߣ��@�.�8���_�Q�>��H���w螙�\gUj�p��O��W�)Z���y �ڢ�������}��q/S����Z��\� �ȕZu�"u�+�Ir��=e5����h����J�{�9��n��`I{7����n+�Y[�oq)��|?�֌�QWA�����T���p/�� 
*)Z8�*���|��!"Ip�)�wr"�k�d�r��q��ϗT%��?k�ː*I��O���%���>'�q��x���s?m�ηnǣ���D�y�~iC�n�@b���'D*���
|S��ӊ,�m�^i�N�O"�~���S�Zտ�b;5��U��
�a�uE�(<���7�,D# 0��rKrfNv,��6�UVD�}���D�G�nCe7�o��
���Dί�`
�#�l��z7FhUs̛�{��!۶�p�˰L��3A->fQ/���Wxͥ��k�kXC��if�k/b< ���ūG���c.�.�X^3K��1�I9T	��&�}��;U�pH(ʻV7��(��;%H�P ���\ۓ멇J�$i��M�vV���^���@7H��/��uͳJ�� o}50�9�^-(x@�T��	cl!,ȎO.�2?�/*�	��� �3�2�渙��ole����(6��|]�Ł�G��!**��� ��9coR�$# ^Pj@I��@�{��@lDՒw�.F܋�~B|��k���ج��b[+�%.E�B^�@Kʼ'`zI��4'5ڏ�K��;����
%�9W�'KFޅ�@D�q~�a��K�un9�K*\�N��N6| l��In���a��JIH׃�[��r���%�M ��F���
U �76�&rV��[�toa�_���|��B�F>�����^E(�Je�$��,�$�Sv�1J�b֗١��.�\;}`�`|>�1����Sc`�_2�	�e.���g�Bȗ)Fw��y4'�N+�D΍��v��C��ed}=��lU:�b��	>����l���ā�e�y<���6�c�g��#簷�dDC���ϊc/Cs��Ëխq�������Ar�}rz�N6X��zj1�Vص�*՗N=�{#��`UɍǶA�<QH+͛�� �M�	�}��W[u��N.�jE������ҳ|�Q��n�z��Tg��|�t�K�JҚg{��=lJ��I�Y�Ԟ	����3#j��`�~	��k�]�W7��ڔ}(:)q�'M����T�U�m���!���[�0�e�� A$�AB�fC��|�v�į���+R~��L�y���/?X�BE�+�G��5/q�`S��]�9�Yؔf~���P�al�a��2%f ����@>���	m}�kSxCO�e���%�<�����T�?�a"q+���e��48�>A�@�J�1��*�:Aa��ic�Dˍ��q�FQy����l�)%4�J<���Qc&<��9���6�$�a��g�#4]����OBF��aW���NK���q���Pް�S�w���M9"iL9���PK<�/���m�����d�H|{�I��}�8��W���?���D�b�����$%?FK�Ӟ3%��v���ʺ������2ZM���!¸�G�`�ּ������>8�LV��[�C�,\�Jq�?Cd}C�-�q �|b#�"^.L�=)����;G�צ�B��ײE� ��z�b@IO�����`O�:��]�����)�'>�^�e�L��h��ʕ�|�OT(\8��Pr՟��jX��Ij=SƯ?]���C�|��6X�V�n	t��� ���4�B窝*G��N���H�L���1�v 9̻[ܑ[�\3���9�"N���#o�i��
���Ʌ���
�7!:�E/V���c���r�?������ Ķ�1�`=ّ-L�9=rVN������j�!�A6k�!�aR��Cܣ3ϋF�XX	��4��B���z!*}���<>Yr��E��K��6�u�,����@�]l�{9GK�Y���F����;CR��~�C�F��Pnf��4�Ҫ3��?���o���(a�ҍ�X����I����v4�T��`\�V�Н�u��P�1h��l#��m�����(?�s�W�W��D��`����(=����(Z��!�&ׅTy�[4Xi�����H���AY�6����;�6�s��t�����i��p�TGߺ�����Ȇ�ޤ���(���������W���l$�lxX��-���ÀJ���~���p(p篈�U��ɩ��@oa4[޿�EǞL���LY�r$7qZ�`���Q��s��l���s!��)��,��8`UD*�}i)�<���i6�JK���`��Q$�Ն�b�OeG6��y��F�7}!��.�;�	�$��	�qJO��O��_�<��43=@窌��$�s/�0��s2������BZ2���V����v���Ij�.:2��sj�ץ���@��a��2�Y���Jo�0���Nn��c��>���s��:�@��EL�1�n�!B��sd��k(
����B� ��:,͏�)��W�-sse�^��v.V���C*�ՒX5��|gzSE�:2Z�v��y���bO�k�����Ā'N��f,�	�	d֎_\C��o����2���"��t0d���|ؔ=�����jC�e�J�Q�2l�]m�.?�~Q�z~RSWWˉ��D��C���n�n�����\�}2�<jl��EY%?�M5�'��V�˕ka緤��?`�w k;$�y��V`N]�Ž��<mn��X�5��#�!(��X5��I����ىQ����Q� �-������I��Xn�8�Xթ������|%������qt��m�$T��M��H��;���D�h%,UۆB,�u54f_�H~�x�S��yZ����(���dux2���JvV,�%�W
������ j���
c2����@�w��zl�iw3�p�-B��c��-�	i9hn�1J_QY?�����U={5���]}#��{W!������8S���R�Yɒ��癋����U���em�����R��Z_�Q��$e����rt 򃬠	��D~g�N> �J�����'OsΔ�eʑ��Aҵ<�l�����J,6��9Ռa���m���G��R�=��_p�5Ӑ'�`-�ȡ/S�5�:��>d�푇�O�1MɚS9A.FH���%�����)\�j	 1�:a�70!�rT{�
 Pfxu��DD�
�	�>���	�^�zZ�;M�24O"
ź(u)Q��f{k���yBv%��ƍ�n)Y�B܌\��y��4y��B�~�1�����r����ϭ�zƅ���cX��s�ezOo���c� ���)�|�H�2!m���z��}S�?�@�hk�'S�m�v{�ۄ�G�%|��ee�U_�wE�Gn�/��-�@�~���M���D2����2Ey����s3?�H�!]A.S�xc�z� .�'N�8�Ά;N�����v��Vm��T#f-��-�0�_��y�/+N���oÅ��w��kbL˥;o�ߌ��$6ߕ���?��RD����j������Ҡ�&���t<�ue�]]D��m�\-ÿ���|E�P�rAloP��cR�Ͱ/"
#'}�)��<�u��&��
���ܭ����*�U�hʨ�1U����)��K_F(�������S��ܟF|��!S%��@yG����j�����L�l�}{gI��.�i%G*����^�r�0}��k�؜�$��5�YMLD@����Q>KZ���0���ƿO�>���M*���^�����]�.�u��r�<�ǲV���	�'h񸖨j"\���������/�����O��K�g.�4� ����\�b� �e�6ҵ�v۱�V�wj<���u������Ö;$N󹅋��N�N��߾#�{�TK����mRT4Kq]o�Ư��`���]�B���M� 
�&z�����C8!�e����+�B�1MH��	��n0��ZZ �I�А��g��6�>k��C�L�t�?ą��w��Z͋jA%���i����:9T����ۂ׀t#����5���U<Y'3-y�덤�P���R�|��<l���mi���BTeg��v�L��;��sU�0��E�*�he^�<kEg�"�f�+�Is3U���ܷ{�ꕄs|E*�f"�?���{��?r�p�
j��rl�b\ﶽ�S�͒�z~��m�9K�:��2�}���r'x���e�c�����X��{z�eï�a�Jz']l�6L���y�d�sh�7J���G��诗p�~*�����g����y��q���!�D�c���,f���=_�΃�݂!�Y`о��b��� �lD��������(�a7��a~G�f�P�F����J�����ׇ� ��K�^�@׌B��~eR���� ' �
��#캯��.���\�G��WE���`e��i�boaN����G
�{�����zZHI�����kv��u��8�l�Ξ�C;?�i�:�E>
��b�8�G�rX��ڳtL-�tm���w>̴̷u����1�o�`=;��ɾP�
]�;J�����<$��s��H^F�\Z���dpA\ �Y]��M����^��;GP3�	�����z�MGsP􆿠�����@?/��1��rM��i�u�״P���k� �M>_�e�Va� ��� 6���m�K��6��Z:����}~���R�B��<I|7��G�=���o]ڒ���yϊ)+�O��:lƛ�[���Ɋn2�9�<��I��\�A4�M\�X���[ pT�N_u��K���.�7��HP�R����X����{b�gow҄� [{�$&���*�U�5)��&���+G�޵��D=����Xny��y)ԄX�ݞC�Ym�5��]��s��4P`���]�a�jaerǦn��0��!�������d��4� R� +\y#;+��ٴ�p`�_�нs�O��Ч�J�8��Ҟ� ���&
��Ӆe2SZ��M�yN����V��� ��[;���Ek�/��~�b"}�Lۡ5s���_=Sl��jg������\-���Z�)��ݳ��k�8�x�E�� }����90������f�דz��M��3w��Ω}i�fj�1A6�5g��V2}j����3�F�PCٽ�^�,'�0�XU,�~/X�2��]p�����-��/*2f�vD���	�r����W�a��OX��Ӱ���\��V��g�bD��+�L֙v;��$�.)y#�n`l�����9�eB���5�4�5j��خ-P�]��p�
7|�����f��3�ِ=B�C��e�<�Y���_�k�7��e�޽�
����l`P=!wd�J�ǋ�֩�_T'/�(6Y�7����g����5��n����usڽ�1�ZV�z#]�NZ��D.I��Jg��e�9\���[�a�)b'��������o'�K��̈�a{��i���M(g��E��V:�u�4�"�|��\�[`�6v|�Q�*TjZS�XJϷW {� *���"D�(�l�qyP���5Է?l�!
��5&�U���E�-�`B.��m���1n�^%�<���2R%��P����j9��F)��3>���W/Z[4)t4����c�q ���w�oL�P�p���?�s�y��.45҆$�!9\����M�[�^��R�NG���hڅ;�We�!M��osR{`�j֬FA���R�^�0���A��yE�G������}W�/�j6�p��Xc������r7%2���C�{��<�������o�Q��V��zđ��ꑟ�&6K�F<��[y�|҈ �+��q��tz�[-r5.�n3�?��A���s�}tfQ�ɏ�k�� ��$. e�Q��f�^����%m��8u3��l[7Zө>�&�y.>��n�X�!fEs���ā�/��6��ܞ��`�Se���Jc
Uv50��j-��?g��p�gcW�O�_�hŸ�8)S�`��m��
�#:?W�0��u6)*��`��â��M#0��z[4)w&�~�L�|$��B�x��I�CS&��e@g-n\�r����fxL��lK�Ëp��"�Z3I�zm��O�?���8��Y��IW�1Un�{؍�JS����س�>�V9�$Cg�xlwK.xL+K�	w�G��Ng��V�y������n��Q1+�ӂ�g�Z\4����Qhu��[v����1q��D�2�*�� 
���;��^�s�/�j��F�����1���ʸm��M�RR	��S�ݿ�6tԬ���P"�c��B�ڔ�j%���7#>J�%�XRH���z�n���,���2���/x�׎O����e���:N+�CF�''�;|@��Q��@I���K���/�y?�+�-L �-$ud��v�횮~�AeZO}vlW�{��6+.�fUi��G64��Ĉ��<u�E����p����'�l�,Χ�j�_rKiټ�"6~b�qf~�(��q�²u_��R( ���ިT�-�	�[��!� �34�#HL�v�t.��%b��b�25zt�V�x�ާ@ m�\��>O{iH���$�ph�ķ�m�T��q�6�d.	�-�6*��~�j[��L�&ʔ�(��^K�wM�Á��o�F��ն(a�Gd_B�9�ŗ�u3�#���r�t|a1���~��m?׍q������?!���3�=C
P����Q�Δ��HeR�Lj�	'`Ɍe|�XP����;��ǀ^�YxB��+W��:[��U8�{���~��qG.;�h�O&O��ͅ�^���G������j��5�Aр7?�5\��Vz�.�+��B"a��;q����B��*�݊ʈ�e�1���7��j��N��7�;�'*��Y]>lUXX���r�b4 >��dQCOc�;���R�`Xl` 6'�R�R������,`�J��"��:0��S��'='bzڔ:��.J)��N�]9�<����~�YD�%𻃹B�3,b��؅����t�����8��'�9����`(�`�\> �@��э'�Kih�CD�lXJ��67�?�T��p���a�ټ(�@�~�,�
<m��ӘM�x&>6�2Z�h��xA�I;����f-x���ޗ�V��-��6m�"�M��̩o(wB7#J��T)㎪�q�(�Սgm�w�W��dR�\����g?VM&/�l�4���t���h�M�H}�٧�w���`�))��Y7�ɂ��L��f��|���ב�=
�TG�MA'9t��VLGGoŚ�E j�@�l+a���5����t�H���A���]Ҷ��Ԇ�! Z�E+�,F�!�V����VV�U�3ؘ��CU���EYTj�,%��8�d����sIz��^T�����L�s"�wNr�V	���M{έ��_�Ӛ� ڷU��^z���k���1�xh%��)n*���Ȭ����R~�۴�X��z�ܼ��k�r?W��Ik
j%_�;��	0Rp�ѭ`B	]�2�G��	I>���{���}+�Ԩ�`� �-p�a�x���ؘ	<<��.A�����X[��a�Z,^	ϋ%"B�e���h�L�����v�@�dS���0ǲ�g�8��&�)4������:��v�,[4J��w���dx�M��ypŨ@��<Lg�=Eh�7��R�b��KD�r+�͌(H޴�wa��3X��$J�k�����-���!�y�����ܿ �J����l�j��b��9������H�T�H�f{M2�;.�l��H���rB9٬"��J�6Ŀ9��3�X�w��+�Sj��l_����w�d��/���b���O�$�g+u�ɼ<�0�Jp�U��uX�q���׷8n�kR��?���Sv��{��Îc{8v'�}Q��1��>̲� �崝ht㹧ݯ�t�tlvN�g��_{�@�(�h��8���h��O��E��m�W���A��2�UQ�>M.Tx�&f��P�� ��	��:w<����-���,N/L�l�L���!��������q:b%� Ȃ�K�"`��Rc�z�.�~V)�r�k�Gx�B������\q>�(�f�����3&e�~��=+��F9`� ��
����m��#r�{8�U8q\�TK�� q���n��̛8h�o�
J�`���/?�(Sl��n�vq�P��r8���6�.�_��n0���@r�̎�� ���c9��6���qķ��[�7ѥI�M���`�ڵ��1�uo�w�'�մ�A��o�'�(��+$p�:J%��U5����p@���~	�F��S���\	��߄L�ed����r��7@ߨZ�6��Aľ�R*A��q�&�}�����q��V�z����+�_/l�aJ�ƻ47/�,�ѓk���dr`!�Nq���֏s�,%���`|ԇ��?L�Is�Y�ز���!s�b��re���X���f���E�a���t3�HKҠ�a�k�
��L�;�_f�)G�S-�c(�$�&"5��Z������S �$�G����m�׾��d�t5���ZW0u,��ˑ�:�Qfo��������E�?�Q�/T-:WhI~�fDN���6���e���$��D�B-��@�=k�Y�l/U��J|R�V ��/8']@b��U'���NI�u����*�AH���LBQvm��A�^�q'Wx�qvq	�h��;sJ�Dl��!͎ 	_���X�#��>�7��v��1+c|��[�p��k���b�+y^f���ݔF�fi�YC�������
�R����E{�~�p��)�
��_�����6#�oW[ ���0���W�������2�#�;ˤS�|��sI�"�/�ũ*�������ŋ�j���� ���b�tv��v�[mʃ�=0�����,6鿝9F�LϐZ�	C�M�?ݐ�g�[f��~����_Fp�қ�;x
��s,�ȵ(���}�=Le�Є���kR��l��=�;��$�U�u`F4&p�ev�<MV3����ג���7��K,������q��O�p�5�QY^,;Sq��{�54��{H��e�TBR���E+XsZঀ<�Tۛ��"N���5,�����M�^�F�n&�-���0&�c�J.o��@p��m�3v��Be��E���N-�X�P�7���r�<d�5DJg4x,u>B�(_$��=�ҡ�T̋��4�ɏܶ-���܇_AD�
\��b�˚�յƍ?�|-��2�����͙7���t[p�Ps.�Yw��>Ƿ�2��.��t-w���/������=��C��֢�8f���k/��?;˼�r�D�:�~��N�)�ޕ=%M�T���������Mo�l�kIt#@��)P�e_3�)P�F�<U�X�����΂���it��^7X�9��݈䒔���s*�=Y�C�vOc�1�m��U��m�m�T�!�^T|6��߉���2��(���>�WCg�:v�#M������m;��%E�&�0���;�����$e�#�{�i̡GF0?������X?�ɳ�}�[���#�k|G����\{_���>�;2e�;����};�ʟv�A�+iL�B3�j���F-��̫���a�Y@��K�:}�wa�{��������M�]�`�t-�~�Κ�k�[�G�9`�xp��*��� 7VGeq��H+0�2o�Ig����qa>��R��Z��IצM5������e��M��O�� [�w��{�ͺ�)���
LD4�)����73h;8'+�!F�'��ε��ӟq̿iG���tZc���^��`]N��"a8���f�`�uݿQPL	�bQ@
@f\>�o!��@���l�C���K��ȘS=nq���� ^(���8If5;��Q�����[y,�B ܎֎�Zz�/k�߃[����޸� *J�C��h���EJ,�������NKVGR>��Q����eO�"_�}�����"�t�:���2k�ݢ.��0"�;��ު�Oz��(:<_��Jn� �W"�~��b��y�܇+��Qf���	p�Qh�Á�w���f=gTm8��> �v^��
ߑ�-�����/Z�>�hd>b��y�B�4��!��D�[wU�F�j�|Zˏe,~w�I�*-i�9+�u����c7@��ulrP濗�&��N0�j�DĐ팈�q�3���^)F��h�Q>?�d���p��H���`�I���S����&c:����j���K�s���
;I$�,��[�"o.fw̬��>뤇����\@��&#��9ӫ]�K����(~̃�vށ~�k�CëӋ��$�.xp��~.5d��(��I���?{�)0�~�م���r9sE���S�[2�䌥m潀I��~�S���Ǉ�zs>�|�ϧ��i�sU�U�hZ�ɷ?j�a��|lxa���v��^/�4Oc�7��+D��z��VB�<�������|�/��s��f������$!���JT�U(F�\�c��'z�^aE>�dG�W<�e�L1VיE�[��pTb��VG�p��M.:s<�nM e���[E�U�㾾�?�9tL'G�8�i_�Ϭϫ�S+ʴs)a���;gL��f�`̭>+^dE���	7�t=��j9�!QO�$��Rm��&N���E_���������0C��d��;��9��>h�����,]+Z|E�Q)��Es��α@-�a���a�y��������iZ�X�n�cn��C����U���`!>(�ȡ���W�(�ТVn�v�/h69s�@Q��̀�C�F3���\���ݱ��K%�]�yz2y;�!�V�F;��)�GmW����z>�#�Y
��yp�C� �����+7o֟>���@��L'+�5�qB�A8��o��CX��Y0[�˨� �y���4���
���:���Gsh1�د����6.���?� 4��� &ßH��M�� �6ݨ#�Il4��w.����+�{w��޵�Xx	g����Ϩ�����I����.��-ꑵ渊��Q5Ŀ����̊Z�sa�r�kk� )�Vb�� ��?�dT�nj~s�e�3��u3 ���@��X�J�}�����{x�W;�s�R�X-..9�q��9E!֫4�U�������pH���s�v��Qψ��"�u2{�Jr���*t`X��;�m��ÜNy���Lo��׎�/��-͗�%/��w�)���H(��R��J�+�]�g���O�j��@q%���'��!��6�����oI�[�s#��"�?�t�����Ų�U�Y��) ���+ǊiÓ�<謘85v�3��'0�������-ו�E���1c<�(��Kxp�@6��۟�w���)�+�]����PR��栱[��T �%�ӎ��G�f�ݥ��B{X����HGn�\�W�RX�y��O�̥vI�؍D�~=~0jH/ׅW�+����w�O?��"dV�i�]dV�N�?�1=���k]�HA�/�8mM�3������t��D�Җ��A�Y�4�����q�ʩv95��}��*��e��Z�0����=�"�'�Zp�k]Ѥq���G��9�2�P��Qå��uE���ͯ���7��w�y����.���z�� ��ؒ��P����ժ"��Je�][>���G�L���L�W��*�)kI�4��G}�a���/�E�2�����|�4��F�Jh���fZ2I�릺��R)UtI���ĵ{���Vg�r����BoF�}�u��eREB�9�G�o�5R��:-@��]����d��zV��8��1��/ljn�,�Œ����>�\B�eH�/f�\!�~ss��:e��ȵ�q�k&�F3*���Ö��n{�[�����\�7��M�^�ƳF�+ �ci��[*L�Ԅ�u�Ѣm�	�NM��k�5����
���jɔz�ŏ(|��其Y�3B�����X�9 �R�:Uq�2�Y�i�z�[ج�{�:&�&i](? :��
�nO(�
��f������	��s�Ҷ7��^�čx��@I��]�����"�KSh��k<R��;�CUާ(u�q!��(7�;S�l�J�_ �ҹ��k��S]��]E\wklf�V5�M�7ۺ/���A�O;�j�����Mn��F�&pG��S�ݴ��������l�N'�!�~�$"����DV%_o�
"A	�Kjf,���`R� �*���b���ⴅጯ�lN�������� �إ�%mrN��ڧ<�["��� �"�^��1�\���H� ���XQ��ēv�y����(:9G.�]�J�n���`���掑'b�"괻vM/��'���h��'�-��� �4�l�{9{^Ɯrɬ-��r�n�����7_[2ZKK�4_�K��9��6��ymq�n*�k:2���Hh�f��� T�=�C<�����,N3�ق[�g���kC��ge[���6K��ХT����a������o�|���/Gj�л��g�{�<N>_I(���t0��Sj*�;X)�ǩ��hP5�uJs��+���ĩ��1�`C�~u�T�C5�~������&Jv���9����
�0ìH�筀>f��)oT���x��������*�d6�WQf��Ƅ|�;+�	-�����uj�LP���UEui���oн%��\��u��#���U�y$ƪlo��İ��G�}�R0x(�(��x�4L+����cp}�!���������D�����U��/~�>���C����n���h���DJ*��E#�#4��C�x}�3�L�X�"�@)�'GU�?���ꤓS&��YD-�?�u+�Os}r�������ʏ1�Cqk�]vcX{P�D�n�1d�y>��?��:JžEb�N7�ߡq/b4�2�����D���g��ڝ2�1��0ne�"���&��FW�3�|��Ծ��j*0A(���p%=�y���=�C��@X�9:k>)I��?�U�'��>�K�N�� �GK�"'����w����D'��<����m���Pܿ�'ȼ��W�'���֦Jr��8��3s�*��Q����:�f�Y�<��ζ1�x]��Y>�-2�(`�hR�e�Z3�TR�KR^��Ah$� o:��:��?vs���y�Z��2v�, ����"��Ω.J����e�h��c�xvn4'����+�� 1����q�]3$ڕZ\_�J~	a���~ZǮ'�R�V��̧�N�ő�,�8 �Y�%�f����rH#�};������n�1��o͐�=R�B���W�X�h6$���^�����[�#�
\�R��
xi%���b���%,[�U9gO�ݵW
�ػgN���s��]
�wL�c1x��Ȏ�u�0���U��;>�@!�'2j	K	�P��