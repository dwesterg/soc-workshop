��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� p�X��Y��!�����j�V^�ʳ��*
�,���I�)/��� �����{�4ePs�Ҋu�b'��j����Bw�>Uug��q39�NPU���>��Q�~�pC���ڪ�- vӏΛ�9ȁ��﨧;�2p�kq̭��cɇW �??J���=�#~�$��"k��,�Zz���h�;��89q̮�b�d*6�5����Rd���S펎�d8���)�p�qfƻ5��Nj{c�I�����eTo�5��XIID����u�<	�1 ��!g�nD�%A��
Z-Cej`�d�.��oN]&s�����d���?�L鐩��ԟA^Q�vn[T�����w���sN%�H���7Z��pz#�t4��0w߫�S�'�]KJ���
���>��u�����u��h"s[:	�G��m�k�w,����1D��i�r�b��zꃯ�, viW����]��ɢN�S��z���E��aTO���5�NZ#�2I�s�J��s(P�7w��lRy'�<�?ӵ.r�ĺ�5180�`�"`=�h�ې3�n�˶O��F'�8H�I�)��]a59��wiﾗ�F�1�ZE�c ��ӑ�ǉ?�Ҹ�3F{�M���A0���_B\jB�Ӆk�gm�?s�k�p�μ[��i�����H�M����ZH׮M�՝\gU����u9�,����q���L�Z�����;�G?",	�:��mSo~�"�<H����7�<�\��v�\�o�@�a�c��ݷ.��])�VO���\���6\�G�P�w��'�Fr��� /U��^��҃�ZP_�[)l[X3����\�+hd��N�L�C&�~�]i��(&� .$�"6ku6�`�#�ec0O�<���F�S�!L�\)S�X�V�L������zr�����7uo�Ǩ�(k�K#3�~�ȹ���*��������;�8� ��ሠ�=w�i7؉�k®��4=����6 �d�x��䃏�G;���5�#{�|�o����� ��_x�����/nU�jM*��д��}5$x���f�#�%&i��;}�"�G4sc��w��.͹#AO"��J4/���֗A�d?4ϖk�i����uC�l��l�����I𝂱l��J�v���a���c-�O^J�ɧ�}/O*������������Ҩ ��s�8S��E$q}-�(�q}��ћ0��X��z�>�X�3�r��9k'���&�%-lY��:zt�LeͶ��Ԡ_{��WˎU*�&�o�H���~�1�Ν�!�kr�	���f�U��:�e]�i@@�O7f@���v\������%Fa�ꂡ뮁08T��)�@��g���sT�l�>	>F��}A�HX�1��t
U��[:/�H�i�<�-Nz+8J�p����2.)0.��M�]��3}�ã��+r��WP!����0#���ؗ�(�5�9DU~��"�JE�� �����9ߪ�,��z{w%
.�'�:��
-�����Q��܈�ۂ;xf��}[�������D̜`@����q�D����lW�@�1<�7n�Gƃ�����􊴮o�{K6�|1���" ��b�f�Ǻ�-�{��K]h����ە0H�H�Q:T	#��+~%}��O��T.�E�5Z�(��c��L�����}1��^���k5]�+J�>~�	hٴ��]����")�����vw���X	S�/�f�;({�uz�q���J(m��JU:�g��*rۜU`B}#�$]�ǯh`-V%c��y�Ϝ���8MD���1��ԓР�F���$��U����c*��vg�X �]�9͹!��(j��G�r�|�_eΫy��󞿡{����zfPPHj�C��{$@@U�Y����Sh3_!��H�!Q{X�K���I�N����fpf5�T-9F���Y�l��{?�(��PPfE�@��w՗�6@d�JU(@�8���0U_��[��y�����Cck�ؽZE��(ȥt��ăA��9_�,Æ~i�h�ܒp�H��	I(x$����}�����sX�f��:���`�5�jK�8*ල�?2�@Z�f 	q��څ{t�8�ǆ@U�+>cms1⪠j�>?�>Z�=�DgI�6�j(�˞나�	1݄�S�C�G*S�ӬQ��W|��)˨�Dm����-V���TP=G�o��h�08@0'楝}�so��(�t�l1`6����g���6����m�y��<K��8;Q�����)Y�״<Wi����ޣrSY�������}�f��T��3e G�
�4�r���վ���^Ĳ���y��@~�΅�|� ��Rz ��L�D��������z�n�DgQĬ1\�1f`*���>A%d�`�9s�SPD�\�z�ӣ!D4Y�jБ�fT�҆�|���8c`OL�xڑ��\�%��B|)�|h�{j:�l��
�H���T._�4�Ew	ڿwW���cW1&�:�G����w�t^�����a|�k����&u�r*�:!�.��R>tj(V�΢| v� �5���~��%)m�{7����Q��v͡ݥ��Q?��z�>�A��U�:h��������H�ۆ~�=Bc��V`9D%k0��7ׂ}����6���ƫ������nv�_l�����s�ƍT���O���$���8�a'l�^�y�e/��A�^����e�w&� �^�{k��<����jY_$V[K�5��Z����^!\[!�k��C�e9���`�l����� {��f�������������e�ԟ�٫(Mx�(YƬ���S
���r�j�q?����U1ـ�b�����Jh)j�z��-焜��v��A;�8���?h�Y#�WJ�|����Z�3��$k�, ~��=������(����	�ir�,2k�_�NuJ_3�'͏��7��F��s��جUa�� ܰ�(�'/RשD�k����.S��9&�0s#�X	N5�L�!-`�2�Q]4g�5aR�] ?2��<-]~�z����̙���w,8@a>���b��)ޘM���� c�����%��[�J���wX������{C��/~�qih}t;e3�������Ձ�6�6� �����f`	]��Tn�АA`��~oj#�~&��!X�0��2F��a%XiۘG.+��~5�<ѩ���Xo������~^��j�	�+f��K��b����t�qvAu�N\?P�5�7�\�&�G�����îfx��n$TT!f�z��Z��~�~�N+�@���o}��c��W��?9���W����z]�$q�n¸��>�õ�����+�c�,�U�\���q���`���_���D	[ɖlM=8Gn�Z �c�#'`,�����꺛Pk	�����1���]�^u�K�&?T���x��N4�����v\��%����5��*'͆"_��(���e���NDn��4!\�U���k!��):��f���Kg��AjLN:`>	�m�Ķ�vFw'�h�f4�I=���i�#��iS�}��-Ƀ���Ƌ�q̀�q����K�Kf���ub�NS|�k�~lO �$=��~�v����1JP��q��i\��L>�(��@ b�S�3�Be��l#cu�G�]�d�S����쿕s�H;�W6Ҷ|�[}�=�'���'28FHH�ׅ�D��uA�>G8J�������ûj��.�uR4��T�=$mV����l�E2FM>�����X����I��O�xM��Ԟ���=��$�?�{�vL�P����[�0tO�MlK/q`�������r�aƢ6��<(_r�Uc�31v�s΄��I5�
ʵl{8���m���_#H�ԗ#r>2��o�l>Yv��ńd��n�=��J�*M5�AlR=w����mo͢v�?�����t##=0c��X��k�y�]=co�%���?T�{�H���4K(�%�qVQ�����$��[�#O#��[>^\����l����l��'���]��z�*�8Lj�]>�|@��U���i���+�BߺI�\�l�uu�@X�o�`��� (U�ld����u��iK]M��@W}p;J�Dj�0��US�ܝ��CI��3�wY7W��3��؃�_��Z�[h�������6\�F�8�uo��"9���1�z"2=�;�0��w�C�V��M�l�'Q.Bn��묿@����յ!�D�S!�?�;N��9K���ǅ`i�JI�^%��A�**�F}���N�q��c�U���z*p�� ��+������?5@�o�c��N�Gxf(`b��0���
�cP��$.A�^f�N�>L	����&��PѲ�S��u�P7y-
�c݂Ou�0~ZO>Խ�|5 ]6!�ښ���C�\O�,p�o���K��A��zDQ�bׇT�(�۫�t����!C�YB}Wr3�I���f���t죚�j��4���`߄��bi��+mF�U������Z{W��r13��#S��(n�:|XG�Kr'�L1����hxw��jv��zL�wW���Ƹ}?�8�_��m���:�]�L)�����pdS�5z������nzL��~�U!,*��8�Ɛ�W��t��?�B]�i4l���Y5������RD*���W���	\P6,�[Z�*ԲUT����X���_�8��!£3t�UU}���Z����)�2��<�O@�V��Qr�$��(���~zI?Q�)�H�+a��5�
�?�-������~\�քag�e\{=�F�>�T",ͩ/��!���Œ�r?͌ɔ�}�߄h��|���������b��L/uU>& ���TVb��԰�%آ�����&���y���(���)�k��<�"֨���� �DE�؊*�i$�@1��a��T��#�ϼ61��oV�m�/o�7�D��a�����q ,�pY���f�N���g5�̣�������pJz|hק:�S�S�8���w�$G��L3��G����y��N��Fm��[/����68�f,zs�w�5�ȸ�e��).o�K��|�7�}&8EBۀ�9�$���
���><�Z�
= T��+����1��X�%���Ǫ[V9�䄕@��N�+���J4�I�Q�fB�
{lغ2�٣sCc-�f�~��z^�VҖ���`6��t��5)��@b�t+��L�=���=���lYq�*�l�cJB�pПl��r�� ^R�?��������p?le1�Iz�|贛�g�dkR3��i�+�O�n�e��-%>��wx&����	R�!�M��;k�bM�0S��lt&�~����뾆][��;��{�acrk9����N��cm�|E�J�""��#�����'��̚xv�ݍ���W �����4����.���g:�g5�ԭ�zd`�/pJ��_Ds-��s:99q���(�t~X��gE�f�n��j �H�e���*-���Th�\���&Z�{��K?���;��w
����,:iU5v>�<�6Xm�`��j�}��s��7���_wh.x˄]s�<��k�2%���Ld�Lf�.k�p
� �ik�C�
q��$Z�h�x� d�ɀn�޲I/�{(7�E��i��Z����v�&~WE�c�]/�< 4�7��u�<}��8���ii6�%��5�McZ��q��dV��Һ@�s����q/n��YKxtEla�d���Z���il`��L5-Cq���ҷ�~��ŉ2ƏT���-k޸C�~���B:��B��G�D2N;ϰ5fs�����Z�=E��/��%͑]��F]��7�&�m�ύ��$y$�f�P' �Ps(��3����/[R����"�ru#��<Cvr9_�y�np�Y<���4M������Z"'Jؽor��y$ȭ8��h��9�x�i��,�.�}\�J�C񉾏*9j>�n�r���d�L��>�$��>���0���6�sU�$h3�ß�����a��� 0��AGy�'ks�Ab��R�<��ʼ/�\�%�u �"Q��&.7,|�I2�w�)�v0Kz���3X��.��
�oZ��W���u��֘�7����Cp�t2�����߫͝F�%X�Z��߾���dE���ȡcwY�B����aW�� �Klo��0j�b؉�� 2��˵�"��k�
)�ǰ��_"����~<e��f��[�	b>P�`o��d�2i�j��>G��((&���q5
�X#��󝭏u�i5�O�n�O	���8�i8-r'f�]Q�����*\u9�V9<�L��jմ��I���NL=�j>,Ŀě�}\"v�;,�;xN�x�mL�=tCA>K�"l�v	��4i
�?��6?�0BI�uT #�S�kqU=BH���	B3�l�\���q�Hl]�����"�q���w{[��P|���d2>�:�&a6��ܚnQ��dE�":/�R���;�0��~��Ny�/�w��a�%��")N�4�O��
3��w}o�*�%3V�)����pJa�T��D�9��X�R:>���wR*g~PN�_�2��2׽1�mO�D�{e�D�׬=�35dv� }�	z�Pem�����\.�ck}��'@�0��є��B_��@��6o����	Ǿ>Ͷ@*����2E��paj�VS��EKL\�4z��(��u`jk��)}��>-5ZO���	�g�s����ns'L�����i�ո�x�����X�D3���w�ʻ@q�})m}�d��&A6�DW��w*a�\��j���q�v_=!�m��v1�\(;sڞ����6��?�zP�`#�1����]�Z���Q#�6PX״��Rq�*O�'�D@BW�M����k�H��a)OEb�!yp� �/9����.�k�tϿ�F�^$�H���x��ҶE,c9eáǝSuY�Lj�\��	��:�v���N�����Հ������K*�rB�ǩƿ�{Fo��G�o
��Dfs����&������[_c1�XP��}|�s���Q�
�.S��a���\n�4Fm��]9��VE�bH�����_9�zv�Q�D�́���Q��ZZIC��  ��h��+Đ:�p�_��I�,��
�	Ȗ������V-��8�\�夰�,�m.��u�ku����O.��8�p� @�D���O����U�3B.�/ޑ��?Sl�s,S�X�P�~g��+�*�'/���pW�Yk�/Wn�����@�ɬ��yjߧEk'����R}�΢>�k�\_ګ3���<�Cm��`�a`{��02����u����aYV��C��s�XO�	����t9!6O�_�O����ݵ�T���ȫ;
}{Ο���Iό'�C�Fw���B�bX�ȸ�ZG����fbEk��& �h�v4��2���t1�:�6�=��3��ЮJu�;��np�q�����U����>���"��K�l��R)�/�V�#��)TGh����'��F3ƌ����{���Zׇ��AX�ƫ���hXx��K#4����5�:1�4� >PP�'�_&Ѫ�K��˹ȌDk�����RT�����i�.?���X���䶿���c/�F׸2��G�s�͜�l�����/�q�)T�q��LGI<F�ъD�mrY ^�öδSm~��37���W��]���&7ǎ����؏5���z�����43�IT#w~������:ߥmݠ_�Z��9{w��-�� P�xW�BZpQ���T]�K�=�vٔ����O�q1Kr7��\Υ��A�,����lV�,t_�r!˚p,��͸xy�Q��՚�rm�O�S1Q���;�1Jl�',sO�2��C���_�����\R�D�vl9+XYX8z�3X����NZ�Ѿ/�_(�V\�$���ڦ�چ�v?�4aI�Ϗ���ǫj�����,VzsZ�4������H�'8WVĝ�|
?4��{`�I�*�}ۡ?�'���������*��Y�z|�1�������?w[��fg��s�����k2x��/��z��͛q���+�2���r5���;��R��d�1߄�A��^R��K�g�#ہ����f�f����,�]|���}~ϫ��L�(��x\݃O׬��Mv�˯;�`�X��WyKx�٨֞Z���.k|���4��O.�SO�d�[β��i�N�:S|0�M �O}���ZX^d�#�B��7r�ܢC�Nb�-�Q���A�-��x�s.o�Y��O���v���e�]���,�z��ò۩�Y���q���=~9��*�FC�����AB^\T�/�^FAb��ض����&��x�@s2�1��g��-c9���U�mͷR�e[qn�iB��pJ�^O�%Z����k��+L6�	`���k:��+�2�)�O��i�� ����W�'.�QH�ifͦ)�H�-����͍&]�z�b��"�w�-g*���	��+��4�E�
3U�s�Q��P&g����Q	��0�aPas���cPj1�H�B����P�cX�&��f�j�#!�ɫ(��]� �/��[��J��~uZS�b��{�{Fô����&�A"*5��� ����j�%f!E�'�')������I�5jQp�V�z"��X�N���R �����3�� ��_rm0�	1˧"R�{�ˉ, �nn�ا�;~yI\�h��i��x�% �W^�/�=�a]#����M�K�f|�>g���YK@�� ��u����l��}<Xǫq��$P�w�+�ZY0jA�
�s��!��(����;��e��m�1�Tga�he��\��晟���6& �>�.�M�c�|�DQR0'��u�d� Ξ�!9Tb�����*+H�.���/{�X��f؏����$$*�j7nt���9@�m;�rOn���E^K�Ňg��v-�Հ�@��8�-{��\p�ĔM���1XtW���#���Y'�%yz,�D��v����Ή|y�B�NA�c���X�����	���`Q�gl�<��KG�S5� 	ߖ�%�鐫10��A;�q��Ѵ�JH����/�P��R[�F��8`�������p���`�ŗ�D�aY�$���Y,cp�M�U�k(͘����p2�*��~[��.��Q�o��I��}�:���߽��B�;:(�ݱ��fq
�%V��Ip��n�tp����ZK7�(�G����KAX��!X�b#%/&s�J�Xu"�,�c1�P�1�W�QC~�����dA:+�Z��z9uNZh9S�f�����OfR���ȖEk5���1�ܰ�i?���v쪪����,�}��{�T-]aa�vݠ,�gͥ_4�ʷ)a��<����l�Fdrzd�\��Y�9���֢�[�JqWy�h���gOsu��-��^����-�?ަ1�,���S��b���{��f�H�J�)�#S��9nM>��9[I9IN8�b=���D�m`j�9�`ue��%Z0s�&�D(�g+�f��:�DI\@�
U-�y����R$���]��~�V2'��a��o��ĪnL}���~jC��2�o>7�B�V��z��2���SSx`�l蘻�:��y?�e�9H�+�#�:4_aè5�;M��xЋ�㲲�+��Ҭ����b2�8��j�Y���t������@��5�
�Ka4�����Y}y��|O��ߡ��[�(��	4X۫���u	�X��Զ<�te���~+�5�5k�ydO=m�V5W�!���*��RK�6c�j} �|���þ��,���f��X����l�oky��ř���H\��P S�'!�oI_�6\3���x��
��EyY��P0	 q�d�
<��*��tyD�E0���+���PzYР�i�B0�3^�u���ݛ䞪�"�|b���$�O'B#e�#�,n]����\�)NRil>��d�H���I��p;Mi`4��ւQ3��/�m�ݴ/~�) B���&adIt:Xa?�lkb�5�����J��zw{�m�����h9K5��._���G�m�~>S��/��JԊq	�[��u~�xVZ\?�~1Х��;u-v�x�m�FCU=kt��f�9��7\wͯA 8'y*YSM��J~/�=������,u��*NC��Q����2��l�P�(��P�+PI*�3���_V'
�>8�䈐�,�W1��7uLJÝ^5(�F�xV*Ս��Q0��<���xoeX`~7������S�8�!ڳ��_�]�E�,��X���J�$퓸�_a�h�l_�R���._���1�#P��vu� ]8sS��Yi�J9��4�}UB`#YG�Y��0K�C�m�x9��ρќ��w!oZz�`g%��Qt���D�[�	!@�=-�	>@m�t���2�`��j��M^/���$��7C�	p��3��	g��(�]3�K��ٖ��ѷ|����M;? �'�60�;��4&�K��7�R8m�X�r���i{3#cSr����L#7�5!&-WVE���$&{9H�٪#�}/C?�
�ՙ^�R���Xv(�^������u���0�){#���.��>3K�b�M����o@�xu��s��D���/���>� ����Ƞl���gM.�s>#!��;��~��H���ZX��Z��Y�H�����([��#�\�� �o�=:�O�Q��Lqؾ]H�{̞t�-�[J�Nfe�"�7o �n��@�6gT�1�!/��9W��t��:q{�@r ,,�ew/L��aJA���~C��@��-v":*�=;�z�� ��K��Ł�C=$�����4���0��a�}"�y���U�K�ɣ�#Ѫ��s"^r�Cʬz�Q�B�� 3��U�w�HqnjW3 ��g5���%#��3����z]�}Z�b! L��/JVӌ�&����~lfMt�r��А@��~m����	Q��1=m ���얺�{ R�k�V������*v5V�&�n�ˢ��@j��-]�����3��v�Q��s��Y�Vdg�˄��fW�DR�}����iڴ�4;qYPeVR�A:���9:�_�ZOS�%-�<��*6������<��"`�x����2g�#( Vv��J��`(�BN
�S�D���i}��Rz]�1Ʋ�ft�5��TKrx��j�Lca��=v�����5g��Y|K��Ql%U�H"̫�3��jA����v<�K��Nd�L>���%�D�D^~� ��s���Z����ހ�0ؐS�ŭ�)���0/�ܳk��@d~�4S<G�~W�0��A��";�kɾs��(�����1OZ`��~>�ki��H�w��r=��H� � ����oAe�U�TG�'�9�!T� �i�/��ڭ)p)�F�#�4�틙�(�j�-�װc&�L��s�K8��l��Ջ'b�z	WF�#��K�aA�}����� �����/�9�f3p�i�q�iQ*�t�a��>54��I��Y����,�s��:�v+�k4�q�����0�\��z���dz�S`A��}?kϏP���l�ws��;E��� .��:W���v>˃Y��^��W�,��	m������2h�^$��xxjx(�֯=X��NIU�.�Ŷ���Z7�n�����~�t�I��~j�s�+`�4t����ǎ֐��85�#�Gd ��j�]�3rKz`*%Uo˚�"��TPޖ�w׾��
^���N�Ν_5����G ޤ���3�i^<p��fkI]V ޳�RD]��?g���o{����jT�s�<:�Qי��8�2Ue�p���o�E�����Ճ0���~�K��[�=K�<�]�s�[*��DϺU�mg!S�����-���8'�Q�b09қ�q�r�_���$��0A���C�o.���)Ō�J1RM���>��d�6`�*UQ��LGzh������|T8��Izgs:���
��&�-cϙ����&�fE�腨��>޲M�_�.���q��V����rZ5���[�O��Z�ϧG���E#�h�¥��ZV���
������6\YX�?J:yeW���i�<����5�d����i��%�E���gw��tl^:�J��p�#�ˬ]���Sja�Bg��e����C�`i�$�3˅�(�/�6Ξ�]��pd�i���M�KD��͠iS�H�*o9ȱ+�G���.�]@L �f��7T�	Ue����#�����)��E�L�~gS�U^��L�]��1�!F�3��:KE���$%�j/g :������j�R��f����W�
�F�|W�|l��$�g �;�t��~d��֫��p�"\t�3M�;��(���f���9�(�ŦFB�Ǝ��z������ݵ�h�#W`��!7�� R}ϕ�'=�	:ڵ�|�T@oJp���O=m����K�e�r�Q�:&��O�	/i ���8�����?3���V�Q�0
=O�|7Y�`I���w	�OT����yMa]9$X,��� ���g0��������>�Fxu�=�ZF�7��!��ھ�V��/.�c��$��1U�:"�����ӴL}����-�T�l?��Z�'���-nR�v�m�vJ=�*�g-��	�fs�6G�/ �Ď���<�7O�RJ�{=3��Xy���FA�|�����mR����_~j�ٓ� >H�z��'H�?��5T� �eY��M�̃�К�j��k���H��B[tV��$�ƀk������K���׭��b�0�/���~6Vcq��v�57�,1�	�W�в:�kSM4@�A+�4�y:���R\��U;4q����*j�I@j��`vK+t�ӧ��-��̐$�'&�&|��#�%o�;���a�؟"GL�+���\LL�ϐ���m2����?#�5�O�x���ै��Z���*$���`�cj�H]!y����@(��(A��8�3h��:���?אּ���b<ގ&rU@��=x���bS,82�_j�H/�����?## ��V�4�t���ߝ�ӈ^#��ô <9���S\�C?�-Hu��MCv��������Ϧ4���h�}����A� 
�� ���,;OW�z�fZ�Z61�W��A\���j��6�+�E�SBP�T�ڣ�o*KI�n��n�,���qm֗u7�W����)����C����bX;{Ų�n�Q�Bo��  �^!QGv�Wgԭ���h�oƍ/KXU����O�.�B�g�tkc�N,�L����O�jǮR��`�
&�	�w|V��'�����A1��s�����?�O�&'�f�W9f>���7����:����M����V6�2J���ܾY ���7f�T7)׿�-R�Wg�
Cd��r�3�{�Cd�rd>)��t�ͩJ1����<�'[:���7��E��m�B��]�d��z��*Ө��ϗ���-�
�"�o/s������B[�B�`%��)Kt_M�,M>gz7P@��@�di疱��K�Ҫ�Ƒe�F5`ӯn�r�o��̈́lq���`b�0��{��%��שϏ0���Ϋ @zfA@�֦R�"A��U�=��J%;�R�J���O��i�΅U�H�����B���ֲqA��/�@4�?!�V����2c�t�!�3@g�z;2l�Ku�>C*�q�l�=���~��Lw�ʻJ4�yV�h�B�5�e����L������'l��T�Y�'��E���_l���(�q���-��M�<������mT���e��޵�
���6��K��~��݂��쀊��K� �8��#��K�or�O���,�h�0B���+`QB/qhS��M����;�@$;0B��-�̻C�"�Ny(�a��Z�@����{��A�.�����6�9��ؿ5��N~J��T}�k+/( ~�t}= 9�UE�#x�n���f�rtW|C�_��M À^��27���ö�{@`y~��_�r�3.G��Ǣ�dp�z����RY�Ab׳n�ɋ����(A�1�lO�����R#5Nԃ`����}<�\ݘ��6��㑒ه�ʣʤ}ft��H�'俞��nu�/��W�Yt�ƚ�	�V98�j���+_��jv`7`���L1 ���/���6��<��$r� �z���-��P�^�y,�O�x�m&E�,�7������4<�Z��gd��6��T��Ay |@��T�8�+{L�7�����8M��^��x�g�!���G�A�%�v��2��X�f�$p\3E�Ҧ=��qO��Wr�rK|�a&�}�z�7}AN�)X��|�C��3���\\`<��%��J"�m��ccҌ�������)�V\��V|T`��ɂU�0�D�{�Q��v���e����C�u�q�rRY����7Þ?���r!���\��eC���.�D�D���5�;W��]�R���z�	����n��r�NQ1��]�yz"�-c�y�v�[��sB�{�k[G�%�f����{P���F�����dX�F#g�K�OV%ū�f��y 8��J�0��Yn���9�w�����F^4|V�ѓ΄����lv� #��+[H �Z�ެ�[|!O��������80�\a��GT�K�X�ܛ�
���g;2^I����I���+D���oV#G]BՄ0���=$�-�Y):�-����x�9�H���B�8'[��fL��6��7���Ux˙�>�V��0 G�1�d2݉��%���sO���x�~ǌ�1�J�kIk��"�|�KO��ݦf!���5�$q?r���cWk�{�����������J�~��|ݠ����<�h�9�E�j�b}Gb�1F�GcO~��=0�Ԏ	U 6?qh�Rv�3�YA��:Y~3L�e��K���o�S��L�5#��xgO9�p���@�U�vI�6X��ӑ�����u���&�6c����j�D�3��z+�	�j��򨼿t��vxFC�dt*e�UzpL�Ʈ��I�FAY�\��fh
V��߫iA��p�L������H�������}n�a���c��!�E���	Z-���C{���a'8t�!���4���|�@��Y���>�X�r룶�b�	�F�H��2�G�2%<��.]3��:�b(�g ǂ|��O��,�y������.�c	��Y�� ���Y�����gb���T�¥~�ݯjЖ�>�B�ڥ��8��MU�ɱGK�Q�ds���$�H-�&&{������d����2�����
H��_*��.��
D@c������������g4{;���Pby�"�#2Օ>�1���0���$m�[e�~�5�KAOX�}���ɸ���e�d��$���4�2��;H��;&u�V��Ag�I�I�3�����:�X�߱�_��O�H�L����ʁ�W�D��Ò!�{�1�Rh��-�T*��ϗBC�_���`غ�FB�_:}H�@�UM����Yס��@a<6z��;�:�ºv�0?9\��)�����2��^��J̗!�J02yL��]H�_$��ړ��g��!�;<Hn"��\�qs�B����,Ǭ�le��h͟�<S���ɕ�z�f�����Oc2�ՙ|C��-[$�����+�'h	qqrj1P�T��;71(��^^�R�.ftd�
iH �ѹ�3����f��8��j��L�X�^M5�, �apK�g��T�\9}<�I�=[i/�[����v1g*vbn�L� gp� DC%y�s����Z��[��c���N�܏�/�uFtCb�Y�rT�#�)c�}��`�\�;�8�j9�f����Մ�Hd&�3]�#j��a���(cc�����?</��aZ5�� �_<�~]�Bog6Y�=�Mߙ�����4����0�&�����z�|���
�:7�Oa��K5֐�m�*�'i�W��������;�(�Q���D�';�ȍݾ5+�`S]� �EG��� q��a=�
1���=��o*Y�Z�-�{�=�Q���r�	؝�r-	�[މ�嬝�t8j:S�D%��O���L}�U��;���.Ч�OP����,�kѶ�ށ����� ����oـ�\\2���Iެ��/�Q��5�2�p��|