��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(��ἧX��P |�`=g��P��F�qW�4qoG��\�ewQ(^n&��G�u��ة,��(\� 6�S������X�'�i�غ��ƝǞJb05���� E���P7�ii�D���uҢ�P�+м몃u_�o��K�9!r}!�lk�E a^���.iO���f��F�I�����u�%ЛӃ1�=�$���V�n۬M���O��og����1�� �[q�-T%�_m���:���YN����7�d�RxD��|Qnb��P��pV���Z����b�[g<�0As-��=�9��4έ+a�b���N��-����A�:�l*���L�%Q"��qmc�l���&N3A0�ZҚ���}���;[����*}�f�J⁓�"gϤ����K�Ln��"T��ѕ����ߍC+���h����|d���5��Л���^#(p�
��*{k��AssM���$K���+
�H�b��k�>-�<H"���%�#ͬq��mmw�x&��ͧ�k��O�r��FPZ_;�Bl�E]XZq�hb�� ���t���̘���Ɍ@Q�L��]m�L��P1�c�a&��f}"��3HY�!�U�xVގ,��M7L)JqNh_hD">>>��o��cV��!jڈ�6ʜ~��!4�?�0��'a��t�;M�Ĭ&:��#�J~���N�9���:0๮W�����1��K�A��p��~+u,!/|�h��l 0pQ^&(�\QD���Lg%(��o\�Fò�05[Q����	����%�$YeVBՅ�[nYK��g6�����8U�sN|�q��?�w������ �]��iBŰ��^�g�r[BԬW7�㖡�&�S��E��iDE�8>%�[\��aKVg�ᆊ�>\B��{2��L���jQ�.d��<�o��F�dY�T�b�Qx�X�`�.�.��b�3\���±�n�`�׬�04�o�ҷ�p�s2~E��Gq��\S�˽��߰?Z<&J�����;�K���:�sL�!K��-�x�)}���T��J�'w��p<�m�� .��I�{+�I!�Wpʓ�:��2�&T��;��b����~�!uDSg��Ϗߌj�6��Q����_�P��O��j��))�.wgai�6��7g�J�	o١3�7 �ET�� �j7��D�c�O�qvG���z,���,&x�p|��q
l�3�P�pڅwP��l�*������>���)b3A�tJO�h��b0���m�;=��V}�{md��2�iw���q7������Ln�3>�|�n1�)�hM���^�KM�n$qq�宝"A�F�o��6�DJL���l;�f�n�%(k4]P��t�X�z�����3����T�'�E�44�� Fyˑ3YsX�ls���	Ɍ��ES��ǎ�(~l���ؒ!��t�@uD}�����H�k�f'����d��V;3�cr}uEp�s�[���ڊ�/](FK���e��.o�(�$��@˲Hؠu+؛G�0�	��畵�Ի�).B�)(���'�iT��%Ds�-�W��1l��u#��#ٻ��qN�7��'N��l�sȲi��BT�J�u���_I�,�l�@d�xJ�fS�!?i�����h_�����K9�'�ɦU������}K3X��I��6!-�j�����F�D������)�����f�@PrǮ�5���D>Q-c�*B��dЫ8{@�pSI�M�.��ɟ�So�b���P� e����w�Z�N�C^+�8�	�EK&�#����y�kb��<�7�g$�˴���٤�x8&���NjUf���,B-xn�C��A��s��:~������K3�ػ�E�ޟ.�D�&����x�����ʫ!/sa4i,uy�,:���vz-��z��t1�p�88��$���5�_]��>%x y(���͎�.�3Y$�2�JiHWE�� ���3A�A��Mu{����'f���g0Pw�g�l�j�`�d{�|~�!����&�Tv�\͜j)���E�w0uBU�ے�g�DHrb�9߬\�͈E��*'�Y������\�k����� Q��ፎ:�lH��%�]҂lHy�37��=�m�I��~J��=�V�y�	���k�����Y�����c;$�'-�l㮛F"���GF'L@
P1-��RQ��LIsB-�}Ç�w�
04��&[[�4�̵�^H�8TD�����K3�H�p�I*-H���*0�S8=ōA�B����� {W�<J/熐$�����z�H.�>�y~#� 8�[k8M,�9�h�y�\�y�z�RnO�e�X=
�;��-�BM�sv���$�&�riU���kQȜ#DlZ\C1�-س�[��yW�Y�ٸAV�	O)AǍ=�B4����g� ��FVc��/�2�z�(��(�uJ�틔/�L,~��̐�m���S��ދK'��.t-�A���^���KG<��1��Ǒ���П��#ZTT	Sۨ�8����N���l����r���:y��NT��(ee��=čѮ��E�`C��e��'oPobT��K2�^U�_V����2'5�=��4�w���)���kq8��!y[����K�� 2�������\,֤&�B�4�dK��Y�y�X�̒�>@)����-R<Qh�����\�n��n���10q`�%!\'J�����M����A�"�\(٠{����܌�=��:y������!^n�h�uBw͔x����l�I`i/1Y�D,�F�uĶ‒m�f��6�#�������K~6얂��ǟ�u�r	Py!�%�OOФ^k+�@��"�� �lD\�l,9�V����<F���r0����(�a1�o��>���DmYD���1eV����_��>���=f�-ÀNշ(�m�E���~	{��-�l�zd��,|̃Du�������{ە�[!2��޽Cr���惿��&p���q��"Ԓ!4�߾-/|a.�&]�ͽL�$\��rɖps�pY��k�%5_�U����J�cFtw7�X�lo\nZ-g�*~��1�U�4�\��C����9ܢ���x'B���mo��1��cdz���2�BZ���x3mt�ζ��2�5|�S�/S
�$|uU���A0=��'�Qj�
 el�����;�O
v�G��`+��h��DwM����8.�^ҋ`6+���ה�A}�}x�/�L.���\��-�p�(��n�r��gwӊ�h�������e��Z��u�P�g?Ғ��<GO:�V���qL'J�/<v9�f�W 6�yz�*��N��L{�v��M܊�?IAewh�x}ƈ1S����?�o��;�����k�ӛK��Zj�Lt����ΠM��>�~dX���_����!`yo�L�Gq�?���|yj6��EZ�/����('�>chl�9+:�R�[��D��Ĭ����Cö 9|�$F�o�	p>���<�[�DRG� 
��_�����^P|̜��v@�=[�MK�,[ƼM�r5W�%i�_t��5*�Od��.�V·��n���a�m���@����D�����W�	��F�M��C�SviYj��o�w�Q�J!���k�Qn/�����\.��s��Z_�iK��������=��}Q��U�H����G@}$��*��	�=�Z�쬱�w� 
Ū�j�X�e�ԁ��!����s��ȩ��u�ƪ���Rʄ15�E����v]r��%�Z��+�̪�SI]PEhA
���[�/	�I6�P�c�%�$L��� #]�Vw/B�����/o�_�q']���{@�Df�Ø�m�Q� �>��䟉�{��|
-�����sU)ˁ����󙧷�:��coj���x=�_�J���P�|�J��/Z{r��Iw	�;N��� ����3���؁~b�U��S�^�B<�+Z�	[¡��D%�`-���A�U�^�x��)a&_�0�=����%��>��P���c t*7��uxm�>�r��?��G�њ�!���C'���ԅ�3�����ي�^�[��u�ŦeW7Be�;�C��� ��s�����xII���L��J4���7Edh�/f��	kh�L��N|M��6�J�%��ǭ���������8���9�5N�ƕ 7B��ީ-���T]_N���E���ݷ��,��Jo���.�f� ��\�֏A<�8���Q��L���&dD��"�G*�`�bA�7��]�w��s�i�8a�%;U��B��'���b��&'oɑذ�%�����q��&}�_�Pm���= ccM;�R�S�R?9���X����F5�/�X����<VD7���ort��9!j-]P�G8�X�\�<Ͳ\c���Ѽ$��$G�a�iLF�AV�#8k[mW�,>�u��W2N�E��b˷hr�ϐ����1f?8�7Ð7�֭J� a+��(2�;W��&�Dm�'�'f�Z�ӏ��"�&x�� a�k�l���[���ܱV)-3K8�aR��b��T�D�6/�Bz�N5~�j�
�pEٕ���P�V���vŃ��w�r���P�>��0�$��'7yd6���%����Xo�zA,H5 �+"�==ۂ��Ӹf��ճ`)�9�޺	�z0BF�0l�ڊ/9v��
�h����h:���4�瓳T�*U�[E����f0l���/\p6��=(���7�C���������פO$R�͐���k?+X����@Y~mw����:��$.��$��[J�ک�<����JL��oĭ�'�!�0����ƍE��6�xH�(re��6i`-�,t���flӈ>����@0�E���.�p9�\�k�}���+�hޤoV1��u�x��W���q��M�;��{�\��o��
k\49M=+�da(�J60�h����E�y�r���|�Z�~{�ތׯ�u���0w�B�E����8	c�'������^)��L�8Wr���{�D+��'�n42�W�gK��͘�("�'*l&�p�Q]7��_��r6TV>�j�X?
�%�,�� �I�eeQ��Ѹ�p���o�g�o@��7�ʣ���Y*�b��tU��$⢾��3:c�偙���x�u&��Fm���n@+�V��Y||�>�I�E+��/����q(�p݇�FCN.dn�w$�W�Ԝ��R������̆�h�j�c&�R����R�$��a�AQ�jV�r)Č�enw��⧆u�s�F�ۻջ��5��>�<�B��T�����cd��D���˔�m��!y9�`o���H��l%�aʭ��ĠF�j+�A�!+y�yW�Kwf��-5d��3x	?�V0d@固�8���c��u�����Ϻ$H/W�<�(&E6'�A��������,1���u�Kg!��ȷo,n��H���D���@� Ձ���rJ�њ����1 ������[�q=�Ǹ<m��,�v����i<����>>2�b]
̚�[�q���c�D�	��ǋ�+��:���ӕw,����f�_,��B*����Id���-�y����LZϘg �`��ق�(22���v�YZ�rg��y��%�:��f)ݐ�1�sZύ�h2e�<6�Xay{�z8�W�����7��Ha�@�OYC`��i)�p ���T2�<�i���ڧc_s�e�#8�ڲ��N�*���j�H�XX.h�թ��{+��웘B%o���&d�Z�+���y��b��2�H�~ї�<��5�K���w��t}��xڃ7V-�Q���h9� ���$^bݡ�M^=�Ҏ۞ɐ�c�s�o�'���؆k�tѠ	O��b��(9ֱ���C�ui>d`oW�'�Ꞥv=���#ע~�XN�N.8f���d�oBd��Efu*?>�R���0'���\�XJ϶������+d�^n��aP��'<=��z�#m��1��v��oCX2�[�4�Y��SZ�Ƶݡ��i����ua<��T�,����"�l�� �U�B��d�Dt�2DH{AC��
��&�YԲKͽǠ�� D:�\��4[�W�њ�pk!�a�ߏ�Ż�zh0�9KY�\�*c�����cx��i��cUY �4SS�����E�Y�*�I~��y�GT.��R�2`�"��X����'�b�8��5��S��ؠ�C\�/V��+t�m�{�N3=��G�FP���@ʴ��G}�Hw4Ў���
<�Qn82xS�ܹ���� &����3Wξf�<���C�QY���K�;"��ܿkK���>��w퐒6�jV�B�Q;�����J��l�?�۱	�?�F5>&�r.�}dO��/���4%oځq�sZ����js!t�5��[�l�1$��ű!F"⌜V9���|r��ݨ�Mt���&9��8W�����t�Q`��ݐJp��g,�J��OT�e@��m���ձL���a�ӻ�G�P�!7D�x������b�䴢�w�U�WU��?U�e�<�}��{���O�8ӱ|wr��R���QL���e��A�]I1�� s?ԕ�s�7A�*ʥ/����m��w�f#���UOѹ6�W)��YFq�&4!�/^�>�%7�����y7"�x�U�XM~Mo�/b�]���K���7�����Ӵ�j�ٮ���y��|{�
#}���J�ۏ)�a�!�9^t�p���/N�΂,C,��/�l����_fIz)��pQ�:/|j���R6hR��"���R��N?n��<���-��`�He��i�s��ȰG��?��d�_�D��n���z�?�l���-�S�*�Y�Е�^.NB�N����B�<�"ǇPF�ѷsf����Wh#Ckp� ~/{� ��
f+����B��wU�5���!��F�����]�#Eǁ���.�3Й�3��7� ��x�4�x)"�=p�/�C�љ7y]�-�C`ˇjT+��3zٱƑ�����s�d]Y7�k����F~8H0������=�*���y�\$O��b��/�ߪAaJ�Y����c.Hͺ�+E�k����պG�L�.�o^OJZsv���)��#<[����R��Z���. ��M����N�O5w�#X̓�,�p6�Z�G�ޜ��jrA�`�OBUV��l���9Z���4�/�8�hq�r���5ׯ�?���UxHFX�{�A����(xz�uF�I��ڗ�؂�[� �o��tI�Z�$bkPC����eb�N~fa?vv�	+�_#��{��3����3����!*pg�o�yD����+�b��-�����Y9���maQf�r�&{թ�v��O���#�j�=�l�����=�A��PyD�A��I�����Bӡ�ġ7��c��(�*\I�L)ʀ�9^�I����(W���������Xp���Վx�8�����붡�"6R�J���:�C1�t��&�-q#ձ�QI�.���A�i�,��,���T6s�¿�Z���Y#�(�xC�z~�e��X�*���R(��/y�3�;�]ּ���{%��|Agɩx�/�N��9��W��ɣ�����NV���#�cZ�៌(I~u���HQ�f��mUκ�k@[ȺkC�0o�g!3��+wT��Ҁ-u���&�"K?󣙒�AX�R���1oȾd�)�����N-H���j�dv7o ��l
Ľ��@a���,��/�C�$�����h�be��i�3d��7�ߴ�`�|�Z,}�l`�:������S��nac8�D�I��@���z��a=�*�+�M�¥��+D�JS��N��xﭯF�د|!TS<(?W���2��U���ޠ5�|M�d!�
,�����|��=^3�L�6Ś�=���ɘ�ۆ�79-`U���C�)X�|n#r{[�/�Ԩ)�ѡ�-��N�g5(`�����,G�C�Z�W�s�4���?�EB�Μx#��[dMG����� D�,�DE��NS�AS�E��Q�.���.b�����*�۞�b$wq�s^a5�齤.<,������/~Bo���b�}��^rx���tg�$�٥�D��Ж]�U��T��-�\GK�q�=�'K����*���F��U=}��X��@��@L�O:�L)*�(�%={3���:��{y`%�O[�1�g�Wi���G�����e0���6i���b���ր�H'����Ki=oF�=8��P�M��>k��j�<����$���>w�z7A��t?��/W�P��ۮ[D�	�t�ј|(P~0x�iK�':^Z�M;��,j�� �=&ސa �yW�ٷ���J���T���~�sI�6,��[��ـd�k�Ԙ��|,L�c���r�f���Yc(+�� �Q�f�\}�/h�� ��7�~L���W+ Ξ#�d4���}%��l9�P����,:��5�{�>K���;ա�C�O{QeX9�tZ�	z�V?|8J2�kY��W�S��
>���Gn�P��~��b��V-F�t{x�Y
k��CT
�����h1��k�Z��[H� _O�L
N��1�E>Qus�
)B+���F"���a1��i�E��W���R��� +�r��+5�������P�]5��۸mV��������cg�H��z�MI2?PX�H��(�Z
{����Pi�٥e�[}�� �>�.!�<�6K�~��F9"��ڬ n��0�L�"9�J*��b٩�i��=ɢ,h��/�- ~��?b����PV�/6㞂���r�����y�I����a�=������1zj��R�N��M������P+>h@���6�@���0}�������7�a����o��1r"��f�2�冀��c���.�V�q�����Y܆�����Q�j
�9f��f��C�3#x-mK�L�f�PNȩ�ؔO/9sl�U05���u�0D2S�o�}���}22 �	���$:%��}{�'��t�.6���Kf6��jLW�w��nx[���<I�u����`�M�}�ٳ����$Sw�c�����:Lb��s���Oe(�ڭm`�v��=�ę��+AOBw:Ul�.'�HɌF��[{��?�D��r���&�H�oq�}b�E(e��(Ƞ�+U��\)�.D8���*�"֥�C���FC�8�W�%���h��t
��J��n�|&�^���_�S& 4;��3�d>����KÖE����ʗ	�U��Hh�o�y妶���5����2�w�q��*
C�r!:3 �B���j��vR��qz�6Z�oX�p��ҚJoτaj_r#�����ʈ�N̓�$���G�DA<���NNI�Z3�,2�e#��fH� �5�5 ���Ƅ�k1v���;��F=��S�S��4��D���c��Ϥ�XI�4Ǐ���ڡy9hW}R�[ yJ�{��~�r5]ϛbCc�-^|kT��M��:M���@���Jp�`���&|He�Q�v!�xF�������	!<���_+��1��oG�(�3� 0�c!_�����h;��?T�^~���o	���IN�x�0C��1��Ӽv%:��� S)��	�����;��7���ŷ>qϝ�;k��c�	mO6dq-