��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd92[
����I�	x�^�s�N����AO>OχD�h��$���q���y=����p�A��$
^�Fw�*r�T�-��0]�5jZH�&�Fy*ŐU�� ���9sԭ2�C�6Y�Iv���)\�A��F剑������R@�b�6�����U���n�5	��M��[� �ѫqY��Gs�D�j��F��,N�v�.�q`���`�?~�\�h����=��zc0�s��3}����Nc�Hi����9�����1v����mip�x]��~u�Ӟ��3�?�ȝ��`��S2@����u���gY�_�\�j��7�se.�{�b~�����QL��'�l��Ƿ/��}��1��Y�=��j�g�k�2��n8$f[��r��8�IV81�����U��oj�lJ�������[�Ѻ��3��N���i��V��_9�><�s�"�x֝�D��2�_X��U�O%���S�j�o�Z�y��}���_�v�&B�8��:Q�/}�d�
e� 1l���f3\|�&!��D�
ސl?n$������k���;[�J\�����$==�
�8��~t���xU�.�gD��.L|r��S*�jnJ���⊋�!�at�"��̆SEnNDą��Ja�>f8�x÷��ы|�q��s�i���E��,7�Ϻ1�+�D���թ��l���G��5�v�6��U���xuQr�x���]�/�]���4�%�EӰ�R�a��]������q*ʈ�=X�k���e�qy�晕���p&��얳PEܦ �⺹� O�8���\���q��/�����$�G�(�����]�n���\�8t�?Ϳ
8��C�� 9��l:�i�� ���#��� 4�dO���A��ͺٷ?� 7z 4��e���c��Z�59�:<P`�FT�s�a8XZ5-���OF7w+%���Ⱦ�M��,���B2�C-|m�� ��;��>�u(��-*���U��hi$��S�ra��>�0q��|�x/0Ԋ2޴}llq��4��hM���1i iTT�8\cD��u���5iF�����6�@�v�I�Z� "���D%I3;n�\.����Ȑ��F���dj�}�<�a���ܶ�r4p;�Rq������ ��4���y���O����LZ�7���,��)�!ÅJ�Q���|�
�%�7�ϴN��z:ӥ�>��\Fj��9$V��{A�~�>o�|�b|8U�إ�IK�Yn���9Zj�߅�wY�' a�N�?��[�Ȍ-�}̳9=~XOh��+�R���J3�TB�Qu�JK,^kp�bR*�fɚ����0���+��sq�2a�Է{ah,���pAO�.��������]v�=}X���1<����@�����^��pn��	C�5�+�ݮ�B4yNR@��X�v0���,z�9��?)�"q4�+ѨY�5���������X���]�_,y�h��p#T��nP<C�9�r܍��7��;X����Q��.���z�\���R	wc0�O��e�Z*�w���I�.�y�g��=�-��s����b�u�c������h�b���|��ـ]4��@��*H���X���xW��*�VTU�;�30����a�j�w7b��3�j~�m�ٯ��vU���E��	R*��$o�����Lh̕Aɰ'q��&++���R02�f�5�e9����5�uP>��@��ܕJo���a08\p~�C֫��L�o
��?��BU'l�?�;#���K���k[����j��,ƫR|iǾ�
#-�@�$j�nݖ�N��"%�1�=���Z!^��gf����k��w|e�T9��V�Uc���㢿R`BR��X#��rگ.Ph��u�"vi �����9?��Zx;]u��n1]k�V@�x��-Xr�`��(,�q�֘t��Cʭկ�������\�un�Jg��������Z�,.cP�(V͘�'JD�|"��4<ց`(e/"; �{��f��"�� ��FqBh~#a��)pۄ��G�,�b��-K߱�����2EN�M�ַ�y2�w�-.��k���ϡ�&-�1d*���|�D��f�,3O��-�x�4�m
|`JP�(�0t��_�[�3� �������t�� o���"M�+�gk^�y��<���􌽩T�ύ6R�Y� ?�hBI��Ԯ?a�g�A��ĕ����_��?�Vֶ&>N����/�}B	����� ���۷&��o�r��AS�L�_�K�*��a`V�٨C��?�X�e�9�3B���'F���$�P-N�X{�6����&M,�	;�;���C�쬒��r��j�!��.���X�&FB�Ҁt�Y��"��1�u�o�B����3� �2��ԩ_��#.7	�/`z < ���g�e���}�����Ӓ/Ao�tչ˘�*�	t]����a�u�q�Fd��-ٛC
� {��:bS0��s�T�Y�n��o�a7g������t/u�5�n:�7d�(LZ^Wv������Y�>٘45��,���I;P*(=_��2�(y��	�y���xp!��ջ���\�of��,��
��2�l��۬`'�ؿu��1	�Mm��3��N̆�+�/?���M�)B.�G��ou������C�N�
j�q%+�w�
Jm��o��(�GҬN�n@UNbe\�@�l��
 �j�r8x��PԘ%�n����=�&G������~��z!'i�ؐ�*�nO�FaL�Z�c��xch1�6X/BW#Z*����W���~=9r���Q�vd�c��N<���3C�&�m���}��O�T-޻1�0�h���E���V>z�L�6�o���3�N�� (�Է�� �1�8�XJ}x�ŭeI7`i�]�{�2R:0��a@����Ѣ�R��cH���;�"�~�#=��������a�t{���y����=�������]4�9ݟ_�A�m��o��>Q�I�3���*y�!�tqa��]��KI�n%9�6�2Ī	P�\�#mV�ߵ4��K��Ͳ=A����������m@F�[$Gq��"�����A������W�bO7H]@�I�a2w%�]����*����<gI=즩���b�w#��y������e�S�N�����Y87a�+�N��tw�fU���i]�l8�X6�����(��#hE���_�pY!A��iX��M��pX��B""��4�$ר�gt������|a��Oޢ'H�i��bnC���s�uD�/�:,�5T|�T���hm�u�������ů;�;gE���it�gE�6���^V�h�&l�%�Kc��=u2ۈ3�Z�2�%��������~G�3D5|M}S�{��f�� Ǘ~S��)d�*#u�0����y�>|�>z��܇�*����G[�-����4H�"��Z7���B��
Z`�v�A���K�NA˼�9�,�Y|�X�
�9RDW���GL$���+�)h}�2{����`�e�).�u<i��Ԋ��N��1�\�lh3�5� G�Lx �_�z���&#���%��U��+0,����50�r����:�Sc}�|���=�\��38��̊Ր�f���ӏk�����_&&�Y��.�~�"����f��������E������_*��#����P�B�|�׷��x��m�$���R��j*���:.*h�����Z}�T�[Ǟ�s[�W[��y��/�"�v?����Zl��,��ϑ�� 5��������w��I��R�����k�$�Z�RJ��B�}����&��F�#|�i�C��%��{�K��y���qt�UVʵP�W�b+XP#6Ў��>�<��7����E�?w�Ճ�!��
Z��#�e���@��X?�V�����2_��*�'�:R�d�����Jt�PP��H�2����[�n#��A��ꮻD/��&��@�����#�b���:����������~�en�(�K��U����KX�O@�Ak���vr9�P�� qæ��ȇ��f�u�ȓ0�C;���5�D���U�����ƿ7/3��oY�ҋa����l"-A���N-w�����eN����#�C
+J�?�@��(/�_���hcZ\>���6^a� ���:��~��]�<,��r����=�B� �����m���i	8.�`/�b{Ivfف����OpAG?}�f<��/����0c�����5$�>n ��MD���<iFa�R=�W��!C�]��9�??b���}��!�k0��7���\��!X�dI���{���	9���	�J��U�����h���b�cg�Qc�#d ���<:�x.3�Y����f1gK�!�g��-j���I�@R�q�����Qn��`�\���%��%4�V���E�&{�Z&'��?����:�Z�J��c"�ۥ��$O�����nh�kS���l�l%�S��N��O��ʫ2I��<�r�B|jK�jz���%k@��-#���}=Z�١`=E�8���q3�xu,��٭
���O;�AL�G<�c�����I>Ke8�W�F�m�߀* G֐�Q�|\Ta����q��GE}T��8p� �Sx\��a2�`��t���\\t�FEo>U�+��=D{������ѕ�Պ�1[�1'��0+�����ރ�;��p�ۍw���I����Ӓ�F�Mf�i%�Zj�W%5�{��7�A5 �z�{7�a_���R��IɗB�0c��[y-l�F����<x΅�H�8@�I:�2Q�@�ї2��eG<����A���iU�~�h�m��A�:�ٹ��(�(�{
a�W}��hG�6Bȏo�z��V�]J��� #X�������uߔ�����G4F����;<�b)�Wn[�+��,�ZȀ�"�Q���ad�dw8#3���̗����8����V�!x�����P�,�-���)��&�s��T)���H+�ߪ���`�8�q`�B��D�q�z����|��x2آ�nu2��Z��o�6������鵍�=.��-v�?��^֗$z�n�W6f�Xm�_8s��x)��,Q����	�ν��KK|ݥos���o� ��i�&\��E(>������GEdh�R
ӥ�����-Y��2�?��(y/*�-�F��9�)GN|��ƭ����t��R�U������v��b>_����GӮJ@��q3q��^�Q�Ay+	��5▱��*�贚g��6xDO��1�u�W��(��&vb��H�Z�sDn��ܮ�1v*�(�"30=ė��Z-�~l=�ﮦ�n���n��h�9z���3�y�܃o��~9ߪu۠ցIkg2�Nb��ύAMd�B��.A���E)�R4s'��zCC �CFL��u7���ysa�12��>E�ys�?
�O�/R�������+K!AZ��ߟ��!H�H
z�����21�msk�X�Se�A��V�r'������)z&	���@~�B_i�|�7JO,եˉ���N��Bݠ�H�:�.e���i~)r�/6�IU�Qۤ&�8W<n��.ƼMu���X�\�܍N��JFɻ?c��A��t�^�'z���k�A���a ��-nk��j�;��`N���l�Y�戚~M���"h�=5 пG�'���X�&����rL�;���$\���$p���n���I&~���T-i9۹��E5��W�1\�_R1�Ρ�C�M�0��'�@�)
�Mrc���tP�Ŗ���e�-_ʾC�9����Xtc!̢֬@��r�d��as>�̿�����I�J��G���=gAY,o*������3��P�G��I`������M9[�P˩���\@DǔceqY�_��w�@s�7����J�ºO/��wL8d &�@���/�E�����W{�f!MQ|{Ӻ�����mTx>ߍT�cR1�e_��=�@s�z�C���?Q�~,~��h]�����R�e��O'��e�~��ks	hh�ƣ��:$/����j��v��i&�@˃�&���ѠT��M��~fB�І4�p�az�
���_X3�o�Z��K�k����#��+ɥ��=Z��U'n�33qƧi�K�t�k߼J�@'��2�_.��ܐ�n���^����E����f���OO�^��J^B `�߯�ӡ��w͐�<�M����s�R���n�/��Ɯ�L��Ɠ�.�������"ҡ�����&�D2f���G��!!��Zg�(+s�I��(jM�6-��l/9�X���T8N��d�"Ϛ,T�Q�{������3�BL7�F��4'Ps FŔ�'*�H�mJG���}��]S��6�u�@X,�B{駣TI%տd��^��t�7�����OjD`��f��ݧf�(T��ۋ�]b�|�y觼Q@��d�Q�*�|��=���)��A��_sh4�8���}��a"7�V0YN<_�h���(�,p��w��0�
Π0
t)`g'�:";W'���|��Q�KK����z��-I���_� ��!'�-}[�oH
Iࢾ)�r7��`:�k���^ ���X��k:���kb!�L����q��:�Ԕ_qy��]d��r�����,�(�����O�d=g�
�i�Y���^}t���n��I~B�Ռ�KfL������("��Ƅ�d��L�e|��z���6(��kW|u <� ]P߈U���^1������# �0�n*�xX;�_�����0���f�Y�M_�U�Z6���;8ҕ�� 7�����6X}H��pK#��y	�b'z E@6|-Z�$s��op~x���:L#�M���e�v��p��2�U���O��tH�?To�F�{���y}Z)F�����yps|�
lO{�#}&]+����N��	�|�ûg�5��[��=K�MF,�
}�ʺ�1"Z��Yq�A�B�J]�9'��D�a3['f�>�����ߚ.,�9�c![-�K��<&��)�<�g��1���������"_ �6�C8�X�є��O=�	1<Q��6���~������D29�1���}V�ls
���������0�s�&��LC hi��"�H�c�M���^YC���g��}}:��u}�������:A �W�&�.ݸ�t2�Ͷ\J�*��6�����O�o�\#�g�$9b���л�P9��=�ؚ��v0�H�a��Up��-�������;2G�)����{\��E^0��$��Z4����8Z~n���X�q�\ǏI�� F<����?Ed%���f��	�!쩓��Lj�D݄�(�v�}*���y�C�МEb�l�3ge���؜yA�p4x��{�#��SȨ��r�;&��9H�?��[�'��2��|�!��?T'�r�e�<����s!���
7su 6h�ٮGV	9��f�cߐ@�L�b�����O� �GǶ�v8j�&�ί�����M�/��W�4��Ii�/_$Ǚ+ZՃ��4?2�jb�l��xԩ>}�lx��T���5e�K��1#*_n��8�D�b�8����M���ͪoG�vEz�ϹNF��f5l�~5">(�Іؐ�}��m�ѧ�Z�>�|q�=�p[�Qlw,��5y(�m������4��c+��#�0~��{��r�(X��eh�.��X�˝�7Fǆ(�/q��6�◜��[������Q:�NSvPN���]�D}c�9ܥ!I�z�i��Yz���z|�x�<c۵�I�k�5C�-���e9|qc�=�'kY��kO��3�8zL �;@���?͡S�ePrV�!t.��@nN��y�ze�&z.3ow2DO(.;#�|���z5Ģe�nLYJ�QP����$З��(�Ty�D�T�0�/�,�İ�m�/@�͇��B|�0�� Ӣ"VGb�n��TM�c򠬡(.�a�]X� -}�6i���j��]��-:�a�^��+�rN8n!��H��]ͽ]J�u3�L��G� �1�����o�	4H�R�~z�)?#ǂ���gELj���U����KY;� �������d`�va�,��TP�	�rgwH��k���2J���^���2�oƜ���#Vᤇd�c��\|5�{��0Zq��:�$QU���7�D0o�f�	zu�
����4_a/ޚ�;8�"�2�G�bA��[�#�oe����$��Gۮٸ�L��f�$?�*W0�I{m�T����4�����i�l�<s"ŋ�c}z�$�=��C2�h����F����&�E��<��(Ά!G�6��V��s��'d�u�DB,��:���!�\N��"T�V����w&n�l-p�V�l�Փ��D��&� ��?t�|}��]�.��ސ���q���.>���)UC��2�y���KJIG���J~	��`��e���M�S�:lw��7"��� ���W�!�L���l]2�����ʐao��܈�������#�Gm��YB��`$��Z�R��J[M"b�~��$|P��}t}R;�T(��lB<+Q��ɞ��C�WQ�`R$+�����-O��3{�]&�emE�}�G�pu���Q���)E!D����Sғ3@9�ޣI�,4��/�X�q��0o����#����\Aףs���7g_��`'؀-Q W�����
�I7���|ʆ��SĿ��ڬ���SE���_�d�g�8�ڸ��{d��!����/F���XC�TStI执ɓ��3�<��u2����;��8y����s!��GIf������Gdgb�3��9Y��K!x�����;?�e�S���o�K�w� נ��q�7�y�z�'d�4t�r[\j2ׂ(��BO�
V������6'@�����~`���5*�������Ԓkh*@$;�e �ƻ��隚��z�Ė}�@�k��:{vX.�sX(LVO;��p��3Dn5.��J������8+W��@�02�P{R�y�0�-asM�c,R��r>Gu?Iىo[�R�^M��CU��� α9#߷*�����;�	~�S}��I�@�%��@�-���G�w>���3X� R�Z��^B\��Hm��@}?�i�m�{F����|��� b0 ��R@[`�P���4PѢp�ӎW���)*���.�l����2ؘ���w�r=�6��t���No�}V�.�$���?������7�q���yK&�]ZJ#׼ͺp ���

)̠@��j�
�V���dj�@�C�@��D���0ȏ�Z�1�����GEM�t���[C�q�s2�v�׻V�Qi�X9��R�J�2�Ôe�~��Rz���'b!��";Z��<�yV�t��nI5�L�|a�Ղs���d��>�y/.�M��j<������� z�l�W�cA�Ȋ��4_�$;�r�3偘�����^4!ܘ��U#S�b;��D`��~�:�tCq_�Nc���4 yR��x�d1/ڈ.��~@��{�FԈ� l�E�2�G��$�K0v�ث�����B��RI�
v&^�b�-~����p�r���<�(km�v �}_�B�U}H̘i�@��T2��K�6J��j�Ч�Ek}��v�Jh�!�����#��6d�����ڀ�H=�ZqC������%�dtT�� �<�"U�SP��l�_�%�����X��X�.�`��<�6͂ v�d��c,���Ċ(<�N���	R�#���K��9#7ӐeN-�h���C���sښ{Y�q����?X}s�bS�bU}�����θC�`Zu��x8l����0���b�G%O�:�-�EȖ��G�w�⫝̸�:�U&�������¹���+���P�s+�gQ	�0lQm���n>�^�Hޅ)<� ʪ�J�O���Ҥ'S�L>ҩ%ѐ�G�&��0�׎��iB��9�8fea;��ANWVE�?;����Sܜ�Z&�EXc,������C�l�cyK��z���®Q+'���x��U�M=E������R�$�������� �tlT@�J"{�@���Jo�)�=V!��y�S,�GpZ�`�Az�o�Y�(�QE�v�bz�|3�<���,�(�b�8�hT�(<�]Y�G�F����Њ��'4�C(I��-�U-[����
��~ԕ`g���`_�&�`ˢ��jv���f�&��Z[�!�mZ��^غO䌁�]�i��B��m*t.�~��mÒ�ָ▞��N�f�0nGcB�ּ"@}�s��e�I�����m���ƻ�F{k
��k?��{w֣]�}�oU��ţe��a^�FcD�}�1��u۬��Nݚ��{��?�C
h�X�w��l�|��	_�{�����z+����A����z��ctԼϚn6�}��u������`u�J�=� B��K��DE�Q��"�&U};gR�붌�X��0�`�h%�z��V����o�uH��C���p6�?]v,�\w�#��N���sT:�,�(J�ܻZ:������B~�lF�)R�A!�[��R�In5@@l��f�x#?�ի}脱�I��K���P�ԝ���o%{ռ�U�}��l��aJ@+��-,]�|���x?r{���
PJ�4ؗ���[u,���Kb_�'�q�fN���w ��ky9���vb�q�A�K��7Ƀ��8��D#!���ש��ȒTď�A���Я�z�Q��˘��߿MG)�"!�̪V�Z�qý����, ��EO��O2�������ݫQ��=!s��]s����z*'K+�Ʌ�w�!�L��VkuK�n���/%TVv�S�|*q���^���5(f��a�S�;�5�+l
V$	�.�i���F���2��j��e�E<nQ�]���|qī�R$A�� ��:@�r�P��ף?�P��vJ�|Ĕ|ɛκa,����|�q� Yk���
��~#�xMt��1N�B%#�d��*�u�Ǟ��?��'�]r��8g��F��U!��>�j5w�&�H���yQ�p����� �4��u�;�`��|���뒈?��.6�U0�K�F)��w�2v6V#��_tc'�v�yg��g�;�`FC�H���7�;�5������`�pm_�\�$���R,����\㒆�^�y�麓q"��L�!�Oc��.�qa���L�W��}wi\
H���5�9�#)!��)ϭ�`u_�x�ˋJ\�g��Dj��ȖYyx?�������*<�Y]�n{<�H�����̻��Dۂ�e�^�Y�M��݄�2��\r�'��0�{䷱	X|�,Wn0���+��s4m5�(��T-$�I�?�W��vXҝ�M;S
E���Pap�<�#t7�%b�&�)+w���l��$sVc3�+Z���c��>���c|�i%�В�90ѵ�m��(��������	�
�Ҵ��Յ�bP��RW��%�ä��Q�hh ��@OWT'Q���|�NS��S������f�=e� E� �%����g�\������V@r+��9�g��巬���� ��K6�ˋٞs⫅ѳGv+?�rY8i�`��1ۥJ���?���3Ċ�K��S�ޜWk"���4���\�Ϗ��|��@��H�G�k.�Fk�}=Ȃ��3�1�	��saߖ�d���Һv�OWڕɏ�l *
������=m���nc�}�$:tZ�����'}=�ߠﱱ�B���Ai�|B�!���F�I�s����9~�B��~�-�j���gi�S������1##9MCfd7��	Cļj�6fg��!8���s�׃���J�ż�e�]�sw�>;�)y�{닗��L�����Q���Y|�X��vr�Q^�\�h�Y�
9��3g�ӗ[��$ R��ז=t������X�TԜ�U��D�aT�l��K�2L�I��=�X��'�
����|}��q_ѨĔ�0�����b�~-��,�hܤ�}H`��J[�� dk΃�ݞ��_��0E�7{�kEdd���ak�\�8�d���y�_œ��	�0adަ�)R'`>�Uz�!�Pk�۹�/��l8qŌ��W���YoBv������TX��TK�bz����Y�)�b��v(P���K��b�`���5�6��gY�wE�������B�A��LR�|��&�"�_�i&�� ���ALaХO��`2�>B���hSBK�%�r���5�dC=�ra��a�����:��b��!R����gB��]R�t�M���a�F�Cg��6f�t}�3�ZZ<r��)^QҰ��L&#�\�N�>�z�~@f���mET���h��fF�*�7#�����sE=�=�~Q�p7�l�eU+�Z_	���xQ�b?��2��e�|��e�R�kv�����-`!v���?;�,��e��>5��b�)-P��6'?� ��k{�d�C��mxo��S,���ш��2Rf/Y�ຮ-�t�����zH
��k��7|�����HN�K`Sˮ��J*iv̅N��Y���-c�aV2�r������������F������Z��5����4����;FO|bME���%L�J�T�jܞ��X�	_q�F4c[$�-�ĮN+ꋍ�n�%�jA1yf�n/��S�t�u<�gO�=��Kҵ�*&ԄRp���#�Ƨ���r�?��DT߽�[��MO�(&��n��ӹ��_|ڑQ��h�QIvF1L����u��h��R�ϓ�G���$��/�Klů�C�M���66Ȝ�<�fxOd��f��$k~֔*Y�o�2%**�Y8�\m־�U¤��C��h$V�8��U\�^�q)ƹ��c�u�U9}{��GB`
�`I��72ʧ�=A+�����[���YJ�n�)BV�R�|�sZqa�+n�o�ǟ�.���B��h�U����l1�����-ua�ݲ��n���:I��
)H��J�+�$eB�X�h�@Q�]���e�L�g<�������0g�(���FԞ�pQ�ŲR�Z�.���Ȉ��Y�[�o�Q�5�:�3W-g�	�v��O�����@�qֈı�O"��a��X_mY�m/L&j�⼑�ߧi�>�����(�\��5�h�yvΝ>s�s��̀�do
䂄Z+������4�����������k�MF�GZ_Κ��� ��0�$BM"�i�O�]8�Z���DC�4�b�K߹Œ^�uKjaHY��E��xI���yῖCsP��[��ߎ1c-*��i�?��h� #��\>���L#s�!��#�Zڨ���b� D_YM�=j���Br!�DƬE�%���g�8/iU��F<�� ���F&�+�j�M QC�DiS���B��P9��d��	e�2����z�yŒ�O�l�ȅg3	^*1�V�G���TJ��k��y(P�d��0s|�R�N�bG��Cx;v5^��짖��`u#�Q�;���Щhn�KW�y5�k[�D���;hۖ��y�Z񈸎m�.���H��(i�%�M�J�ق_Lf��b��sF*+���54'�Q!�X��֌������<�].��x�D���E~��9��Z��5M��O����pe	y6��tnwA/O��t57H����'�3l�:��7���x/~�XN��Y���/d�1MS��v�Ԋ�*?��R�j�ʯ+?���4$�40�F|l'��&�^�Q�݂�#��0��J����ϱ�Ɩ�f% �"NJ1C�����:�/Ay�c�_}�	�h���P�	�tC7��{�e��i�{����:-��7����k��d�Q_\p�6�|IjӀW�e_6���� �AZ���7wR5I\���y�?��������Z�d��bBfŉE��.�JJa��(�Y�x�d�9�d>kz	����� �u�ϕ�����)4���9PH��)#�q���w�x�I������P�)8yZ���S4�&2��,��F��ݪF�Q����Z�p�ዝh(��fsTA����G5�ـb�Է��tb��m���8	�&i.�k��En�ٹ&K���<���_T}/�U� V���F/��9'����	�� 6��61_|Ґ�٠��|�3"t��y��<no~��� �4���pV8���l��o����9�=��'��x��e�QH'�4�g3�[ɼ�č�Z�߽��5��l�g'��
�d�<LJ�����E87��myC 渦�v%��c��y�*Q����_3�]��2���@�/x�<�`iX۫آw���eNbLE�� ��.MՃ���R.�@�mb�t~t
`;�j�kTs�G��UB8{l9�]
e�੉�}>,�T��J�y��K ��CٯC焿(��QTޏ&`�Z�G9У|'{LCY�Kj$�h�m�?�F\HVeea�՟�
�ꢞ��ͦg緡?�Mj�%���'�Y�[߿6�X��J;ɠJʷ{�D���W����@���~z�#��n����<��e���b��I!=q�{��8Jm��O�����1�Hy�6�3-�r�Z@q�д���gv�¸�X�F����ցE�d3����\+:J��f��3�\�O�,+�<bH�1FX5�����gک'�[���SԮ��)Y��
Ѧ �o.�-<�KC�Φ<��\}?�0��>��Rr� c�\ޑ�!�S�s�Jް,(�5�]��~�:�gYz�&�q*�d�k%��f�~i�l� ��4>��$��?�,�;�H�����+�����7o�w���G.!$&ƿ������T7n�c��<NIQ:C�^"|sB1ۏ� x���1R/w�#\�2�qoׇk�����6v>��jd�i�K�g��|��y�UUZ,n���&���z�Tb�r| B�GZFwN���xW�N�;�\r�iq�} �t�73�M�*��_���/,�)���k-�����W���Vsv�-�p �}���
�sA݄�Od�[N>�t�ԫ��DO�����չ��Rݓ����{4�CI��W=͝xZ���Kvo��yDǭT�u��xʹ5��0!���yM]��.�$�\�&W7bA�9�����`1��To;ٙOs����^�Z�s�ӏB�NX8D��Hϟ+b��YM�^jh�>x��f�h�JO��J��cVV̰۞�	)���
W�����+�R�LP/5�z�i�Ƒ�\�7��t;Z��v�W��
>J<<���#�q9y/4�Yߺ5�c'n{��Ɣ�3��i;����Ԝ|X�����˓����_�_�ø�ƃ�!H��3����05PO����q���E	���ny# �>��q��m�pջ"3?C�>+p߭I� �K���V8?�e:�x��$(��#Bt9a�G�
�ıN�6q#x����u���N�3���g�]M�laO���(��Z*�&\@�]��G�֬�oCt-s��7P�py#�9}S+
'�TY�o���W�q	�^߫�s-��&ɖj��k�ţ
9܌G��m����Ě�l�p�Y\����u�<�ȸ3Fsi���;E�F�S������4kA�2�͐j#�Wa/0�MAX1`�A�2Apt4����F���͉��1��E�x�U�ی����Y2�e���5�~H)���)�r��<w?1 �h<er�t$N�V�	vu�-��ٙ}A(��L����1F�����N@fY/y��w)�X��]�?�����̩�M�>Jr0"�Ĩ�; `�J�NwbEq��Ke.s�1��l�}B���5��������rO��^/����Y��K��*�\�_v&�^�e_Z1نS�o+C(m$�f޴��dS������'GKߐ�]W���q�Q��5�ḕ��X���f�+�S�e�ȅ�Î��a8�5r^���N�讞��A�Gi	_�@Hq(��;�U����V��"QQ��B��WBh�q/ڒ�����D�"�2j?U��l_�x���I6��p=��)rх���R�"��vF��
t�JÆ��g�����$�GmG)e���j�x�0��"?��#(���i?��o�hʇѨ�8ܩ\k�� uu�Jp�KCw�/�v>l���!I	P���'���V��r(Y�����U���
���"�v���6�?K�	�����LAE�����<.�/N*�T^�<X�ɕ���-u��?�����?0k�L�f���|�Xl/�93����+F:����(æ�F����*,b���6F���oCu�{���?n��>��X��
��1���4�_>x�r���;��/m���^sC��<��<@��V��5�QV�:�֑��'�m�Q?0�q�����X��q坥��vzwa�&����IV��>SA�-R7��W	�%5���j
-�s�jM��
� i�9�y&��fW���NX���d��W�v@i��؂��Lt:��'��+�J��WSz��ܨ_�wiT-Q�wÚ��wT�P��G�1�XA*���i���c�d��a���A��`*�|O��R7���1��>g�-�p�HȯG��*�BE�[�|Ŏ�W�3-�쐫�����Pc5j�\�{��m}B��@�Z8��l�7��_�5`D3Zܩ%D�7d=9���Zٝ�g[�<�Х����s1L�?�~wV�4��4r�́JR=J���F� W�����Q���I�����o����X����I����#�D���F�*��~#���)���`"x��-q�@��zn�t���2>ol�R����g��Ќ��(ԆM1o�Ow�N�B!kI��o
���V��X�ֶ +P�pzҪH�,q���%L��
{����lc�BH&�wu�#������x�O�e
�l��}U}�օà&>L.�S"�V)�e�'�f̤�Y�����$�%��{��� L*P��k��"�`����o&!}/)�sy�B��:x=�S^�/��=5�/VS�T��is����-�W7IF����f9���D���+����cusd¥"(]��JV:�[����Q��F�S:���#����J���e�%�g�l��}��@���舓[��H�Ϡke�y[��B��@�/��2��BR��.�F|g4�^Q��$+!a&H$��A����"!E9�f@���>ْ�d�y�Ԉ�7,!$ALV�޷7��mƺ����P��;��)�H\=�߻��C,���T�Y_�AW�{r@�'F�+�.��
zv��/l�.��u#�Ō���8$c:	q�X_^���a�{��]�1��fV��z����hZn�
��~�G�
�J�OQ��.r�
�����t�*� F胘67b��Q��V���ǠY��]�V3��<_#�8]gz�� �_3����k��gf�e�P7;�q���'H{ֳ�K�^z�//��i`vm�t�b
"8���$�N�ٟ[�Ӈ��Mt/�1mg��%�I?�4-�2�qvO���<�,����<U�ƻ�0 �	������i'l��E��^��<��@aՎIbn) ł�;�\oCS1$@��y<��rS�stB]}0��ٞ�̴U�x���0�e��1zw!�n��nUv���KDEb
��y�=*(�:KsqL�q�!�c/l�
֫�9�����5�s���ْ�X<��$EU�s����`��&��l��ʾu�Lh��tl�ͳ��|����@Ϧ�������_��2��?�O��%b1Ӕ��x�S�6�t	
o.K�$ғ�l���k;Җ����Zh�X~��]�Hޖ,�H����R�6)�V
<��(��ӶE�!|����� Y� 髉Jb�l�:�"���I+.�\��H�	ܿ��$�V����H�@�����8,ine���'��o�s�B� I�;b�T�c���0P�J(��ix��+�{�j//T�Y��}cZ����d ��BS�����õ��l2-7���7�~ZgÛL����r�˴Y*&5���ܳ�Bѽ�ylt�D5��j�]p��Ձ®;},:w1��J %�|>���6+@�'��(����(S�&΂iW�|箣�^��f�j�YH7~�O��	E�����Ѐ%}�$ӣF�Kz5��'��sk�Q��|�e��+Wg��r�,q�|��y�46�7Xl�������'y��H��_)p�y������غB�?��'!	B`�f��L�>�y|��p�2&.g�'��E�����t,�*�AV�%� ���F���v��l�34@u6�w����$��F����hi���5�|�^��e*�2�h=x)w��ŧ�M����<�
6�(t�GJ� WC�ై�d�����U��'I求J��㵞� nS4E�� <��"-p;ʾ�����0�B-��;�4�).�/�o	S�@�Ħ�N�7��r^FĤ�e�R_� u*�s5d�����ݑ�
�Lv[�ET��cs�ka*y�����ksw�g�<?5��J��Í$O1���4�۸����,��ɰ -���Q��Z�ˈƭ�R�Q���j��{�}<�c��)�CjqLs��J�S|�V�r
(Q�\��w/���ifN����n�>��Ʃ�&���C�eU)����b�ɂ�1��� �� r�cd���j@|�}���*Q�b榷�ʾ�˕�*{��s'U�2�1'i��Rb���x�gյ����MG�A<zer��Ȫ�Z�k��:x� ��z�D|���J�vC�}+����8T_�?R��@KM�#��+0=��P�C2�8jN�Y���B7��8�)��OVΤ�`���q����U��x�%(��ʮ�����l�W��Z��7���͝�8��S4��RV���<��Ž'�<�=��u=1��'���%����+���!�C|�Q�C���P�<��H�z�L#�ɫ6�|'��?'3�����K��U�(��> ۉ��Ŷ�������a�3��ֶ�&�=���]؃�E�^_�VY��
��1��o+IT�JQ�Iw6���R	P�SdZ�!�bA.�) �ic�*M�!����ε�O�(�$�W�$Xȱ*O�'Z�I�[��~'r��,���Pb��W�:�A�����W�xNե�F����ێ�Z��M�%����"�����XՅ�"�;�U��Wu�w������\�Nb6���	�Yt�O��W@z���=���=�0J,zy��H�x�7�%+㼹${гvĮǏا�c�Ʋqe7*w�%��kq�raYIX���7�;�K�ݓ�^�\zC��'�/�4�
�5�`���H�h���Wު��`����s䧅y��á]�ffv�!e���k�NC��%�w�e�k��E�U��Q�	�Pb@l"�BK��T.->��&�P�e�&O4n�����H�?S��HI[Ax]�8mO�po�N�ܢy�=��%��Jj(Ł�rO'y2�4����j�_:��|�V�䉅3�k��PV��輝8��pS;Lt���k9g.�n�1���/�Jl���-%��S����5�e8?d�~���v�`���Z�!����]W� � ������'\LPe�Q�o"���ݿ����a�2��令I����r�x=�}9p�aj����n� ������1�s�.�i.���l��.��ߖUǗ$�SL�]�n!JR��J$8R��Z7_��إ����`S6�c�꿏.H[��^��qv��d�����\K3|�䤤^2//J?E$�4����x��o�A�+�u}.G��i��n�(8�dr7���'c�
�9Q����HJ��o������{S���#iBo�pFe|#�<)���1���@q��J���Q��~��G'��H8���M9!a�BlB�I�t� �^�.@(����c=L=2Q|����SkTA>Ǻ|C��ֽ�5��;������g�hh��U�_��w��u.N"�O}��$0�~��V�pא�� ������"zW|o��&�I���i���T�)~pO�"v7��;�Tw�U(u�[����mC�+�3NC��L]�"�\s:H5R����­<��DQ�
nD��V"�l�c����yv��v����[�q�g�<�ꜹj\��}َn�[8�}���V��.P�_fA=��̷_�;�0�Pvb��4,fKv�䰮�m��oq�u$[
�=�����8jT�%�g(4dI���T&d�Q��Nq��V6CrX���Ȳ��b;r�A{�>���z�G��6Q�gL79aT��?�҅r�_B��G;b-PR<�x�$�e:��4�5�ˣj8"��a;e^)G�g� ����u����AZ���(��e�8W��X�H�=�$���k7#�X}��ԣ�G
Ę?H�REQ�숕gt�c�?�:�;2�Z�n>)�l.�+�6y��j��RD0�������<Kעk;�����<��#$$�#�8��!	81������<�q=�b@��F�H :BdiG��!�q��U G&�`9�g�ضĢ�Q����^�b&̷��I�"N{a�=\��]�R���Ǥ� �Ða��G�d��j>�&)$��v��:~���&���`�sV�������5r��-�YD�����>�n�7���:�m�-s�:eU�O�����y(��iϦU��E�V3>'*ˣ_'獬�E L%�y�K����V|�D�(�͋Q����@��p���ך��A�. '���F��ط�R�l6�\������}����ap��?�b�A}K���S4݅��D#[rk��j~>�b���+:s�F"�h���ֿc�*6��fk;��\%-Y��K�o��B𲭫�6�BwʩU���9��@�eb�e﹂�C��{q,q�QԤ$A�py^��=P|��b��Z˰D/i-��ȷ�s/P͐�{�#G���m�en���Dտ�w@ռ�_np���\J�Y<p q��`P0_�[�5
���&G�:�%�;F��A�V������*EI�-;ʲ��͟�\��"4a�K	�Q�1!p22A��T��45��5R��դ�͝O��5�F��_X��Y�<��LlE�=�
�5� 3�RX`��L�75�pG#��ㅖ�����yr'F:�>|t���ީ��%����f�'~��`2=�ǜTԜHN�ˮj.&�����h����b[��O�#iq�uKB��u*��z����%>�������l�g,���3�/Ob�l�G ��!C	��>)�	�a�D3,�5��>�Uhl�q�U�}���YK4�#�m�:�	�sJq�ދ�ACYZ4LH��&G`��R��Rhԍ{}�2T�q��k�o�ח ����]
y��H�~Z24��z�8��2`X3���M�v��̑�gcN	]�����e�Zs�L�z��4��e^
���ם����fD�@�F��|� W-�, ������4��vY:��� �D�Үr�E]$4*AY/°�����W��9w���E��4��׆9��X��d6�D�ŗ�7��
G �������V�TO����U��@�H�l=\[O\��"OA��R>Feo��%};z�M��9�8"H:M��{Ɓ��l�߽l����}��t�D=�ˉ�6ؙ�lâ���Q�����TP	�IW��0�.Z�3L|��B�����.71I������I�t��̡
�`������k�I���x�rR1<��\����f�ڛ�"S4y���z��aG�f�+,pr��{����Q͘Y�%p��)x��N�z���p{S��Y�O�~>T ͰCY�����d.�g�@�$Iw'Ѩ+x7�I���mW9��<�T�o x\��~�Gj�«���ł�M��7R:z-Y	��m묯zzn|��J}w��*�wU���*��~�5���Iy��e��ȃ|X@���Do��%��z�BM������L�I)*�^�"~z��2��?�����	�)	�dj�b[3��7�#L���W��`�gP� ު��@��sG��N%nl~�U���������xAE0z2�z�*3�y�9��pN�S����Ia?�̕��S��L���0����cJ<G�q7�ok��o ��xȳz�;Ry%�Wrh&�I��I���m4�O�����%<�S� GM�ю+���iV�3?!�3@�p���9�Oj5�j�Z�#�)=�ɷ��D+�V'������Ǩ� `xã�XH�ۛ�.�=h���H;�1��J*Vl���0KJ��}߰#Γiw+dYG��ngf�eGn»��[��r��t;���X9�ū5�jM����d+{�24�!B���Di��e,�Ɉ���	�,�W�u�1ӳT��	u��yN����o~�@���ˣ���f�C�qA�O.W[�v��Z+͸ɡxG��,�>(���83�����@u��*�ej��Y/0&���@^���ŴP ���@<,�^�E�#C2���PyE�"d����NZȠ�!�nH��\��ˤ?����)m}�1e"��6�̠2U�f��b��nN�����~����Ɂ6� y�u �SNU}ݾg�\ =����QU���"�т��|���O�j����B
��ߌ��3GmC�q�)�ë9F���H��F<
J�L��2�=G���u�`Y�[�k=G��[B�FyS8�����B�^�H�@�,��s�K����/�Ԟ"7)����t�}��Z}�����=��7s�Aj�h�a(/s��4��X�� m[�V�5��aۘ��e@6���ەl_�ީ���N,�����d�'
}�`U�lс}����;\b���8��xD�'���o�����P l�7�n�XZ��G
=gd�hZ*�m��.�!�jp��vE�z���PCR7@��z�ȭzh��� :�߈�W���)ݸ1L�vo��9c��5���3�֪��;
=a8�Z�yd]���{�z��"1����PH���fq㴏i^�ԙ�/������J\�k�+�? �QЭ=��%<� G;��2w��8��^�JB/KF�t
��\���20����l�8���fy/Zw�ha;j�qm{�:<��b����z�)�P������k��[=8�m�z=��ب]*�P�۝@'�UV�w0j}wK6��۬=`�v�>�⭌ğ���H������AĀ�f$��!j����C;N�g�Z��`�	%ŹHc�Y����H���4�p�gq ��/�3��g�T�q�������D��͝��I{�[��<�,XQ�[$f���e�$���8g�����N <c{4�Z�;����f��ҡ��\��\\=�GL����*�O�j��LNx{:��������\/f�Yy�n�E���e�(j{92�d�sc~�@R� ��Ƌ��H�s�A���[��_�j�e�a��t���8�Y5Iqԥ�9yNe0�����>�kb��_t�ϲ�z��bn0�5�_{�Y�ߍ�ϖ�Kɲ����,^8���|W)	�.��"E�s�Hݭ�������{���Y�yDO�me|]ù{���Ae��OÃ�L5����ש`��GJ	��G	�ŭϝ��K�JV["�	�͘&8����/Rpc�Ν��oB�s�d~��5��B����T��-.%��A�����Vg,el3؎�T>����Nm:�r������8M(-�n��LZ$?x��u�N,j{�#��]�u7P�H���H͌�zE�Ug���d�.ѐ�7�^/��1�a/��⥐��"�*�ܞ�7�Z������y
�sk���!+<~�]}�s��.-FV�כ��h�/�
��m���Zo��|��g]ٷu<g��3�H�H)��
�^s�5�1�(���
����0�.��O��i�D��Q��cd�����ꦈ~�w�P�� ����/ .�wq�<O��+"���w��n#�qk����{؛��2��`αS{謞/�R��D�X@����N����+P@�^�L
�u����sC'�����Ϫ^�n��pr�\H��;-��V\f��[8KMfq���Z�O(*�5��yf��J�By$^� Z����YXkb<K��:�m��SÛؗ˔�t�+�1?�z�ڊ�W��r��G�%�k�Ka��ݙy�����y��z�%#�� ��[�
��<�_�.a��1G���d/WG���Q����W��t����k�5�r5��B�f�"2*a��Պl!��+$2.��o{�
�k��Ń��|�✌�`�`��G��+E�r#�$ ���V~v��Z��p*�TNv���m:�ܮx� 7��1'�)�����FzԘȽ_)�ճ-��6�}��-ns���2���v*sZ���<T� ��1�;���~Q�q���KF��(�1�Q�Bo/- @��i��M��J��-��5��N7ø[�"K^��Y���r%R\������O��Z�J^����� @�i�Ju1Ĥ��q��>*lǣ� IN���q��a�F���w�g��6�T�Z���NϞD`,�1�p6��|��N�U���}[�:x��|��E|�-wɱc���k�T���V�i�
ܬ&S���JD�?�d�N���r�>,5�Dj�ΛBs�HT�������vc���ř��EDN�;���z���|�/�x@��@�M{l�2k/L�ѻ��e�Ň��Q�A�m�Q���";�?Ԡe�������"�TÃ�̀}�;XyF@�H���F�sM��<���x9�����MȘ��"��l��]�oč]�(D�Tqƌư�ǯ
$`ٛ��V{��̢J���sc��p�lƛ��I��NaB�;�^�����ki�s5�~v�Hn�T�\R�Y�Z�P�Z�\�Zò�4�9ʥ|*ǭ���f/�B��Y#L���{���g\ֻ3����������$�ņ?�b�ӿF�B.("�Я���󉾼[���T�vÓ�uf����-�4�Z����� �j�0N�X�"��w��SHZ�B~�NK�2?�
��I�1tfx���߳(I�-[>�[�aa9��U�D�!�}�rK�������2�����m.���ԟ��JX���9F����g��"k�����<J0C���Í7�9��(ZJ��DY���L�7_~_��۫��-woѧ�׷��6�5�(�r�mDOGB��$�S�d�:��<�8oQ�tOB��4ˠ�		�a��UKȥ4�洉!£�|��C`l��vof1Bm��˽�(ƥ�钢}����8>���	��L5X&-��ńԋ���W3�08ڱћȥ�Ixu��@
�XqQ8��R��T������Hx�����;��[�u����1;���!�b�=�j�p�ŌI���;._fnс˂`n�搢Xb�mj�'���y�I'?4�ZXVkKϚ�L�d��.��I��nS�o{/j&��41ٹG�U���kz�|�jq͗�Dx���nCIz��U6�����D����`��jN#�,}���C���+��ו�"������ƚ���s��Ft-V=$�l�m	��|,��c�C��*������j���{�<�zqM���ݪ�(Q���ŭ�t7�O�&T/ݔ\%�'���w�e�ݣÛ�_�����)B��C|�͋�*_��SP�Z�O�b�r@>���!�_�#m����ͨЋ��I b�r�`�P��%��Z��m�*C�.����uPS���˵��$,��	�30<�/*�JP��$��~p:�1q~""�k�@nS-��}����J�*nR�XR�%4�q�u�4P�����i�՟������bb�[/:�v�l�瑶p����m��j�y�r�6�l&�.���JO<��@�aY��I�:�YN*A~��m���g��g��ǎu"<�V%X���݀�9�Ѹ,O��\t��i$��@���F�g�b�z�V���8�i�t���D��s��!�:��ɧ�?�!���vvv�8��brJ����戼�u�dX�8��@��1��M��~+�1�r�8�[�{���W.�T���p��9��-���L�:�Қ6e���5cL��p��ג�+�<�9�� �dg_$d�%��]�==�_x����O>��?z���BJ���o��S��"�j�>3�wO����S�!�����",C���P��� Y��'��	�V����l�i#��� �*�>�A듴���*p>������l�9���c��t�rX�H����.-�cy�],I��������B ��HY��vJj���H;o�CS�߭�����I�m؞^>z[��uw����Q���<X�k�2@����%M�2Ce�)隝̕[�R�/4iPZ��&,q���9�@�9�HE�[Mu�1i��f�;��`��%i1^w��pKZT�ˤ����w�]��ԟ�ڙ�6)�� ����f��\�dT�_ a	Or�_��*]ֿ� �B�L�4��y�}��h����`i����s�d�w"�n�9��)
��O���sg_�Q�/�_@xG-�E��Lwه��}�η0������Xe�j�^�'�̠��rf���*}[���Ӟ��!����4�l)��}���sZ|,�SKg�ݦU2�{����gpť2MfT��V���)Z6��g��@9�%��f O&��)E%I�Vb^��i�t�.BeF-~hy����Eu}��f�����ÿ�㐘vzuY�P�'��o�ݙ�m���[`�����0��>5�3+P�3<��`+�:�I�u�'e�$����:�ľ��?��=^4F�72@y>=0ƃ�D}�wR�{ڷ>�y%Uz����н^�P����iŇ�O����3EʢTy��}Н�ԕ������xZZj� :EJ�v34������7Y
��Hd0�"�
:a3��c!m��+��jюz�P��DG��yחe�:3T]�c��W�o����g+��@b��"�֍E�����WX�ƅS����|�ӑ���3A�_�en��У�¶MF���e���n�*�~���e%���Ae�0�H�|���J'?�ĝ{gt��;0y��K���{�ݍ_�Ͱ����f��Ut+������ �
��O���`�������S��O��w�DC���m�^�7��	��Bb���7�Rw��{���B�4E����T���F�9�$���h���]�:��a����Xu�����w")x��~���I��x�O���%�!��U�ю��^n��N���|�Do*�����p� c��m�w�(�⏫hHN2nP��#�?��%���V���`
>�?Hx#]�jU�.�Ym�����S&b��$�X������Gнa#�W_�-:���n�����9�T�j�Ȏv��9<�Á���I״>�_��-w�Om��w�3H��銖��@�X���]1Y��7��a�tNikэr��pp�+�a"i�qb��� ��$l1�|�.�M`����i�w�_�*�VU���׏���.����s� �U�0�$
'	���3�����ɬ����ZP�>��y	�#��7�&�ec������p���f���ba Lfh�j���DR�����{i�y��hXi�gw��y�xt�[Ǹ�_&tf+��F��O�x��>#�{�����7u�,>|.K ������3 �$�@J���@�9�؀'�2J�9O/�n�m:�k!U�*�%�k�g�oL�=j�;���ց�%�׷ex�=��'�1�l����?��&����@�3W��̈́��e3���ɹpM�[X�l�@w(A���f��?�(��RD�5"��>M�'mj�G�p"��O��!�K̇c/Z�;V+�9y�R�.f��q�jq�A�v� *A޹h�����So�s<�[sљgi���$ea�Aň|� �vTA��n((�H L������1!�fh�о�<�2���:�H�,���#�L����fA7�լ� �\�
���x4 �m�-Vm������޷j;Ꭾf����Ý=��Z��:�:�a�[�)���T�;��3Yf���jW��lS����Y�J�uc4Y�Ʒ�"�F����2�1��A}Ӽ��y��^��9wt��P[�ߺxC ]0��5���v���֮%_"rq��W
S�� ����j�bVÙ�$�5�];p<y\�塍��?!3�qrjjh��B�%�O�4���D/��u[��*'^����h��,pW1��!63U��0�0%��e��	�Z򳒼Yk��}Z�N_�o�Ҕ(dD'����gyJҥ��uzgrgG�=���v2�ʟ��ric�y����/=ÿ!�ž�Rm��`@���S������+q��n�yy����8(>�p���Fu!Է�f�=n �싽BBF	�GI�8B��f�w7����3��� ˔#z74\���A�N��[��L�-��ި4Vt��3���ʰŕ�Y��LsZ��T;���\�3fG�j�M���gg��Y��\1<e����]�� ��֟˷#J^��Z,���d����B%D;�CE'�zc�O]몴-е�*�e#��$]��˟�y2�@S���%��9հ�$�������pi�)����r�p<$���HN��x�nE��걍���%ina�F�Ͳ���Fextg�يb��@?�v��Y-���3yy�o��Mia����Ns�%U�qЊ}_��Ӭ�Q�{�˯������P�,�C�������>&t��"vH�.��K�z�"X�F�V":�`��"]�r��؁�6���ژ�UD�5�=ɬW�X�3A�kg�b�UU���n�\����-��1�Z	��-!��a,��=�o"I�M�P�����adW���|��^���B�Q��gQ^�ɦ����`Ɣ�V2���)���})����l�ɤ�� �9D��>*Ү�G{�P^F�����!�Tn��I���O���-�.*<y)�V���W� �F��Iw�8в3�OS�j[�'�Q�_�C���,���J�̕F+Z�_ǿǠ%��,e�L LD�o��B<T��o#d�6�����ʓ�<��⪢����Ȥm�P���ɳ�+�ZC-Fz��;[��[]�U�2�N���L9�w�$p�n���Շ��:~��dH�K����D�N��4����*p�p��j,.�I'�ң�>�<+9 S�~γ��@��*k{��`> �	�
��?��G=��Y���m�5~B0�ث���X�54�H�,Sm�M�=���=bk��X.*�Fhɻ��~�,�G�����\�� �ѧTO9&���N?wxI�G���+bɍ�� �p="s�̷�
 w��N~����?�f�k�<�����;%P��FV�R�X��+ҵ��{s��?=�6vd������Tn=���b�M�L�.�IT��O��:f� ���}2:a�@�Lz8*io�M���ʮ��f�(i�<��)�y�\��m�����>?�د�*���q�E��v�[�U�1�B�_�ʡW�;��MgT�?kن�+��V�����̾���i9�NbP0�q���{�����GDPQJ�[�r���G���6tm~�>\hv8ι��Մ��QV+7�{>OI`�k�Z@#���/�Y��P�u@n�[���x���3�	�h1Q�E�ހ�� D�y���R�`6i2�I�=� ��P}/���5v�	�TA��tę����"�7�-�ӧ���4�Y� :��ЅDM���߻-~�s�2�§뚰����J� �{�W۔�H�N�dW �s�?!&,'e���{"��j��JyR�,z�07��S,7����q����N}�)�
@rw�Px/ �['u�{�ʓt�Rq�!^Sh��;'�KWy��o~��>�%�p��&JMK��\��
���NSx�K'Of�Z���~GA�%H�h�ڜ��rOf�͇�8��Z@C�7��v�G颊�1��|��_į{����,ĥ�f8����X"� )��f�uڻ�Z����
;܎�]Es7�1�gZ�B[�
�BWl
C�Wg�Шtx��*z��#�;8f�5��1���>v厇{X�ڐB�{ƾ�N:�����J3�}�l�/. ,����ٲ���fH̅�)�?PTi�I
H����:���46ئ��PO��͸K��[R.`g�02�'sA-�,�7�'�a]��^l�@�
�_ ,E���T���<�7~}��9�3�z�\�p��1���6�R7�^�VxZ��R�ͭ��ǌ�����~�c�GC?uFK��P�狈�/QQ��!���3���H���?Ը�C%EӲ��B-�(M\��U%8>"�K�\��2��V�ᎍ�B�<��D5���\�MQ�$F�����X�>��vy�I:�^�Ie���s�{��@����P*��e�n�������	��T�R/D��o,�?��y0��*�����e���1t$P-x�i�ߕ����-�X?:q�f�z%^���CE������iγu<��&#�ұakOo�7%b���
�p�g�9�`2��H[j9���������cU�@+ɞ��=�z!���c�gQ����1a����Mɥ������ƀ굼��q��".x�IH{�G�|M���U��9ʼPV������j��p�#�2��,� pH�)����}��6u�	���󦔙�H�FH�.M�(J_8�Zݪ�G��Fz����Y,5�aq�)sS�ڣ��%n��y	�ڑ�_�+],5'��nI��3A��r^�-����^e��-�? ��j�ICS)�8�(LGU���F֨�����JZ.I?~H�0�$;���R��ܯN�mM�S����y��/�O���9����Q����Q皇��;l|wt�@uZk�J� �\�+p�Z>�Qr}��8zb�L�\IJ�#�HQv�(�2��a�6���c���"Ѿf��YuB�����B�����޴��d2�`�+�9����;�,�:���h_B�.�T��ɒ��Q�FYӹ�+�,���K�ULc���CsB\��wyt�s~�D6z4����V�G	����a�r�E����9�M7�D��� �J���<�l��C',Di��8h'� ,�P�+`�(~�*���\���I�_�`i��p�Wq?��!�5E����l��t@��}͎bf������T*E��"w6yY۪��B��(�B���1�(�GSF��w�s���Kl���Pϑ�T��s�q��N��X.EY|8�򌖜S/͖�6Y���#�\j��.1^��o�c���z&)̷��;�)��/��%RDK.�!er��J0q�"x��!���c-�.�c+`*�]���Rf�����Y�+���pY&�~s��i:J����zv�Os��Rm��@��_���o�+șP����ܘ��WN�K0��%������s��������X	�����p��Ա���p��"�	�a�R�I�y(A"~;��נ�r�����.Ƿ��&:��R�E~�}d�ub"�� ��cr6�:�u0ظ.M+��������H��� ����|�f�S�J^pzmԳ	�R��[��1ML\��4dU���AOؐ���0&���`-����-;���)�W'��m��qRq��ܫ#���9t:l�CcL,������`0ee�ո�CU���>���
���fb#�&j���3��:!n��&8�^���_�o�v)��>kА��Ywq�I.�-v��|�b'��v��]��&Aw�&�P�l�$�Q͚���W\��t��׆)(t�y��e/�����ET7���kڎ���\��=%�g�w˸8�.˳.�� d�P�t*�^��K���qg^�Q�U�n`�ګ��\�cN����+r���CT�K9�t��W��AURe��g�W'
�0=̍p��ɨ�lSr 7u� �\���k�.,*`�*�kNݬ��⥍(����:����$*Ǐx7ϡ��]Bo������������ޣ���f^}i|t���VR�@H�i���/��1:-���s\�J��Н�9�����J��XΠ5�i���[��F�,_�knX�ą��i/��t��q�V!:����n4>�/S\}�b�Ռ���ϛ����Ɂ��?�t�g^���ޒ����9!C��6	~�7V�������`�{�,���f���[0�Mx�dS����G(�^��QF��í��s
���G��ȳ+��O��s��O�3-��#�+JlBk�CH��;�	#.H)������r�s�T��\�Z��h~�[�1�O�`�������g<���ε9�*O���F�ҥ��Hz�͕P�q�N��HM,_���T������/C��q�h�!�t)��|�[%��g̚����5�b���y����� 1�����aJ�$~�Z}������ �4u=Wз8�XI�&�!<�.1�.5����C��$leG����D���h��� ~l�
�ՙ�������~�D���.��|��s��=]$m��Q�Iɔ��R�-���#�Q��}|��=�~.��0 �
�nv�8�:X�!�h�<
�����ŝY|7���]m��wkb�#�+|B�7��S��*�� ��?e[q#���)~�� �>��?Q������Q�lV�
ʐ����C{fi��K@��K���'OQ�v��{��?
c�]E�1,�o��`v��r�wMӻ�&�4�c;k	�����E��Hw) ߨ ���u��:�n�wȸ��t���:�MmN:W�9��b&��p�e�K��/QGc�-�*�&(U�r/0�u!�Q�T<"���9W��x�;	گX�Te��_�{�8;�cu�B�43_jGG������׋��-�ta���I�C�F]ӵAx"���U{�Q� ̹Ǆ��m�`U��cbQd��2Tðb�W.���}!U�`B��נY����l�C���8���\�)��`y����O`T�$ผ��!��6K�9���P7\��je�}4�G�p �}@��\���U�wQ����J������7����@�=i����_���f� ��ʯW������_����Ru./Z"<��ً*�Ee��dM�9�7J�&��3���0=9��]��`��
KT{�$N�"t��;�(ٚĪ�f��Zo�+P����N���ݑ�~6�v�y�<]h��~�2;�t�-�@���K�#����͋�����z�GP	�f�gЉ;��N4�,H~���r��[8���{��Ƣ�ljb��/x����qi���=��tp����jVF6~z��j�ϖmnD@9�3/��Jd̐��&��?�����b��̝'���v�&V����ԸSZj(LRR@�[�$k�ׁѹ�Aq���m�LE]��gJ)Õ�!b�5�.��鉙#l�Vc�~s{�g;}���GmaL�\�����P�(�zu�'��Ds9fyp�,�@mV�q���0���oU�]4�f�fYٹ�HeL�UN&�[���kS��q��]�Kk,��i�;Z���z�(t��>뇅ת���^�v��N
4p�N,�ʘ>���.&�z�H�v��9p�@)���<VYA��n�y$��{|�{g�_v!�
'�䫖Z�"�(K��=ՠ��+!�k���kʶ�dU�l�o"��وrS�=8J�}����p*��Zc���Q䁦��������p*l�I�%�O]}e��<���
a��oTRČf�M�@��[�P�)t��%A��Ġ�zK��}\�|dd�����j'�J�A�O�N�.�it����/C�(�Z%��u8裟+��J�����
�p݋���=����г�7[_(P9Ǐ��3�K�����64%g��{ݞd��VΪ���+eT�$�_�s����H���:�J���=�J�k��s�A�p�����;Z�Z�n�,�}m���CG���d��������+M��9T9�I��8gB˒��M�{�Ew5<�d����ת�B��2�q ;���X{d�[~�Ki!~{����l
�5�d2*��������c��¢���.:�8"�h�j�m3�F �;&�8���ڝ/��M�mG�j�D�kL�]��4�nSa�`}����6:�2��L�X~�#{��?����a`,K�\(T�@0s�G��0ס+U
!��kI�Y����7I6���@0�K����7��n����<�]G6빇���+R �n�H�T�K��eA�R?|{x�yP�
�cX��eV�fųGx��~P��*JRj����%z���4��7�F�ҔaǦ��g���M��a-�l()�dv�km+�
�	 ���+��ȹ\ꗩ&LO�Z�{�MZ�b�.e��ڼ�]���V���^:�\�z�E~b�&�K�L��8'B�L�*�s�C��`���U�'�z"�!h*]:�x��������"�y�fORA��ȮcVe_ǞH�M3��&�xj���u��;���	t̗���j���<N9��������.��x~A;�Н��6ݲ��&�y/��t�"#ң�+Bk�}�s�^�<sm��
�D2���|�u�����O�D�gz��m m��n*RON�:�6v�]�����'���I2O�ƶO�i$�:\�� ��'u?�A誮O��U��[<�W{B���!h��+UͰ�}%H�T��ǂĴĜe�؋r"�黪sO.@ �zP�3c������� �Si'�J�8;F���v6������@��@�;������{/�B���� 6�(b�YW�u*�V�?)%�����J�N���}p��80�>�sT���5��	D5{�?��R������)^%�k���t�<�T� 9eO��Q�>����<��d��_%D�F�)C�]4��:�Y �
�l�F�A�f݇��9h��,L5��{  %WI��9���� VC,M�QA���u�-��k��Ssֽa� q�=���w.*���IG��د���
�L����[��##A�2��y}Z}z��H2�:����e��V���赣���js����/x�-�`a&X����/>���&C"��M��������}pFQM�hZՋ���L�zPc��|��R"o�	J;�/Imv
\FOPɟ�.	�|:���i.Q�!��X �o�Cx�.Q,[EZ��M1,q��z1�|�_F���v��9�~����jc�~�6�g���AZq,D���Q�&xak%�%5��1��Ewg&�-��I�usS����:V/��D,�IWq�y�Vx��i���jL3A�'R �>av'�����//�D���[+D)�4ɟQ�PB�CES�nV���հC����Jx����<g�ݟUqt�����lƽ�{��Q[�Y��PZw���'�"� �)��o��Q����S����U$ ��[X���z�ihP�`��b���~��/����=��ƛ���:���������k���	$���k��kTS��2P��A��;W�%���5�����9wdrY,-<�w�����x, ��7Y��D��{d���Q�Ư�4�m��HO(>�Hq�<"@���5��ꌖ�#RY�dݑŠ@�@�{S��'�l������.��\�ua x�W[�wT�
hf��r�����NN��W��]��Jj��_���*�W ��CW�K�cu'[�(�����Wz�-�]�u���o�"���c2	i{2�����c)�M�Kc�0NwB�Z�}e�B�ߣ���g���1'��`���^�6��*�Z�˗:���y����<iӛ�7*�w�Q �>e�U��l��%a�c���G[��rMBe��J��	�į���m�t#�<���ڞ>���ٹ�g����J=�N��� ��׎A�����!=~�a��Ld�@�v%�Ҕȼ���J8+��6��x��˥vK��%["��mH�#�W�����e
©���Ga��G8��?�\��y�Q�r�nR	c��MP+p����Z�z�s<+<��2r��U�e^Zk5���v�}�$($ʶ��O���}��滛��>*z%�SR�9�t��9� Txq��˖�x��g��[4����xV�=z����x��0�lE�y�{��7q]����9(�[�.��-X\����%J|`����y�L��7~�T�C.h�p�O�ơ���U��)J:�GA�L��ԇ<"�k�#l��Ηm�t�Z��{kwF@��*� �.^Gd��}��x�o���U�@(�
\���q�������1GM&�������D�\�l�Y��7��H�:���V*ZA�XG	�u^�!�3�yd�L�/��b����Q3p�T`_3�c��ײز/�
�1y휲�J�LC9j	���sT<gb�t&L'�;E__Q��;g�8����.��Ȟ�#�x���К}��*�KE��1��'�=/Z�H����= (=1v�a���M���O�V�(U{ H�}xǒyT��.�-�q{�R�O4y��q���c����6X6�*��p���ca�Z6��7ͻ��cO(3�����@�<�-�f]H�)w�M����C�}�ῠ�"�SV�:ٿ+�Ò�y�p&6������,%�/D����3�'�pk;�Z.([��D���XpjYk�x���k�����y�7���s�Q{r:�ұh�v�ل�/̰�O!e�Y7��ݾ�q�4J�Iy�ѫk_�?�z��2s�m0\�r&-��`�V35�\�����&�.�!F]v/1�r�

�^���8G"_����Z��ĺ��]��rx	$T����d9m�ʔGE�5�$hנ��K���P�T����A�iC|�R�uco��;��]����_�Ca�����>c��˅��v"}���m[Rk9�3��ap�.8��u5�֖�;�͇e��K$;P�p�Qf��f/p�q)�r^Us�̀^���� �5��Qnen��O��p������x�А����K���ȒV-���8���8�u�{`�K}�q�/'�~i�M���_���Y�)Xy�+dBFi$�a.�z�o��ŕ��s��a��.���U;�����Ux��R}Ňng�@A������X}���-���'Ȟ`i��RY
:[�;Wr/���z,�*0������ڥ8	7�K4�9ѐ�X^������î��г�O�=��+[�������:����^t�
�G�&��d&��;z���#�Q�Ű�Ȳ�H1x	�S����yȓ�=�N�ZB��9tkW��V����&����}���d�l�-�2w�.����Ŭg�=PWc���C#g���r�� �������1�w�������I�d�[!�!;X�&n���'�2�3�g�i�~�@U8zPA��P�}b���}���6����E91*h\��%sRM;\�[�O�v���@s�ܢ��s��<3a �,��~�3(����&%��lǚ.�JG(�稗aE[�t�"�*B�������w�n��#�)��_CQR�����z�`�D�|��=�B�<���X1�y|"���e��5ۍ򎨲�r1OqΗ{8��a�7E�&�~h!Px�W�Z�~���$A�$~8	���(Dh�ś��D� yk���F�.��-�|HDjWt����:��J���q��-�E�D��L��|*v׫]k`j���}t	�_��:t_Q~�ۄXP���
q�m����g �� 2/V�ȇ���j�V����`�RxT���R"B1�&x`;�+�ϴX)�O��G��Tu����E�ӓ<�o��&�4�=�OB��A3�w��=_�Q��AQ&�T�4�B/���'���[H�\���iR����&��vB����>vqO$�gt�Jin���-ȁ�t�J�&2���i���t�6ڼ��#�VE��rA��X���s�iFs�9lM�t�a|�ˍ�;�{�VFj$�z����}��mr��l�HR<�h���Y�,1��fz��_MS����j.%ӿyǋ�ã�������Br��[X9(ݾ]�r�����Z�撸��4AMU���u.�`T>O䫑���S�mq˜�)�� �v�=���,y�T(ݹ�7�F�3X�ۑWB�3�V�죝fz��YM^:֌IX緸�:��T�:���F���+�Nx�ǆl����	�*M�Oi�&e|i���H�������`�r������v#�W�oQʤ��m<�����fރ�l�UZ8�w?�P5�k)�pnH��H��� U�*�B6����᧜�<K׾�H�-C�}�V���m[��n���_.�����<��3S'Hq'�@\NW�ǹ&F�W�W��H�O�&|#V����\8c��U��/O��B�M��q�lC�w��l�ȸ%b��g�Ƈ�����&�@yՀ��Y�}B��Ô��:N��M����wd�S�0����P��=5��Upo��R����,}��b�#��OqlH��6� Nw�|r�#D2���$�)y�7iެ��O��)��N�jB�D�1�C�/$w��}pJ�vg6��a�׽ ��r|��&��֒Alq�X��(�3Es-����i�.Cc8�Ƈe�z���O�좊����{�B&��R܁��ne��h�M. ����
� !3z��CE�zJ.Q��E����"<V�K����F.u��-��1���83� J�E�'6�����o�wi�^���8Z1w�eڴQ������̴9�(��I�ɀ�"��V3��-�WHN�ȴ��$î�Di����?���-�z[�"�atо&���yx�kQI�2�UX�t!h���P�/EB)��<�N�_d~�=�]o�qW%)zO�F~���XR�I��u]��z,Y6?���Vn1�
�O-w���TB-�W���i��2���=S3�� ��q{�q��AC�o�Z�s���i����7*�ij,�E`�B�瓌������/VP��4Ռ��ghfT��]���-�K�]�a��Ac�9gRe���/��l��Q�=��	,��x�X�.vm��������3�\F��z�uur���a&=R�*\H#���v/B�ٮ����Q�H �'Xr�Ҭ9a���&�$���%��� w�kT[�	�x��U���@!�C#+9į;� J;d�E�-ӌ����I�O$.g���m�^oU�a-�05�t�&J�_#��YV'�K>Y9��:�� �%IN��&~W�����s�8���:���O�&ؚ���0�}��b�sO��]Z�1cDM}����R�����Y~����a��Bꁛ%����"��4:v,�$��F�6��?81�gx��qw�#�gu�3��Z�!т��d��i=h�L;�,<�¡{����T�����*k5��a�I&�<T�!�ì�v�9&���ҮR:
`b:�t����v�+�5A�����6�7ͶD0/y��f��p�g� (��_�����F��lK	�EC�$7��<��d��#;�g���'jx�c�l��~(���>ys#j���Iwc8����Ss��K������Ƹ�~�J�*~�,���׬^<l�#�D)-�1a޺��{�%f�����\
����,���(�����Ē�Mє�JϞp!�J�>��×�o�7�z!; ���o�sN,40�[v�ª�;5�xA򔎇R�x�9���Ek������}ō [)�n������V�����b��D���� ��a���Q�#���Uf�v��#����M(d�Z���H��G�� 2|���su��H-x���s�e�6$Kt3�����f;cԊ�f�d����յ������~���s�eRC���ֆ��]���H�9O��+���]ʘ��L�=y� ���	9lL}Y0���,	0��w�t@�w�U�*�ޯ=uo�YV��( �GnvCK�����'?
�� �춫T�[_�-�!�]$�e&�;q2b�����?�yϏo�Uc���b�3�0Ħ�3|�|>���L���p\�@!	I=��dLkb��U�K���3��ʸ6�n��A����x�����'�(چ`Ps����W��J1�/a��-�:���W�s�Վ1��w���,�a�yCV���-�[�7��'��!�]�W40^�e�WJ�ef�ߍ���cvM<� E�����ߦ�;n��4��?,xq�	@E���q�:�k$�[������7yF�UV�	)�k����ې�D��0<`j=���w:$��e7�cJyM����E���Ӟ��\c��ڈE���O�PRƳmgi&o*�YA�+oa���ͥ&���?��t3�(i="aגR��@5B\p�\����	�!�wCk�=��L�Q�X�!�k���Q�`X��|�����&���Bh����7xsPͳ*N�o�
�_�2S.&�Ӵ�~�0\��� yר�J�����nPH����\��5[H�y����L?��&�Q�d������I�>ӧ�N�_"�Z�4zM)>?�ͻe Pz��e?h`�A�|`|(/GXv�w��9Y�;����χ[ow��]�U�4ٜaS�2_=������n���1JKS]z[\I>D����=�A������"YV���#���T_��cB���0iW���'=��4-��&��S�hv��dI�>�{(2Di(�*��L�;�Db�,�>�f��J�fއ7����
�p+!���D�,�����ɇgm��3��c�{���!�Q�,�0IW=��L�Mҙ�-���(�@G��,GRDq��oV=�5��.l_���gr���%����k慙�� �e>�y6���O��$L*�Jq�.��Iг"���_[���d+i؟S1m�v�Yziʹt�}H�-6��0�P�7���;,\�S�[!^˼�0
��*9	�w���T�7MCxL�&aЄ�3����Tʼ�z���Y>}Y���I'X���Ȏ��|���꙯L����y���v@W<�s�A����#Z�	���_f���l�}��&�'w��������?�q�~ٖ.#@oq��-�\���f�#�ƅE��2�V�w��z���0VbGSv5�)C��½k*k�I�^��y�㮗�~�a�[���b�2p�2 ��! �&8@r�㠊1�P��(J	��Æj�.{�A� Kr�W8as�	�W�u��u���e�A������/&���zDA�i*>�Y��(�Pq>4���C����ig�s�-�k�9?�f��:4��  Z���7�l�Z4YP�`�-�L��1tq$��C���`B�����8)+����mͽP���Ihi� 3Y,���2�9m����)�pB���}׷qى��AiE�J'G{�@k�Z;g���_������o�>�W!��X%�Ui��^�q9�L��c��9+��kVd9��$��~�?爲� c����W ���	��BC��<B���@Pдs�oم�k����l���UD������: l�8�K\%�Ժz�/��٘�Ӣ=�>�
FIgn�q!���Ś��L�#�ى#
�"K�1$��υ��CX��Ϲ�賿m��/��|�c�3��:"M�^����[�sg�3�D�Wůi闤(8SlY�{s}�dʪ�g�-�'�ɧ���F��&qJ����ų�Ƴ��N1�0��K��h�����k����Ʊo�:70���0��Snj�U������pt���{��>�Y�0T]z�1���o����R���>������D&QZ�\��Dk���Z��O\n�\s��A�����(8D�.�x��ɵT���\J��0(���Xf�v��8
z�َ����MR/�%vO��M3�-�jݰ�1�^;�
	>+l�ٍ�@��R#�"篰�y�o�^�z���jF7ɉ�����1�5V}�5>� ��� y���O<�� �5�ι��v�N���m�S����f3�`��ufs����K9����ι�uL��`�@�@8�A�˛�T4[��;UR>��MZ=�k��oѩ��u:,��1$��3~�q_T����O���-cﯓ^e�_G�J8�ې I��9�T���4n��6%æ�\x7 ��1��Bl�gc�<gN��7�jpZp�Yu7M�cM=䯢BPM\n�"�0��8��H�	�	v�� �	�h���s��ӟ��m�����7�8��/:4Fɸ���X�e+mŠ��cV%4���/��0��}r�RTd? �Daw���@�2���t(Q�A�OSX,"�ۑ����Mh ��;�E��T�L9�Y
#�n��M�,��b�����k�6��y�����*�oe�H�7X�H��������ϘSg�`��� ����V���n;6FI+mnЄ��Y�ꍙs�OG�d��4�l�o�Gɔ?�T��R������&z�P��l���MT���$���/a����9��lg�%1*Baf�FJk�y����p۴G����p*k�#x3�k�5oC n���|`y+�p.�	����K9X�1�W6��8�J��Lux�O��4ӎ��0�~1��:�MN������II�{?�Q0C��Gud9��e�8Lh�.��`I�(KV�wl�t�\�+䦨c�%�B2L�X��֢�/�N�Y"tGd�ZQ�ob��?;�q�#N>w��{�@~��IU�2����i�y��7��~��n�&�S�ʻ�L���1о���ӗ9]��%UKX�
��ޥ��4-E
�C�cR�]�+��!�TzЇ���>�s]�K���3�z�aJ*�U�F; $6	��HR�����{4/�ٛ�h�'CD�ǻ=���H�P��揖#�s����j�q ^>X�7Lx(�d� �`��>��o������P�Q��m@�0�NOS�^�ڈA�4�RJ��}��oU�.�2)
��IBG�� w�F	e>4�B�u���S�A`��3�	���v�>�]:��k����W��G�kZ���Q��-��V�$�8��c����ww���3I�=�{o5�Ԃ��+�qKU ;q{05�t\&V�Mk�2n]`�ޮ_ʍ]�U�Ir�(�R�M�U�������^���V�T|�e�pr?%�3�5�(�.7a�pl�֪�	�_�9WtŶR�Y>/�o"��$��Ⱥ����fG[�f����D%�mq:&������)ah��WPad��X�/X�O�U`��&��|�W�f(�ӵ�o��v�M/�����$dm+�]熔����*�Ld.m�_�&I&�H��2n��kǜ���v)�
����%��|q���OӋS�@:��X�k�t�B~�}cW��b]�iq";Rx�frrI�wNM+5~(�JD��]�K^�=���#���i>pCRU�ohݠ��� ��עR�:�J�|G��D2��i$���X��z�*7�J�;�k?ͩBF�h���<_r 5�R{����s�6
���_���27���?A1+�;����[z�&0��s0�G��l�ca�K)[�K7����t�X�a.I_�+�����f�lq�9�(v�����=�<��&�=�'��o��.W���r�����~�C����b�sPQN����k7m���lw�<�9��>��v�J��!����nn�쳡}E֮��>[6Nqj%V&Xշq�I�B*ǍR�wf� 昽��9��\��H�J~�,�Co�)=x�Z|��u"��#�(ٛe$]/,ǻ��F�{��  �[n�I�E�FV��8#�|��66��c��w����k$]�~E�`h���1ħ�������%ǧ/�}>LX�DQ�2�V��7IO��Y`��_'��|�����X��"����~���t͂�%*��Pg;�D}��	|pw��,��^��Qi�9ڙ~��w0Y��%�#�ϟ���%(��, ���~��'�=Z�����ؙ;���{T� 
	�0��:%*0ӫ���)N~U�*�"r�yz��L�`#���܅��P��q�E���.�l,t��"�jI�V�lN��fپtD�+�n	�E_$��c�D9SY�㸞a���09xR�P<��& �krp^Y�V_-�D �������Q�3����-.�m3���i�G0Θ�GP�yd�2��pg���jy�L1����Vf���KDi.�@;-ȏ�vh����Fj>#N[�[�6�lr���H@�N�~�{b��b���/�-�%ϖ�A��R0h�Z�4M�����{�8�m@�h�2j��cS1mƗ;C�ֽ��@�{�,��2P o��/�'=&"��զ���r�Za��U����3�o�n5�I�%�7ǰ.�.q�Ĭ�gB�T����r�[ #�/�a�$m;ڔ�=�>�}���;ލvXi�o�}�A��&yU�V�rt4L5�s���KXԊ/횱w����E�Bpa����މ���֏��?7�Y��,���D7E2�z|���o�e���/:'M��\�!�&w�����:��U�ǔ��n���	��c�<<4�0����2�uHb���E�~58Ez�S�1��SD�d��4�AN�Q����l���)��"Vm�XE{rw
,�դD���0�&!�#�|�� b�/oz�a�=�o;/�j���O���Ph0�zl��B<lZy�hs��F$^��:M\U��+֘w,�(�.P�4�e�b��I`���e[����悑��_҈�Vĭ���@���7�5�(��A �����sL	b���w�n��¬>e�h1mn���\��9���ɅHI���(W�r�2���X�-��-��Γ�6��c�c��+�C$B�I6T�������t�W��?�s�b>���zܺ��y<�Ӥ�s"��_e�Vsfa���x�Kd.y��붥����O-��U�٣3�3)���) [�j�̙;5Nl	������3Mt7����G���}t7��8CA-"�S�2� ��H�K��모 ����y搚���>�Fm#��̨�����Mb�� :���+>�](��?"��In��ֹѕ�$"��g�7��Hο��b��~���DS���}9�hA�{��o���u.޹:�r3�� �1���T��poǾ#XN��0�O������d^�|kb�an��08X��8XX��=YxO��T�~���\���_ҙ���ws�]�P�Wy�w͈���yE���_����ZƇ�82×�N����A%�ͩ����M��FP��
�HB����2�.��bV#�$v����/���߹g��ܤ~�d� S^Q��y���.?��;��tc���p~A�FL]��3R)H<�fi��N, Quy>�s�^&j�Q�M.��a
,!Ai�Ѻh�&.��Eh�0ؤC�:����MN�w��7����L�TO(ݘwHTy�ƅ��uG(	,4F�nmo�0]լq���dH����W�?��������I7�2�����E�����ӎ�����M�3,o�3^���Z8%5�]��UA4l���,}�}����s�O:~��pv�߹T���5����|�?�������h���Z����� �v�LC֣��7hq�_½�,�w�X�+�M"�� @�?�X��N�+�j"(�>����^Y���d,�����F6x�é�L�j1Sm�hMFW�m%��6���x�ƽ�V`+�Ҁ\=a1:����u���g�}�I���A�B��o�	�+a�Vo�rZ��A��h�7�W����$�uэ�<ج��	~�HX+8�.�Zq@��=�����6#@[��&��'T`1��žY�W�V7�
��(�@B��=�B��Bi� �[ܱ�V1�!ʘp����c1!�v_�Y�C��y�w$��M��haؽ�H��� \���k]͖C�I�vwձ� �D���8��dc@)�
��[�Ż ���?ʧ�#���E<��8��kap�*�$���xt�; ��#��-T9��i�>��(��߅�=<}~��1��w�z�MQ;ن����6�!�ɺ���f��Qs�Wv��6>*Y�;��s*�Um�mda|������Į���t��:̡I1��������z�c<eg��?J���K��T>�_�1D(U�_a
y�~20��S�lrR}��RH���$I���~%Asl���S�bٻ���x�(q�ʎ]Rek��8�P�g����lz#��讧���1��)ET��cD[�Z�4�<��e/��?���mzHmݚ�E[�8�s���"N?w��B&�hZZLx���p|���rDRM�4�]�A��"\gA)�H�8_7.VD��ZO��������r�j7η){j�K`m�T�	?�������)=Nؒ�ɝʳM�^`�Ӂ�#k2N'-y��ȩG���oJ���>�`țV���9���M=�2���������vc��#��JG-�¡�D�)�#��Q��W�{�I�����U�̣ ��ƍI%�v�s��*y�:x�
!QK�9�U��D{NwgxRW:+����a؇��(BK��YsKo�g�-�a�+}��ny��&䕁�Y������ͨ�i��|gM�@TѮ/HkBL(��sY��&x���s�0��w_-����"/�NR���+�0ʏHL�UK���StB��>4�Uj�:��g�~2XT�<iA������5�d+O��@/s}6*��\��T�Pa�c������Mh��2�#�'#���	G��#*b���Y�L-Ob��pM<��0p�	\�hj5\�Ĉ��?x�>�y=+�\�y��g+l4���N&;�"�����G�H�+�ݩ\�l��*�Vv�r���G'��mp����U=�>�����_D��HȜ���{������V}3La��.ߘǇ.��+�:�x_Kֽ��tϴJ��c�Q9p��>~j�ຐ]<-����%�)��q܃���`SM�d�nQ�e��l!�h�VLm$i���q$C��>�wP�tL��� M!+%�xL)@��<3��w�P��WN�!��d�����Qp%U�<7��Z��o15�,-̧���|3��F���Ig�i;l�cnO�ڋx�l��{(�D�5ʲql-�)�qh!X�(�#���S��!m�
d��7����� %i��L�gM��y/�������8K����!�a�/."���1jb�����X�9��Q�^�][��@��dD��H𸬲�An��%d��瀤=r��pZ�(��æ���3�M���|K������p��-��[K��n��y�ɀf%Vf_,��]��+�슷����EC��p�P'knA'�d5�+Ys���o�n�3�!�\i8y�6U)<A�`���G�A��9?'RW�JֿW�N���ъ�kq��8�@n2:Vv�|^èt;]�#�/��`��K�o��ln`-b�e�Kḵ3\�vi�
<�6=����U�C`z�v�����I��L�0U �6iMg�h�[�k<���V���fSmusz�o�*�!�"����Ӱ��<'�Y�؉��:"�N�*%�`�c��ֲ7A��*=��׳j��5��q��ط�a�H���kJ��[�x}�4�CjE,;�l;�U��=U5-!�Y1@�g֞��;I�AW�\�X��8������ҕB�;����j��Tw�]�쯞� �����oW�ۍ:/`z���A���hqJD�u�o�<`$�M�
�~b��=�E�&�T�/�|mY����hA�]X�)a[�(��1�Dw��B~
ܑ�ZƱt-�ʫ�e�"��-���pn�AGoc�­N�)���G��[v��-q�Z����=9c�����7�Ʌ9�W�������0�]C��C��(2���������;S���lk�p���@/�i��=�Y-�;�q�hЯ�<�i�8ڝM��S����dD^���`;�ND5����Y��� "�%V����'
�)X(ީXT"pݥ7������Յ���&��ԨC�gO8��'�e�Ujq��c��/+�Q�ZJ��<f��I��`I=g�ڟ	�n"�{\>V#Uh��Os���(q�(�~@���3n(�]o�Nf�kJV��\ӻ.h_��9J�m�m���QR`����وL�Ad1sK��ϫaӁGG���s�x~9?�$����������Ч�c.)1�	�����ϐ���_���D����a���
�ä��"B� ��C-ԅ�M�:rz��s��X?�٤��Ej��P��&\��;2����m3�:�<)p�f���W�E&&��!2�N�7�B̭ܶ�9$}<ޓ��������ret�w�!Yۈ�{M����V�� r����%������$yJ[�PO/�"��]VM��\Rry��������c ��U���Rf�1�����J��a�a�,�uȊ�O�|ط�͡�a�i60�5�fK�9?�Z�`^��X��ŝ:t�Ͼ�S[@vIw� "�w0�bJ4S�˅�AX�����W�ʸR�'"�.0��[�;�Tj?o���j� �xQDpC�|2#4�r_���G�sk~���r�	HJ]��x����&���F "C���j+b�4�!uZڗU��	��������^�N�x�{:�]4�%K�� �C%�<e����7N�����T��N����DJL�ta\�_�Yǋ�v���~%��X�w���ʙt���_n�Ѹ���	�g|��]����Jr"���ml�N5bT:� �M�Z�6AV�P���T�� �w!�A�6��~[m�|�?Fn
5���g�&4Y�T]�1�IyD=)7��aG�ꅮ�q�"-�۴�w�p��S�XŔ�*=��W.�]N��f�,|@�W����%��)t�j�
���l;Ɋ��H���t�Cw�\��BHu�f��Q��s�����觚$,H��h��*F�U]*���ّ,.�?z��6����Z��+���<�?�Leš��e��j;����+]��^ƒ�1�5o'�˟�N�����n][�VQqH��}�6��i�B܏�z�[t�:�s���]h�����2� �v^o�����#P�]�ˬ�sE��t�D� 8���f��߻B � 'H����æn��"T��9�>.=�L&)*xy������: ,���M�9>"<>��)c��vI��B�p�s:G1f�F��/[;��b���Zz�(����Ѕ����I��Ȣ�?d�8)�"���wԪ�n0�[:Q�Q$22�Y�%]�ET�Ek���M�5N_�5�ex�2�Ƞ����JyU�W|4��k.P����Į�8rf�͎�7� �p�FV]/:U{��H �Tw�R;N���Cj�=�[�'�L�ğ��)�5���7��G��ghv6�蠑W9]7qH��"���Ȏ�ݱ)�#��#�ց�@=�J��D���K<�67�z�Y����?tG�|��k�)Hv�<4L\��.�3�*LD���@;���S��:7��0�z���VO��j+fQ�Ӳ���2wf��� R#A|S�0%^�Ъ�"�8�N5��4����YXT l��~Q�/V�@���ƛx��`z�RL˒�nn��k��Z�QKe����r�Q=Rt��ϩIrE��̉�WQ�swz�	"v�Yh���{���]�Vl��hD@��A`A�����P���1���#�5B+���X���ײL����{��FE����6��ǈ���G_�֝��u�����<�V���~��
`E����}���:������~13�����ɂ�|a`�J[�&��[�a7X���~��k��e��;.�V�Fa<"i2�������A���`�
�����������o����D�:�����B�}r!�Ʃ�0�-��7_���+y�#�O���ٶ��V���!�55/���4�̞0L5����u��v��4<�!s�N*�0ӡS[���Ǹ�����gC)L(�7"��l�����7�	%���&'+I������p�z��'�hqH��A�����|lQ�e�b$${�����ȥ�q�qM�K��v��m����(=���-\�e�C�8$�|D��O������y&�I��dNU&�����¹+���p[ѽU�H. oA�{�Sx�Ȭ���_�(��tYx֌��,)�XB�/DUz�G�3��f�a�z��gL���1�W`	H��w�l���:��e��Sc\��ʮn���H�Y��_ը�YRy�Z�,��I�耺��sI_sKA߀M�; Vt�������������;���?��Z����%i~������^ٗ7iU��!EE�[���~˫��T�^�t��A�釤)���C<9��J���ǾJ���Hh宁X�긾�[�]�j��� Γ����e����g����lЃ�ǳI�ӏ���/R�h��:v�ć�Cb]�2��j��~��b봩��ˏ�_�l-AT�uV��Ju�0��j Fsc}��B�TA�|��̺ן��nK���C�m�< E�u��x��)�����Pth)j��(�]�}؆w�jؐ���X���h�F��UA�O5��RF�~�����vA��6�'��Kv�MoY5�w����h���X��F�s�9�����F���K{���W�P$O��c��$��I��v)����׾�XP�6���e�Xō�P�q.�BE@)G��ayB��{�|����'�ח��l����d��Fᠸ���/CR�oZI[7�P?�,��A��X���4����%e5��g� �`?��r��� ��@��-�d7�}�����3���(�����;����؍N���in�$
��#�TK��i3�BnV����-���6�GP(N�n�fG����4� ��ɰyn������1��~�@���w�_��r��f�*��KR�?��i8�]J�:��
5����p��J;�,��p�'�`�X�.ϓ�T�e" �m�	�+�B+C��w��_�c1%y\V�C��c$8<8G��{���y&�\m��NPX͋w�74ɨ=6�HUK�%~�qAZ���:��d��8�L��ρ��l54��/_��gaO��Iԙ��ˎ��:�*�����x󾲝i�Y~V;���I�*#B�V�Iv,j���g{p^f�؈��t ��ĕ>����uY��n�W��:Yrs=~���Uf���ϛ�P]�F^�&�~���hx(5P��� ���A�It�U�Pqnl�k34̢̓M���KL�C�/���{�g.V����u������>�i�-��=�W����a�:&�rK���'�`�:{f���7��14�u�<![�G�{���Q|��ާ�{�2
���D�|
�G���O!�K�1Ѫ�xU��s*:�J���
�[ޢ����Ɏ@�ْuqr�&C.&��nIj�� %�0�W�8�'R��x��[�đ��n��LB������.�q�B������B����h�6H
C��Eg�>�|�A� ,#��ڞa��TF�;`�ۋ��Xk4�%)�����
��za�\�W-;)��ȹ����b�oJ�GY?�F�\���Z�� �P��Oȗ\p�0PHQ�׮葒����lm���&�^��8��T]m�;6�L 

!�ҸC��ޢ*
�:��t�Y���Q�K�O�/��!3�:���*�O՝�н+��#��g^uh�|Eܵ��V����gM��7��̍������Q�~)�7E�H)χDV(�~�y�]���!����<�� ��F>�ky�$�;l��A��1œ^��B2������a�q�`r�D��u��!�<��阯�by=�:�J{�!P�>��!��}�8�ؖ�7$lL�4)\�˔���f�N
�̔�ը,8��t�!I���2�&�\k����_`����(�k�q���N]�)B��>��"���0Kf��Ӳ�L��ʤݯg�����d��"�*GudQ��O7q*!�����m���D��}����j��t����2.�}V�p�elj��4���5
���Ė�&�tv��U>��P��Kj�Į�@]4Ek����s:)أ�����6�ّ,��r�U��ڧ��6��P8h���l�$g58@>�npkXg(~�Yd��W� !�q	�.[	�|,V�&�  Qv�\��Vh�必S��,��"�;���1�>(�iC89��s�)�t��xX��n]�d��Q��>�&rd��=�\&�]p����J�#☆@���7�BbPcn���#����7DgS���K#f�����0ݤ����9�Є���`����w�%��	p^#U�i�?��:��v��] 3�;v)��������t �,�܏�f�管?�'К�4$�i�#�g�Ό( ?\Qb��ޥHzQ���}ԑ���������ܱ R@����ki�L�x̝���
{"+Oe�<�57��2mTLP;܆�qi֐C�I>�-���`�B��,�.rԅ��9��p@1�yQ?n���G�q3y�	r�jL޻��`���	��^��o���0l:�U���Ya���z�^A�^��*b!�t�����A�����h�2�y��T����s�ı����3F�,���.�A@}�`'n�3���u;�?�^ ��Հja�%U(�`uT����J��9���4U�����d�T�k'��9���:��63��BA�ׅB����/��!�~�p��� ��J.� ��gT��|��VG����ס �]��w������0�$�A�!=�ʠ�c�63���ƥ����˹�4C��by���,�@��j6{�o����=ݽ�iE��mF�+����i�QX��~%����"3�ާz;�l�����*��)w�m��Чq�ɺ�1Ng�r�J���1_��_̋}�-�#S3*l8߯��T�+]3�;D��y9Je�?���<]W>���e[��W�v�;�Y��^2XZ�~��]�w����B�s���j�Ee�������e��nv�������g[{npV���>;_e���7@�vR �՞��i�B@�_�!,ݩ���l,1�Q�Fy�І����N�]Y�%6J'*�{�,�B����	޻���h�<V��g7�*�.��ށbΖ�