��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�Ǖ��[�K�S�%J�L�7�@qM��M[�ߎ(��.��8�M,�t�e�r����n�9>���E�Fjo��g����ȋ��T���\H|%-���?"ӎ_؝dwƺq��[��7'��P�t!G�3R��Ϻ�<���j�L_g�z�ݝJ7�ATD�cs�⦼CXXjي�v*��Y�n�"���P9����E�<��d��Q��7{[E-ý0������^,K��i1�]�q��:�(��U����^�d��)�i�݁`���"�~��D(qav�buZʍ��@���2�fi�|�ќ+�~6�}�Ղ��{�ʱ�ڼ������ܾ.Ϝ��Ƅ�;0+b<��gq�W��41��
(�,�p���%���j���k��K�a��J���Z(�,l[fj�;�J���Gm��m���V�� b�{dw�̃�?���L��mʆ���9'�9K�@I��wf��k9j��d[�x ���l=srEba���f#�%��J�2��*��ezL�8���#�ut0����@{Cp��Ys4*��Dro�:ݘ҈+|��њ'�!SZ��WE�s19��,P�M`�� ���M��_�!���r�d��ي�֞Gy��3ױhwՈۙ���s'e���1eE;������ua���pq	�;y�'���#":�]�
 V��v^�_pT|5<=�ߠE����Pg�g7w���8@�纠L�z#-Nt�� E끄���s��~h]��p҉�Tɬ"5�����&�J��kE�x�
_�,�42M�Y��?����}�q���82�ͷ<
]����Z�K2�*�1Y�<�h3�f�s�Sl�*ߺ�[����Ҥh�L.���/���
��mp��(��J&����Q�:����C��F)��v��{F�on�� ���k��?��v��V�9�;�0K?��Q��h)��ݎ��j���S.��6�9S�N�-��4�6�5K����x���'	����=��"�ީA5�a�(s�nM�['�s��u|켷�j���3�y"ʓ�,
p�k{�	�Nh�5����ʡazI�8�'�>�^�{7���J,_c��b��ά�ю]�kS:<_�����n�D���lw7���I�"����bh�L4+_��v�"m�m��
���\�3��=�uM�EF�R�������^�*Y�c.C$ bڸ�AJ�U�)�1��ƅ�jb.Oox��M㫞�t�t�NVW5}�MG���ԓQ;͏&$�-�<j.���ͿHH8�1����zw��B%3^���c�t <���Zd������s�,��V���|�t�f��^g�Nx'|L�Zd��4�7y�h�<�Yʕ�y�C�0j���%��*���;�S�e�)���j�-��{�N
@3Ur��z��]a�����A/��N�k\gfex��$�ʴ�&Z-g��@�v��t�'
{����#N���Z�W.�y�F�[N��Z���-�R�N��,b��s/m �y���,��*�T��Vo|����}\�A��:��!�AK�(f�&�t��%<�{��>R�%��o��R��z!�ϩtof�C�N�|�u����e�<�8@� �R@H��)��/�aT7���^�č��/%��,`�p��݁aЬ:�$RHXbOج��wC}
�d�����1P)�=U�:RN���P|_���g���RI�Z�3A�ȓ|W#Ӳg'Ō�;��}B d�!���[�ǣS�G�-V\���2(g`V��vv����T�W��.3���#E��:YU�,�tG�Rה��ӷm��`�| ��٬-���9���i�D �w^��ZU@f�7z\�IA��{�K��m��1�I"����H�J��S`����ђ��[�U����0���}�L��;�A#�O�k�n�{�=z��?�a3�m���&�|��IvL�O�]�)T�u��?��=������FX����?髦�~�F�m��ٕ
c�7kP��Y�m�V,��>�r���o��x�|t�!����1�v(������@�
5W8�)ckOuW�ǹ1ϠO��y�]����.�~������;�wG���\:h/j�y�|�����{pՠ���L��c3�;�K|5�12�N]_ge����8�������{�����a�8�}oU7�'�h�P�ؽ�=6����	�Pn>�+�^ͬ�'�r;j;�v�.b�o�$8�f��<�@�.�������p���q�fť�<tJ_��j���q�v�yݱPlS�1fE�x{��������e����s��p�~�_5K`2�0�&��v�����dEuX\�⧬�	]֛�O��(,L��J%Jbۉ1SYɭ�ۧZ�<��$C��
���9�#��Ӗ�g���g�	s~�,�����c����:5V�;`�s15���h�/E�t�����
����ő��+�L�=}.n`�~QW{]npv�xC�X`���e���9�R6z}�	}G6s�i^�A��CѮ�"(7��i�	.c�h�a����*���Lh`;�DZ �
DN�0�A}���H�\88z���xR]s�o�y�)�=���j�=���p5�����u��)!a;��9��
;}����h��:���4�r��_o� ���V*�bpW|^o*3���p$t��1���t2S�
w$S�HG��G��s�x��lƘL��ɎW�+�9�=��-C�>,k���Ilw�i>�+nQ��8&����J��~t�nH����&֜|0�7%G���N�ϯ�fy����L/T�VI,�Nrl+xR�q���n_a.��h���}�$6n��Q>�K��3E��v�=(`��})�ft���>P�%�0u���ޖbd&a:�+Oc��i�Л��ژ��������N��ϡ�A��
`%dl��ZM?M;Գ�Ą��[����Ff�<zD;�fO��W�@&2ǘ�Q�9���-@ћ�
�"�G��n%�Ӽ���D������ؒ΃��fp�/.O���Q��O�C��_�h���ז}4�k���i��~@pp��{���%)��謁h��+D���O�-����<.h MAU�v�Ņ�.lQ�^�`�y� lj�_,-O�Y&nX�'�֟��8��L6�6�@��[��b�Z�Ԃ~G^�%����ұ��۸�]~2���^R=!���u.��I�3��v�k�Pu	�({�<h��!o�D�n���,��KgoSY�k�kO��j��<
[iX��EwC�~	���Nƿ�I�Gl���W��jh�hqWdkp����� �{�C��H0�N�����V%�����
�� ��Z�M"�k���Z�?�_���3Zq_l4�N���
�Bz�Q��)A��f_@���4j.�?UkD�[�����䥟Жi<��l��-�<�Ph*����x���>Y���Ȑ�3nh�>.���$�+��5_'O;2,�S�:a��<h�$��H��@�2=��^�0�s��у�H/衢$�%��"ް����]&N�M9����Y+`��0����ҷ� �-�ɒCo>"��.����g'@�FXv�:
�c"6�L:	�@���;u��E�j��V"M�rM��"��v@p�*�:�R��ʧK�,k����hg#��Ŵ�X���-�~p�B��U�5�#��TR��0�e��/ρ���l(��wy�����04��t�+uy�ŏ��`��4ᴌ�$؆؅�5��O����Ȉ�-�z�ܙ��پ
}Ѭ��L�|"�sE1��bu�|���^�Z�w��+���ℿ�����ɉ)��|j�;���x9�B�,k�t͘�qBlM"���v��Ž|I��֛�^T��[���@�,���n}I����ҕ�%|�� M�+(���{j��Ȏ��Ɍ9�����Jd�s�ɐ �&�/�����j8�Xu/��d��>}{�te),��Z��B͟ �}�)X����v��O˽"��c��) ��N���g3�������ub�C��d�6Mx2'�Җ5W�\��8�N�-XϣEw�m!8p�rDM">�$��lg\1�y���=��M��0�yN�����2�C����[�so�g���!��?�;A1)����{�9f)�Y�����:A�����B g�FB,ئ���h�|hH�&oFCp��w`AeZ�ف,ȯ=�<��gD�텸g|��RW�e������&I�^Dx/�d���A�n+�=����2|K����G�N�o�|0J4f�a[n�A`sɁ�Յm��^-�䅒�B@�E���$I����J�|r��id�!3�b`�	�| �E4w�[���l@��v&�9k�AB�E��VįЄ*Y�Y��S�&V^��z��%#��"��,��&�&����ͱl�����RD�f�?�i��z�Ҥ�+ �B{���Cv�]��A�+,qe��h��z��b)3������i��`{2	O�y*v|�bgEU3U��8��!8,��!�	�7��y*��E��`��IW�?6����,���m��{����^��H�N:���Duæ��:G�J�S�K�7�jc��f�+���� Z��v���?'��\���=1�XĆ��a�?��T�3��t��T��3��9w���� ���´3:ln����ur�9R�N�-[A=��Σ��-��}���"a�0?ؙ��cjsW3[ŗ������s��'++�!���G��~�fcO��Щ��5����L^NX2�oM��t�ZH(��qN4V>��R����UUXOA�U�>3�����k�(Vj?�������DA=?>|<;�ɵ'�9�����r5Ɔ���\4bQ!�˗��p�&5�@�i�ut�Q�D���"]έ�K�����"+xZCO���R���1��e�G��D�(�+���4��*UzW�kL��K�y��	)u��u) �M��)(e�:���[ �zk����H\���X��L,L�h⫈G�,i>Rf'+y�A��Z����%��Pxp��/V��|��Ӣ'@Y��`Q��L*�2��_R{*3�ђV=Q�M#�l}�+[�_<��5`�oꗏ�܇�[m.�a͊fl�g͕���:�.��@;��/�����?�V�`,���/-ŗ�'!-U 9a����3��U�������%��ȉ��/;�9�C�v����#�c�J̹z�yc��b1
�~v�����)x2��\X����%-_m�)�=	n�V�O�m��5ai�f��)�E���L���gk��8��s�M���E�_*OЃ��s�TA�k7CH�O_����p �ve���������ٱœ�����|����hlD#*����_ �
٫�
�?�����4-^���*��.���Qҵ��An�@c?���4�8�e.�b�"�/��3�����go7x˶sž��Tv�-VL�*\V�'w{`��9@��8M;�C�|�M���� �����!������}�{��My�x�)���p&f���rb+��}��v�] S_�.e��lqF��BmV[SV����ڨ8��Jc�F�%�IP��t?N���4(-�F9g!�%��`��d60B��vs`����^H��)c�K[,~���Y�^,T[�|�כ��`��6L� �1 (��c2��6�׻���}����<��%2�(9rq�/Zu�j�-���n������uU#�~,�������:v|�p��ov�~#� �r@����V��V���0��&���\�E�D���	-5t��=ly�[�U^~��ȧ''�#䥜;��YK)o�>V�b!�*ye6p���U�wW>�TE�cy�D�0��Ek._G����YA˻���[m���;	%��G���sTp0ր���*�V�E�VVu�τ�_@���b[�ɪ�ÙQ���嵫�ˎc]snkw�8�k�����|xs�ŰҦ?��I�7�q���_��g�˶.���Ss�S{�}¨n�	���]FR��ݖaA�1�11���J��+�*0�^���3�]�z�ȂB�ߚjM	.���Z���<~Ў���ʬ>�xV��j��	��:3Z�&o��8}w�5'I�c���	$�=?ꮞ��}���֊��o�k�a��-��QGMmO�gʹ�"�ܸ����*��jLOh`K�>X򖋬���wԊ|U�ssz�O�:�b��)�;tT�6~[U��Mcl�"3Y��9���%�	��9@���� ���G�q�O���=��Q�eH�O�jv�d�+�5����8�pd��M��i%H�`�[��.z��^isi��̗�� ��޾�ܩWJ���)��]P��H���b��ֿ'�Io��2�Ņ�,�
��O:B�6�U&������
!�<^Ӽ����[32bG~�I�Uĝ�Un��7�=A8e�Ĕ�<�|�_ȵ	
�X�T�'�p��.��Q?�O�g�Q��38�NP��>��&\i�m��
���Y�b�Z�0c.�>��NN�����)j@)�_�	�#�!�L�x������G�c(�	}oei��k�p��q�"5����6w��`�Ñ�Eբ'��"��-���N��J|�:AT�R�����c���]�*'17�B���n���f�>j?t8�T��yS7���L}���G#�M�NGșv�����o��-���k���lk.ђ���\)P�/��5���!�/�H[�d�����7IwN@"�kr���,!�в��;sB�J(���V�C9�P��؂Cl���1f�8���3<�ǃ�	)1E�:���s�)�_�%zf1El�A�����2��w�ѓ�@<r�خAyˍ�a�-8�󣡆����h,7p[�W3,q�8F�Nz;舮{�>��~6�j��E[��R�}������_J&E��uo���6>�*Q*�?��#���k�]M�I���+�߾T����:���,����;Aԙ28Ѧ!>DP+Y����0#��v=r/����_k�����n5?�x���=DF�����]}y/+�t�I���K��]���X�^"�L���n����9�oO��Ɨu�_�#gs_G=�y��f[mhl�Y
�aM,���<)�z���)GV���\��������ɾ��gp^bi�Xv�%��)� a�>ώ�����E��Ò�u$xL6e�C���UWD��]��6�V$����+�'x�?}�"�i5�p�+�?�v�v�j�kE�冪��������Ʋ�Um.V��Ĝ3����`���aw����$x�
3���|�XO�t��M��h��rb�~����E��	%��5�(�6�B8�E�R$���-�JqƁ�ւ��*�y/B%?�(K�s�V��99"/��a��M5���`�Qs�ķ�