��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t��"�>m���w-\�A��@Mp���Gq�1��HQy��:�/W�0f,1A�2��Djج�mW�$!xzWG�pc�$���;�%��!:ۮ���4��M���}~>���?�g� ���G�cEi9�W���H���H����P�#Ei�G�O����JV�?,��\��X1�D���J!�����Lz���%%'�;��Dl �	��E���W���C��-��3@�������EV@)��t�f��z_��V'�X���#�	A��tcB]�=��m��"ϴ~f|S��.�q�"�٫
�߂ݒ=�әR�bà)m[�	��`�Z��m3w�"����'9E�gB'w�}oWzHڛͯ%~��6�_ޣ�RT����)4o`������jw����Iq���r�~l_�fz�?����.)F�^ǡ|G�@J�[}!�2"�u|�a��j��t�贾������/hnC�Ԃ�>h��Wɱ <q����-k�s��kl���#�����6Lm�Xko+���M��Xx�<�6�"(G~<z�q��z[3��+��>��?<n�' <�c����`'ֿ8��m���2���Z����`_�z8��G'��NÛ�1�y���n�ڪR)���9�>T��ؔ�Œ�����cҔ�1>i~�mD�	s~�X8|���t���
c$�� xH}cװK�(�G;�Jv�X"?���xs���)��tg_�9�(B1{�������|��=��h%FŊj�r��۹1��M:�v�e�y#�j�p�Ry��-���m���vI�ΤW��c%����A�J@���+��5�2Z�j�#�~E\a���dm�_���Q������3E���!�pI9S����a�z^W.�q��Q�㩟Ŵq��8��~<����+piS�P��!�"������*�*�e���E�m��/>�o֞���r�b���:o���i��'��ؠ�kxN%�!-5&�6�eD� ����&��"�v�����)�U ��^�(h�6�c�'��G��R��2�O/>dC�
�Y��(T�@�-�`7r_�2%��>���NMZ�nZ)Mh���U�����n���C͖���!����2���V��Jiv�9ׯ�!���$w��ܬ@� ��m��]�o�Ư�R���V���`Q[|M�0��6y��̈��U$�h��x!22�u��E!��1�	Bq�Ү�:�f�(F�L^�f5J��IOC%��w�Mo¾�a�*�=CIþSeq*5��`���^�C�2^9��a4�Y�%���\��i�Ȁ���Ĉ�"::�S��F�� �X� O/�Ec��3
��oV�6T�0v��B�mцh,�%��4�OĽ�s/�n3�?B
�aV$%ݸ��ڤ�r��Zx���n;+;�Rg���q��HHx����9�z�?�H>q�Aw��#F�y�n���r`�P�u�d��TmU0>�Ϛ�[�xi�T9�n��Ц0�t1�~�:��e�!*��W�K����xdZY����^ɟ�s����FǦ����RW�$�ft��or��/s��G֪�tĽ�E��k�\T�½��u?6`��>���@����*�>�m���,�Lݗs�x�da�4詾zV"�xS&H��-2��cKU���7���3� x|��ѵE�?��-��@�/$�O�*��y(27���|�@����]�XD4�3��w֓3ij��YW�F�������/�<7�>-��(~!�%�@�b"���/f:g���B�q��j@�n��-�z��b<qD�XsS�G �B�%$�jj$#s��U��_��D��<���$�2�"�KE��l�%u��m��g�Ec@�>'(5Dg9Vˏ�� �#"����T�𹚸�4#c�%E�^�.� ���v:}ʜ�
 ��͔6��B��2H�d�{v��l	��'5�>'=E	������%�!��&�e_�4�2_$+m�v��FX������w[ڪw��_�X4Q�D?�K�j1��1<0�U�
ʰ�lK]�$摽��L�9�1�Μn���E��zL��Ƞ�Tf�;��ʻFBǲ��n�����w�C:^�[�1D�j�Z(7�(j�)���jz��h7�}!�2����ꥉ��C�"�-��a�ۚ��SV�����-1^"SP+V���X�Z �B��?d? �f��=��T*���7������r�L�D�1��l+��QxRNd�T��l�Q�&qDޑ_��(m�40�$M�Ѷ�Vķ},!<:Ƈ��
d�Q��[��dN�����ʍwkv���z��	�9q��?m�T#�g�H�EV����``�K}1�I��U� bbkY~M1�bY6�K���Ƙ�2B U�{*�;��#aC�)[�����[
ӻ|��[!~+�@��6C3��Ứz)�B(YS S|�Z��*�v3�0O�	}\�1x�&L��`�;u0��lط]�0��x�Q0���k����G��V���['�H��Ȕ�:˯o������p�;�6�]I���'	Q�GtD�<�尣��i�ő��>�x�I� cȚ[\�WM���jKި��<7���^d��f{�G03:O�s�y��ٟN>�p{?�+H�濫�U�
��,�=�y$��tW��J�"^���6$��f;g����0�=����_��j�S�1�ep:��T��X�$��4p�;L �}�!8'!�~��kT�ƙiw��6(�R��Q��ց{)k�#Q�pn�Rvɂa�R�>�v�S�#)%Q���#�̈́�cy�RC����U4w�X3�g�a�B�s�q�/v6<�\�]B|�m߼�Bc�?��U��o����B^S)�0��m�<�ό�a���,��z_�v8Њ~6���=ʹ݉�c����h7LKהY0 ����1�b8��� �U�S�l�-u��Q��α�y�2TpK2�W�O���݆?@�a��s];���j^t��(�F�����Z���(�\xz���-<�_���)X�D���� �jy�V�wIy�P�IΨ.�`�	:=1!����!��=�{�߈��P��1K��E9�dw5���q�B�妱{),��J�و�0�� �Z��	?�������S]>�t D��'�(\}đ�{IN�X��@��z�.&m߫J�0d_���t�/�������Ǿ�����h�6�k�?=1)�q�^�� ��P��ٱK@�#�RLi�2>5�):�ZJy듈T*t��k_��#��U��й�PN�6���G��'��ϙaI��k�aW��9�p��͟6���)ٹF��k^� $�8}}�p�kg!�����nx)e����׮:&#3��D��N�΁�Ğ&z7ϰyž��0ގ[�s6�C�|W�D�%7fڕ%������a}�V�Q�3%��D�� ����]������9�O�D����_���[�ؑ_�V�﫲 T�l��i�f��N�S�D:�ndO�R��TNJCcJ�II-�\���,�ux�U��A���rF�m1D58�E��x���UB�O�����:Ύo� N���:�l������{�_�}!@�]�mx��jߣT�!��Z���8 �v���K�?O|�e=2��5�OoI;OM��cM̆/�	�}n�"ȾJ��::�TAn2Ij��
�E,�����K�fff����5�G�*ۋ���a;#����e�`���Udۤ����?�Q��`?�~��7x:����ڦ [�ch�`���P}�)}y�cs��	��R�+v�x�*PUح6L�Y�{��^!"��
�NA0�!�'Zm�/DF�^��>��g�&7��]����N�%���" nY�M𾖶���/Ek��:����C+���KY`�{�8�����$�/�����1��M4�M=�%���aܾZjX�[��M�+�M�(6` ���o^r�����\���m��;�2ޮ�m�h�m��@cX���q���"���^�r�/'�]j��D+��b�+�$ܻM|�]͘�Q���,d|�N��oD(�DFU>�{vd^�����nXt�|P
s�b�GD�<d�9k�{��eIH]6��4!�O�M�^c[�i�i�o��J[���/��Ι|7�a,i�L����XTH��l���o�iC��)�`��O�t1s���J�Ї�N��N[��H�i�o=�2�FF�	��.�L)�}�I�F�Y��3٨& ��n�|��/��"u�6�>�	�	GcvYB�3��%���=�ԱY�
��哎���"�;��RR;���tr�F�(�ً��E�5y��\R�Z/o��Q?�!�9�)3b�F�>�|���[PG���`�����1Eg�_�u�U����R����T�	��%uk��R�ϑ q�1����c�QB�J%}�#ɐ�D��<`fM�����HY�9���@Q�Mk/S�o�������L8V�Q y*��U��sifh��N��c�U��"���i�߂���Dc�ˢ�hQu�|^�O
{FK=�A$�Sv5+~dɽ%i�OJ���j�-�LT���cR��NS�6�tV����xg�S�]���>E�#{-�����#T��T��N��3��u�]�G�y{|6G�K��\���"�`�zi�6[9��{���3�Oe=�����V���4}�2�����I2�Ջ��f���5Gyણ[NC9�����y��?�V���˄l��sz�DX3���MH`��Uz�qܥ-���(�F�>"֍��m���ב0�e�J�9����Q�`%�GF��^ϻJ�`r����H��§Mh�^��o��zi:'/0����^C�r�����y��E�vﾍ��B���Qt��ЃQ��L�@F��~�}����#�G���G�L)��׹�+.��T�?��;��e;�sR��օ�\M�_�U��Þ2�1g���JԤ��bul�E��8�{T��p!a�e��kF/k��Ч�?z���7� ���]Q�v9m�?�I��Sp���n�X,�d��MH���b��vT��d������BBRE���Q������!�/�$q�z��D�H`���_��$Fw���;l�i,����K9���&�$t~�Q	ׄ�;e�Gn)��L��Ij�r��Ѽ��P��kf���z�I����5�B�j��V�����w��5�����u����N�97 /*�8wᐏ���^����~���e2�S�����[���h�D��ӑD���k����b~��ȯS$6��������)���
�e$�1��x���Y0�h���7�G��9�'�C��
�(���*P#<��$�"�է[W�=�0tdB����3�q�͗�����v�y�Y��}
i�Bs�`a:��{��G�Y����zϖʎۂ媂�~�n�}'���U���l(.,�(g��S_P�E��螟1���\ Z�t7*Q��G�!j�Û�|eW���N��Y;�'�iZ�&�E)�����8{ũ�%R�����.��.�O}�`_�0��6}} X�H��a�Z�)�W�HF�zf�*���]�����ɽ��(�����k���j ӑ�W��(�)�b���#`�?��տg�Q�z�bb�����B�='?�n
h�_�t(-;۔kH��k̾<Uη����c����02��W�!�q=rq�*�P~`��۪n�>�h[������'C��y��>�4�ƅ�٫��#�;kѕ6��V��x�y��m���)}������Up�&Tk�ΒV����)��5����Ҿ��u\��ǎ��A���y:`Q���@�Vܼ=3�0���]ÌSF �f����` ��J��r����q���ֻ�)g
jPp�ޥi��|�����;�*[
��� �D��p:}I�.�-�psUQ�ǣ��g�����"w��4^�����0F<�W)���Wލ*����p��
Q�MqU���*���DrA��s�R���f˩�ZF�����a�y��Eٰ��P0�p��1-�tEkShnҙ��A��G�֏zf���p������W����.�0��b��	�UM,H�8��D�Ć;ԗ�]��ڽ(l铃$���C{�5��k�'&IxA%=�HЍjZ��?�Ir����]�d�}Տ|�?�:��6����E����O�F� �0x�y���%����M���ݜ�g�׺�tbĕ��v$_��Z	t�a�0�K�4]�Y�ɖ�c��'��9�Q�!2�h�qO (�����v_.f��i �T��"�xe� �
����l>���j��-ս�d��x�k=<N�}�����/���d���ɸ0�I�ʞ�#4�A���XL5]�@4�0"��ZL���&>���X���u��]?��h*��4��f%��i�,� V��B���|�J��3}U�R7�F��w}����,&(p
�J��\W�p�}�Q��g�G��/��b'�-��c-��sYڡ%�ed�Tt,Z�k�e�(���vg���G7.�bF5�x����,쓉rX"��%YY�a��ꪌ^%n�a�<~����Gɻ�S|E��8~-XC{ n~{^{S���p:�k���6�O���_��:�����`�$k'��{k���h���z�������]�<�O��1P,�?I|^�+p��d��ޮ&��d�k��}�E�v�l�Y�|�ʇ����X�Xq���	s#2�)
	�[L �1t1�(o��hzLNe'�st�K�MrPq�Կ:I G0~i���,uԙ/�2�ϓ���\E��`�7���D?1�};X���(y@T>!�jQ��[�Tt��Rq�����HP��&��D�ML�X��W���2���ψ��f%����a@��=*2��=�Îa��(��J�e>�88�x�o��<�N��T.Ohr�@���C��*�����a�V�#�uB�;��������[��͏��'�4F�b��}װY��q��7���7�*���p��0�#����	�R�(�Q��Z��?���$���gn��p�Uα��g���/E��B����\o���w��d�0#t�����_#5f�\,'�@<d����%3D)�5�)�͐ 佝uc8��{R0��q@����Re-�#��P��,,{��w��DI7�>B�sx���:��H�[���]�<�v����������&������T&5g�6��0r�D鮦�́X�L*�Jݗ�-�B-���|L���+(31���ƈL�6�Bʽzl��#�u�L�aͲ�p�n����?"Wݚ5�^�c���+��dy�����VX�p�e��=i�{?��9�[�yO�	�/�
��EP�k���6��v)����]5��ڌ��*̍�y�/���� �e�8��<��H�nLA~0�v0ee7�'�{����9���Ӱe�1bX	B�����;sϵ��jw��xZ�e�.J��6d�1�
���KD� qau�M��`��C]O��T��3��̡�IAų�0��X���$8�nX���|����y����/,еb��~�>�pc�i���~�%�`�j�2	ODO���g���P3��\9��=�,QZ�[v� �cX<������7���I��΁��e�M�������3�k��J=ScA�,�t�H��ct�.�נ0'��<�c�^�K
�xn�;��w�nzR����l7ihɀq��l��D�+	��O��J�hː�;L�v��{b|h�;�Qz�T߱�����27\/����F��Չ0!M�Ib�p��$�;�/�hf�x<����Ç�J���G� n�m�
c�J���5Ng]�_ss$��Nh�f+$�wľUI��-��'�G0!p�i)э�=M:E�B�������H�U����qB�=Z;����$���}�5bX���?��:W��J���bX�0��� F�k������8)t�7퇲��S'�o�}u��Y8�G����n�Vu8��rX��Ij��էV=5d�0G'm�=Yz��S��j)�S~6:�f�@эh~rL��XR$�E��A�غiu��;�^goٻ�G� ��H���yϏp�0�a�8a�G�=tmc����B��V�N� �e�i�g�����<\�_����A��r�N*l��[ߦpajiN-���Q`�k����Z������*�%>���Da��w���Ge���S����D���,����D�?��`�1C:w.��Drn՗��P^B���Se�M?�/���F|� �v,Fp`��-��l�9s�p[=��dm:5���^{`�c��k�k��K[)؈�Zs��Å�k�+�ru�+`1	��M(��m����Cg����Ƥ�x
�bT��<U2�>���}l��H+	&\:���񐷆jlƿha?����R=�^�$��??餓��F]��(��G�qV�����M?��8�� �҇c6J�Q�Jf	�>�8	F�X�#��w���*!���G����-��0�@��vn���O{���D%E@:�\�`�zeW��5%�zmz�+��l�(x�%p��9��rzcriw�� �و��.Sq�����V%��h����V�cg)9�+���Z^���&����?"ڲ����0�Y�1�\3
�*L&� �p����՘ #`�8��Q����)�=�C<$���u��hd�G�z�p���rep��w)��'�T%�gR͝�q/��#�	��c��
��r��A�jaDc�Oª�ֵ��J<T]��j_s�!�X�������Z��`�ے��X�T5=͌�h-�����Z������l�а��6@ �^��G�shr�����>���Ͼ������[s[����O}�)���1 �L��(C���)̌�pp���(m�y����Kz��DX#mi[�%ߔ�Y��{f���q����s�H�d��M?���O��zV"�7#;kO��qXf čV��0?4�_��4R����G!���ӷA3�$r���b!ɒ���׹�0üx^e{�	���sU��t&��Q�ǵƕy��s�_H�ώ��P�	���]��<ɖ���(d�.Ž��~�t0͌]�5d��M�3@����p�5!A(+qJk��S6O�2��A">���O\���D}�2���d`��H�L=���s��'U>#�G����-d�U��x��t�#�7f��.zH����{�sh{O�A��q�5{�Ċ-�(P{]�����۞��+�ά���k�?��Z1����H(�T\�!R������'��g���]��n&)��2��T�#��ّ�������B��',�� ��1柎_R��g�B��ė �>)��	c�,��iԪ� �!��M��DcG��0��>���O�/ߴ��۫�zbM���Ϙ�bA��!4Q]�h�N�ġ�ɖ�sV�x��%����N�W���	�2��>���|�I�x�%:��[!ŏ��ŝ[�iҎK��J\��SJ�/�<��p�W��]	��G]-���iM��Y�)�2,�c� .dX��e�'��8��5�ir���}"��L?R	؇��1�Q�;��l�8��@��
hV�b�;�E�_^��ds4�׮�=��%������o �U�Pu������Â:lIY����t=p=!{��ظ�Նs�����~�)�L���b?��0�gc+qp-���~�0�j������Q<�ƴ|/�<Q���fylR���7	�
������plBEC��td��羌�
��{ip��!��T�r���ϨU0n�	H��b�^Q\H�7��,�`�,o�j`r��^%0݀ 3�ڀ��f2>���Ϗ(��h�̴�Q4��f���㔣{SI��8�x[���b�QU�Wr.��lo"�9�А�m�Ji6�荭�~_t%�<j8�E��H���9�R�g�-���������2/�������2G��t6���:Z����Aݳ��B�Pw���_�}o�Lͦ�d=�ct������9�k��U��fl�|�����y�r����	`��7�1
�Udz�kyT�pX�*f6�sb0F�9-ъ�{Y{��3��qx�=��<�SP���n|�7p����ι�-~fd>��[����ۈ�rW�@��k�7Es��<x$��e9;���R��)��pF��-�u���p�k��/��~3�3Em�
�����'��鹴�Rivn�gy�섳6]�ɠ�i��e�ةG����oxS�����)j,��F��qe.�LϢ���7����<�v����#yo���[(�)lWW��Q�9
��3����$�'�}(�d|�b�Oz]"V'A3� P&U��aZ�8�ڀ�mJRj����`JS�s+�{<ʠ|�_�W����;�k"�4��D0k��(�`�˩rK�~W����OGeW*`�\!4��Y �p�����^ߠ��oݮ�qs��ď0�P˃׶�3�p�=�'�%+��z��C��p��_Z�FY�?��T���H覛)>C�]�}����/���� �S,�4Ok�k�=�
w�]��J����s^Ċ-��o����B��#v&Ϯ�r.�UW �cv�� TR��&&��U���eg$lɌ�YE	��#ay�ae�QI��EvѦ��s3��y�x<�)�G�D� �-O`PU@��A�h�͈��T��_�kIފ�91�/3����)g�����h��5ȜŞ@U�:�y[z���#���C>N��)v��J��lp�N��Q$M�1.�^9��#���N@��:J�/3����Y�o	R��������3"\��L6tׄLD�̙\�+��y�u��# %��%=#>m��:qvY�ǎ1�0�]�-}�yW.�r��BqF/0m�������8P��	�?��
�Ъ	OW�~E�Հ��1j���Sq_�2��k�=���Pڋ�$
Jz��E���j�0G��x��n�p(z���6�Y�)�3�Z&x� ��(n�=���G0J�����cDB�o6^�y�+���K���L��[b��to��H,:���qwA:�@�];�݆�'>���c��0/:/\g�Ӊ	q��=|Y����?��a�7f$�C�o
jf����i1w���������3:����x�?D"�6꟥ץd����o���{�'H����*-9��A
���[�;�訔.{�2WL]��l�%�0}w���f������]mߝ�����;�l�T�*P�{��2L]�Q� ���5v�|`���eH�3�TzM'�L/�?*Ĥ� 1��9m;]?����q��:�e�i��x�.f������[��x{dr71�ca���l�����z���Q�Ow&GV:�O��į
{��u׿��5��:��=tXLPI��2hH%�ex�b1L��Ȫ�dk���x��R�@�J�ޣ��+x��L�y��\���|x�Gh�q��	�g�p{�9�߿�Ce�E߱�-@��/ [��º��#Ŷ�+�#���en�@ٖ��N0�{�*z�N�@\��gJjs�a6�9�s���G�����C��c�XB�(In:��.(:  �C�k��$�m�\� �Gd�39xT ]Z*�_�J����M��ƫ?�����1�]���~�E���˥}����UxW�����h�&u]}����`7����q���c?�fP#]X��h17eD3��=~%V��桰3�%��p�0Ƽ��g/k<��8ߌ �ˡ�4�0��|�Љׂ�n ��Hev�CK���+��Pb^���7��<嘆���~S�[�mx�������w5���K I��M��K�p{�(.���z䳷�m֊y'��5oވ�V�n�Qp���IT��Ɠ��v߲�m?ԭ��v�����]l�t����_�-�{�Js��
�v$3Y�ؗ:l��ɢ����>a=�3��e�'C�av��]�
����ɿ;�ڋ�� �������N�u���	A�h�t`���'&�'��F-Gy�h�׎�m���:���jA��wH��Ŷ�������4ּH�)�̔$��nĘ��cB,��Z=u���1��n����Y��86�Ӳ�N�S��������]�@b�
�*y����/<��@�+����;-XA_�������$������Kb�p�P������T_����-��E)���­�z��\�F�4�� ��L_F��.R�O	��|-�R��ĝ�
0#I��*t�`�o�E��y�I@�HR�Ŏ�y��z��|�.)��g�o��Q�9����=�Qfr�2%��¸��YZ�b�d(8��NH���N�������Tl	�ʑ�ֶh	/��0�"����"�'�+gR���,G��z�fc�pX�^G[�oR�4�8����B��6M��dB��������p�C�w.�	l�&�F}���U���=M��8�'�׻yc,i����>�obhT >c��5�x�
��J�4w��jW`�r���M�\���ѝ�G��:�!����P'��Il�@L].(����z���W~{)m���wI�Y��.�A�G" Df��	Y������2ZRn�3�&fǢ4�P��}�gW>�JA,6��[���_��o���Qt)UA�e�ƨ�z�e<<���0�$�)o8�
� ��P�@�)v��R�Ȅ1�DHg*PX	,��2��|���3�#�l�IK`�G��v&d���M^��w4hڂ٣�.$��#vV;$��U�q�Ā�N@��f�P�9Db�-ND�kF���ϜJ+� �;=}�	3~�飳� �7	��*׵�l�����]��ۋ"/K�C�2�!��殘�v��9DDZ�Z�e���V<��n��xR�b�m�|���z��_a����P◓@� �$�I���D�HR����">��'���2`�.���_Dg����;,��J��r�G�+U[��TI�pb�s���K�z�x��H�ᡕ����)����ݵR�����?����ɕ�aJ��ƣ5P������3����-9�^�z搔�uY�H B�pg�Q�nف��y�|����tQ�F�A�l�頿݄�X�ƾ�;k����ilw����T��P�۳ʎ�Zw�%u��S��h)EXSY��_h*^mMS&4�u��j"z�W;M`uG+�w{#�ُ��F��e�ᄺ��Iq�� )f?�w���!���|��f%���~�M��xZzWO"Q�#~�������B�z�|8�h���#�dW�fN��4����t;;�qߜT��L�Z�brd.�8�Tz;�`n|��U]��Gg9�����N�w��KQ��Ǵ��5�@fmo�Dy�K���עj��!��Ȍ�gv���!�Lk,�M>Е�ΰ�k�I�{��F���ŅSF��P�qu�V�;"q��h�^�4q�I��!��/�A�� ����������TW6|�ɱ4���TQ%���o���k�i�z� ����m��j���M(�Kh\R�JM3������:�n�Y�ٳ�\Y{SWU��ޤ`0pƢ�1n{Cؓqh*k����[�^qzi5�
pL;�-�F-���'v�;�E2�$���Y�j�A�������� O4}Pjӑ��&)9�j� -H�g�4hQ�Z���+��d�;��7z7&�b#�s �QY!�ĥO2�L��a�����	8�-+��g�6{���Y���Z�A�9�Um��'�����(K�T���/���ee�ߟ��� g�|���?��˕��l ��`��.���w�������ы�D��R{��w�%���͸^�+���+�1˧�\�5���m��W�xu�3.Vԉ�?ƌ����8}4�'#1�&�+�/%���(C�q����}�E���e��e0����^�7��d3b���_xZ3O�X�%/V��-j7��m����%WP��d�P�x��D������wΟ�i�U>A�����-��l3����4@��J��_�=#Y0���8��W f3&���.���y��J��I����@Rj�c���3�F���
��
C��������g���;�S�� �,��7n��?�!¹zX��,��h�C��q��pkX�����zg�	S�H\�\�+�P�eC^Wgz��ٮH��tn����M�w$bL�ѹ}�뱣�-���W�uj��hӭ�^Mӭ��M:���#:e��/�F��("#�(~�T���������&�S�.��\t4o|�V�s�{�5٢tX�[��8�!�Ǚ�é�#�kE�4����G�#�A�+�9�l1X���H�f���'OR ;1 �g̖~Za9ݼy���}@�c�y��i�8��}G����wE����D�Tӎ�����+f�i��x4?�W�ø2ũ��'Ш����
!���H�Ii$� �"�@���ZPa�A7!�����#�b�@ݔ/a��&�uQ��0k++K+���J���]+P��v/��*���k�uyղ��1���l�շ���␜.����X��EJ �E����N�>��L��7�p���>��������:�������I�ԋ3~N!�֛S�+���/>��&P��<�I�}�������K�EqY�N8]-��3�c6�ے�X^r`��V�`�@�2>s���3�@]�����N��v�!:*(�hSO�?����R�DY��Hx�j*�A`AV���ԟ�蘱�H�b��҅�G�� �sfևY@�h'A'�a���ؗ�� �Z���\�z�tp�k�b�ڨ�}f�kI�b�к�#v�&N��0��r���˱5�#��^��A:����e����DZ�ũ�R;q5i�N{��x'�y�q�/���&Β�U��w��l�U�q`n�E ,�l��z������������Gs�7|(q����]�"#�Dvw�
)X9����_�輫;�W�jɎW�Ks��#(�#�ħ�j�1�U�r�/|��
�4.Q�`̒a�E�����8k_�g)�����Y/V����~�k�na�����|p�����x-�1�j3�b���@�d���Zִ=�Y3�B���Z�h��O�R-y,ަSǩfg����H���b�b4���o��=}�'j��GDAh_�;C�l_o(Oh������´�b�U���,M�/�~{iw٣R�Y��b�
AǒÐz0���Ś3V~4!�c\�{F��wv�M�O)���J��[�����6V;}��8϶.�s�hͮ",�y�J�}1���/ة^�I7���u>�Ax����(�6V�,�QuJhM��I�C	?���'�j��v����^�S�	��9��'�RjErl2�� �Ls¯'�ITx�4;`���r-#���,�$ԓ��gPf�󫟴�(�D��B:�*�u�-�x8n ?��������&ĩ�~�Х�tL���%�+�\�
�SJ�>�:�lÃl�fz�J�X��R9E�t?�-���n������Ϋڃ˫���7�Wx�[�8���;�q�53��I~���H���˘���M7	�;�VeD}^2��
Ӕ�0nE�����ί�E��ݞ��l� uۨO�+�[��Z��iK���"����,�0����!�N����O.S�fϞ3`��Sض{�j�Z/����BMպ�q�w^��2�S��b�lAJ��]��n���*��R�׃����އS���KJ�%���2�#�&�����`��D�R,Y�JK �K��*޺�Nĭ2�&���Hx�I)2mF{F}^u�Bw<ɡ(	�6�t}^��4"�s�uwdo����5�I<+7�,����Ӽ����L�cL8uzT��X�D�y��k��ߎ�V�<��~��.�܃�@�&Y�_�����5���\K$P������&�FLEP�p.+��S �PZ��������&��}�%_Y��HzW�])錠��x.��t����&k}�7�6~Z�����iHB�(��J�0Z� J]�Wn��	�1�f�����D�4a�SaO�Y��C��fUP˷`��n�_���� �;d/���b�4�����[+�):��x�^�:�}�܌W�9xe��,�h���y��O��ݔ���RI_˷��kW��C�u�#&W�%��%���m��)K�t�w/�2�A%��'����۾у����?�/,�jejĨ����es�}?)e|j�$��B��|�~��L4�Gf%�d����&w<��qf�<�#{7��:f}����#�0Y��ʵ@��_��0���B�96�p/I����ܴ��]�N=�d�<k�#�M����y�I|;C�	:$��k�0890�_��׷��к�PFl�2�["O|����٘5��᫛
֎Ӯ�I�i�Dr�b�e�gu�`�"����څ�(>�Y�4X)�Ɣ���pi��ܒ:��B��%�!Q���"���~Ԃ��FP�6�M2��<7�̃�w���C�9N����� ��bez�%0Z����~��~$d�'�����]a�2�Q�Y99:�\e����H���x�U�ӋW)m� �_Џ�Lof�3cޮ������d�뗄��(�:hK2�7�R�`�dtfQ�S\!� ���: �l��A΍�H0-�a�����ʅ�@�*�E��b��Ff�FL^+�A�����H�?�����v�_nڼ>pk�2�Μ�V!L�;�� �;h��؊����ʯ8c�PC���JQ�S����3M��$$% �3Q��x�0j��#�t��<�������,P���۪���jS�����^|���|��K�1mS,na��+��P� �YP� 1�ij�m�K�9�2�W
��b��{m~�w��A糩V|R{�S�n��{��0����r�����T�+Y=3(��B{�t��d�Z2���̌��i��S�"?ñ�*�E|�$A,w��0<���V|�	�-�H�4�(�]���YaWoi.Q�D��TYա)ڑi��j���M��;Zef?�GeHgxi��{�e|�[�![wU!ޕ��-\�/I�Yi�������2&�ơ�+Hi����}���Z�M�⭢������G��!I�y7+�,�V�@[ڽ[�*�����ݵ;�JX���DK&�p�7"�,ۍ��z�[���Sv�ԫ��ST)�	�1�J��Y�d3EK��J��o~��<��%�~�=:'�ҙ	Rۡ@�>��(t�y �9a�dL����Α#f[Ȇ:�P*��� ����Qn��kc��G�{A
F��Sz�5�a ;UbDp�`3����ǀ|�Ӏ����1Q:�hut��a��ɳ$���k���]�ko�����-~6v�0�3@wu]]O 8�!ux4��喳ss���yj�w4Rd)W��څ @�H���"P� ]�����ZG
բ�|*�/���vL�{0^��j{���0E��͓bc�>9W�ܩ6$4ޔY�6�ё	�ޚ4�^�j}����fyH�\1��r~I�]�
����Hh��]n�`����렭�{xwQ_֧��љ����C2�4؉�tAg�'�Ыr\��]6z^�r�3 z���[��(�@Q��R�^�c�eӶK�M�uOKu%ګ�ĪBv���-t�%e-�sx�[oy�z:|}�4�#�	�����L�a��^B�"P��Y�?J��ǯ�$]�MWw�<7G�<�G|ǻ��ښkN[��lw�L�z��ˈ��������ʻ�e��ŋ�9�p٫y\�ۦ38n"�r{!8��hW&=�d`W�&��9 � �����iꇐ��k.����	I��Ӥ�Z��1�/�jԐ0s,`�k����b��A��)Ϋ��&�q?���Ĳ�"pn�'4ߗ~��!䖀���6]�Ą>д;�����E!�I}�,P%����^-\H�zI�+
��pP+��������ᵊ�i�R�@2Ң}�\���Z��
��X�Tb��O�������)baf��J4�T�	�"��q�T3���z~T�������z�q��K�4qr`�w̧E����ˀ�<��0��U�{�����cf�3���J4��6�p�O���
��nCt�]��F���#b�0�c~�9ca�3/Y94j1�!TA��jr����4i��
�q]V���eI��?]"�t:�T�(���*A'�k��	�1�J�A޼*��u�53��\����W��ޢg��|�2$U�b��������t�s��yB\�
������)*�:�.�Z�>����i8W�x��yYZ>8���2�_��l1�}}�W-$ye3�Wc�"�s,�a���"�sus1hԺ�_k���؈��Ē�O�n΍9�f�P�3[��{K�E	ً��p���#�C�iK�+��`%d|��]��N�i?��iH���	�Zl��c�)���b��RW�~<��������6�-m��(�����[	P�:����ue���w��>H���	�	����Љ\o���؄| �3 UD����͙��\O����H�@�̜:�������t�+��7��H� !�\�q23�����:���:�7���1�����$�q�d�#��������f'r�)mz� �e����7�0^�~)v�
�H�����B��զ.��d^i6�o�����|�8A�rN�T�{V���g����ERi��_�l>�!�?͜|tl�T�Ro���qՂ��P,Hc�~�R��fE;�`5��Ou>ٲb�l�+q�R�䗦\�I��꾳�.�"n�'�GV[y�f�B����R��'��k(ã*�J�k�u��5����4�_�ap������?�-s�ڡ�MCŀ��$9��u�WT"q��Z��3�9*6��L�7�_|���6�����O�ýeu��MJw'�H?�BK���3�쑀^+,�S~w,6��6�	�l���pcW�rJ���4_�7�[�uIƥiL�6s���z� �D?.��X��J��d��+0�L��ߧ�?���EqL٩�B�C�$[ч�6���~O���1�$&!�,k�[�X�D�1�|����r^�|���O��)n�Smp�If�T<1�I�@¹����O��O{h��� jm|6�q�Wc��[�>�4�І���b*^d)��jy�
��l��{_j���4��\aD
4�of��b�>og��W|��巾ã"E�CvU��4��Ը�6C������t(4=ʿЛI��8w���fRW�/F?��NvVڕ��s���<���~�z%$½�Z��(%�_u�&��RP�\��wI��k�d�	W�K󏆦U�΍"����S���LsYjZ���	�����=�귟���cǰ:#Vɯ�ɳVƝm��ٙwƵ��^y���k���AB7.��5��-�J�w"�RL}�%�Lԅ>��i�쿖'�^.N������������l���ݯ�i�n���<�-�K�։��%��=XU:�e���`hg�a~\f>K�Xv9���֥�f�,�A���MjH�R"m+��o
5��|p��$��`َg0(��\�]�^�s�Q���NCe��i�Ь��H�t�F#�hN�k2���k���bluGc�x(g�Ԃ�ANa����b�����?�^c_�#n�OX}p��,ɏi��v���.�$�/�����0O�F�OUE]���7�a.>�f�Ht~NM�\K@�[ �ͼ��K��2��I��j���Kt��60��%�F����-��T�_��sEcu7�I5�m�ċ�Q��p�m<iz���Y<�$�z4*�c�.��Qi��r�GMSh���i�hN�\�v ������{�S*��Ҿ�7 8p5fd ��є�����ÉB�
^ In�����T�.�9�N��t��^U~:����R������c���JImٶ9������l�޴�m��{8(V�;.H�<ز�s���gZ=�����*R��ߺI���y� ���j*�@�Kv?)$
kIV)�>,����y�������0ͤ�۝I������S`x����z�aί�V��}a��B�|��o��z�cܤaӂj�]/Q�!��ئ�<�݀����(�a���Y���]�.z|)I<��EIw=��QҀ'�w�=H%�a�籱+������T	�\}���O6�?L�_�p\@��.��rU2�%���|��r��%����/�R�y�j�������׋c�3�\����;��7�dY��6��Ή��d����H���kz¤��ؽh&�% 4�:aX�� �KII�ɚd>/��
�4?���R��%I�-�Wi��O�7��܍l�t�1ߝ��`�W��cʠb(���M�L"+�����yn��1
[�D1���D�J%��S��/����b�ώd�z?,劮�X���,R�\���M� I���W}�C�ݱG�HW�YБ0^�����5� �Pz���R��z�v�2Z�b����B��Y�<T��x}�{Yf[+ݝ�I�S��j]�8G��)\w�����N��&n�����],�Lrĸ4cmf~�ʶ]Ʀ��
n&���V��x���i�z��zB��ئ� 1=���zP�X�R�U�Հ��Z��4)v�ˉÄ�E�<k���K�N@$O��|�t}Zv�o�0>(4��8�U����K�+0��R��$��m�hs� N��`�݁�A�ځ�Av?l(��5a����fۄ���/w�l_l(@~MZV�g����P�a�P���*�l~��u,S�-����L�u�@,`��8�1�;��
�%�"a����	�U6I�E)�pc�9S���H��2��P5$��!��j�Hj�o�4�����0�����,���p]ֽ�wy&
�r�z*�K4�����=�A��$%"?F"/� 7ZX:�6S�X�)���-�1��;>���J�I��So�v!��s9�Ƒ(0����i ty��f����>�Ư�S�j�؈�V�"$Y,�,�(]����� ��e�;����s�h� ��WT��+���&x��W���� -����_,.��i-�Wl�N�ں�|�@�:q�G�=:��1eS �F?��I�ץ6�<��烘���K#H�񽧙F �
D�B*��7N�	D��yRpE_�A	J�qH�zW�ؤ����D�WzU��q�D
�W�j�o	D�=�C��LT��ꢷM���ɯ�U_����� g�Ex��q6�й勼O�8?l��m�)~<>if���۬$�0��83����;ĀR�� )��*����� ���w�PK� +�iG��`-dF�������D�b��F-YTr¤b_5	��s�[1g)�UFϳ�^(�|w�MP�x�%���#]4o�R��%d&�#���3Q�߁&0��}��O.���S�:��zLL�h��`9+p�άD���`Y8���B�U�g|��tP��V
�����-��#}�8j��;	�_]�Bƾ��$xX�#��9��b���ͬ�ON:v��,T��n�N�+D��пl�c�O��<�[�~��?^�e������%!�)��350�;Vm��'��mu��S�-(g�@f�~w����r7��]�ފ�E�����)"%�k eX��|lz������6

J[_��\��RngI4"�hG�?�F\	�����8���<B�#	+�V�SN,�m�20�:��|Ƚ
L���7�Ĩ�����,�Ԡh��Y-rhf�����|[eK�1��8D׊%�=<�jr���!�߾�F���_�S�*m��������ֹ:B4��>wb��  �BfI�b�j��)����$��A�ʖ&\{m��+�I�c��q?�ͩ�t�V�ga��K����܄�-rd^�je���w-	-ҩʷ��$Z��j��#Kn����, ���x���!���"Am��0:VLu�1�ښ-�^?|�:@�lϐ�j򦩑1%0p� ]�)��4T�b��'&��������Z"w"U�M3z쳢Gu7����=��){=��n��s�O�Uj.�rw$���%|҃^�E�:I�)�k���5�����PRN#��Kc���TA�:K;�7z)5�)|?{V�u� �=G#0�'_Gػ��j�Ov���.���p6�I���X�[����W�q��D,�ܞ�S��S�"i�Fn�K*�HN�Za(���n����s����8��E<G�H�E����˩D��\r�4&M!~�x�B�O!l��A�3��� ��Pz��*EG���Ć��{Zk�C�R(�e����OjX�ܛ�������dnp��������v���a��:�I���&� se0g��K:O.u�j(�q�S�lP�Z��р! �gA3E���X�9n,����+�h��b����0՗���6ڝY�`�h@3�X��˪�x���lŞ�.0H$��)�TcW�r����d�bkb�͑g�\�C[3��]Y@�liح@�0�ra�zX�Rj�-��?�&���@����.�r�^+��fpRk[�s�"=mu~X�e����XD�QR��/TcQ��l*�0?E�E(��$�^�u��(��к�I�K��a�k+l��P�=Զ`J�k�f:@ �&(�jqlP�Ċ�nYOs�e����W_Y�<4�_׳�ؤ�ν�)��m�o��{�waa4�\��c-L^'�mAc"��t�N��pJٔ=���&j:�'O��v�>z$j���1��E��ex�=泟#�K���=���Q�<��Սˏ����b\8�/P�-��q'3�Q��SV5��9�>�C}���|X�QF�����	n7�+lmC��ʼ3L��N+�dZEM��)�{���m�K	�	t�'n�q���
A���PIYy�f�ӹ%�+��>��.&�9J�m�=����	2���5�[���y�~q�6�b&�N��߀.i�Ǚ3(;�J�|hss��\TZ:��J��K:�6���B�ߤ�<��U�K���Nf�����F�Y��D�.�(t�o@��W��j�D� �W�j+~����b�0=%ouy40�Bf��t�g�$��1Q�`sɑ��-T�\P��9�jb�`�q3:��/$q���j����j����0�����]��n�h�&R���'�����
���Ů�	���|�����~@�~�T&�?��H%����6s�˧���|���\�to�R
F0}Apk���R��#�MGO�~#q&5E��]X[�՛U�Uc;���:�%���tu%��G��)�3`3���1��1��v^F�z �/G���լ�1:9Hx��/��*�%�Ηa@�H}��"�ov8�S�Dds�
pN�s ��m���_�L�>4�E?U~ T9�E�A�b����'i�����n\+l�Q�^��������	^�R�рAO�>Y*Ҝa����J�C,����no�`�e3`ڼT@���mH��:}����v�p\�����*��ك���C��jZ`���㙲�ϳ����Fw�B6"�]���0χ�H|���K:seC���)*��E=��d��a7�%����@D]i5'������UZ����*=�QJ����ۄYd!-99��mO��N�����e%wY������Pq�!�?p�񼼛k�&�bԥL�kR�Q+�����Y7U_s�U�)�
[����*��@TD��>�F)}���4�=�8���]��!B��	Z[.��#�{E���9?��;9v&m1A,�uc���Q�=����ܨ.sl����{���u��_�X���rheΎ��ܒK��>��d�9q=r�o�[xX,�O�����t6%(. ��D�Duk��E��2�V͓mp:�pjA�u���e�	|<���F���,��Q\�2�8�76���TGr�ٕ�Cؖ��(�#��2�
c)B����!�*�Fi�D�6��Hr����I9��zp�1B�I�ko���E��ػ#��>�i߲)H��"t�W��Cs��\� @<ؙܓ%V���3�W���|5���/��F
�wEiِ��)(V�0t��v�W�$�$�)N�~�=M����,ɆK �tq�����gr���>��g�ޝ'�r�S7�m�����d/Y�#����������\�����R�ӺmR�{��|Q���W���;���c��C�8����я2\���d�v�a���f�z~b�q�T�֧�Dv����@�� ��hk~�O������F�!ok݄f��fm�Q}���aK�5��V`}��<W<Z8�T[�ڂ�sR�|���ذ��E��(�*�K%�dt��@�ʬ��QP �h��� }�.R�6�����_M�0Ei��[��5��(��^�,#����������=���u1cI8BvD�W$�(e����1Eg�������%
�����6�Z�l�~�����1�|Q�����i�$v/��j��2�>ӫ������G����|�v=�Nʂ�El�z mD$�ȼ���-�@E��G�l����;ve�-8�K+�G��A��7��ey��l)rWWM2�������>����:���6:+�3@���Y�Au/��}:�j�)&�З�O"sERzd��A�geSm�I'=8��FS|���$|(E�͠M5+�P1��p�P[��S��G��.�ՙ6�!q* K�t]����n��=S�7��m&�?x�����G)��X������3�@4JP���dpN�{���Mp=�L������h�q���]hk�yp�-�D����BL�{�n��`��ę圑Rw��Z�3�z;�D2oL�#}�Z_�hs���ǽ��c����E����B0ؓ��X�b�����'*ű`L.����/P����$����r�{�}����.�$�tÞ|Y�g�f<���@*����H����ؤ�Q*1�W��H-<-5���<rz@���\�4ڻ�:݃���x�MB�k/��f���7�J�td��q9\a,��%���#���eZ<��U]���d��F���+�W IԒ��?��V�SA�4����r]l�b�gHH�oo��n�T]y��b��3	a�/5n_|�h[�ۤ�"6IMґ�%��4>�U��G^'Ť��nQd|�R�$�/�2������[xd�U��
~�h�#��J�vNS���`INuv�?�b��IE�ȃ���D�x�Ȅ������HpUR4KMpa��%T���gV��w�lIP۩˕�����d��϶8p������U��6�ݻ�������j������0��l�;��,x���T�e!���On*Y>���e4OM~�u�V�'/����s�R��\�_��S�H�ӡ�aJ��%�<1S�>�S�Ե���%D���������}��b|� qܷ�;)�@�_����z��m�����������jT��R��\9ܹ����ކ��r��4?�`#��oأ�z��ΐ�wv�[�����cě1����# 
T�������ܘ��g��H��� ,��h���$J󩸈����Kǟ8H2��� Szx[_-b��>Ӄ� � ���b������u{T�(�����6������*@�G��|;�P3^��I*���N
�a�����@��uF����Ā��4>zH��od�e�a����O6�x��"g��2�r(�I2
W@]�	���k�;��A{,�����g�D�u��!l�aĖ��Bָp����>{^�bߪ��4h��,ذ�#�����S�QQllL�_2�343_�je�(���!���W��=�.��/W��U �_$�kA8"AV���1��`�ϱ�}_t78�*P�^b�ƙy�������q���/����A�ޖ��#;z�dЕ�tmI���(�5Z�NX1���χe��>��R�P�a�ĥ��oN�C�k�?0���o��Od.�3���~���Mǹ?%b��a!w̡�U�*���n_����[Dʀ�	h�~T���W�z*^d���:��G�B��O�d�[�[Dc�3����u���T�9B�9)�,sԩO�ۅ�`�L�}�S|��	U�y$��~��H��N���	�}��*����r�RR��	��Sl�B��˶���zH�6.� �M��U�8)Ģ���\6M����U��>bv_'�b����M��}�^@��l����c�_㦔�,X��]�4{�Y��hR�K���=�X�S��~l���Tӿ�sL���g�<M)H��Pb������@@�J�ኜsY���<�Ҽ&�{�.D���;R���z��,֐#j� �/���J`���I�z����)Q~J|�!pi��"���Q1��2	�ш���i�\���6ug!0c�Z#:������uYb���|� ��R�wT�}p珴	��0�g��Iz������C�!!0xE�vO������	p�tc �Zȸ효L9%� ��ۢ*�ўAn����~��i��b\*�ag� ���L����eZ�(x|��9��$�|~�u��@��ku���C
����X�C՘��,[Q;I���x�l�^�QY5Ȩ ��P#��]ȭ���K)$f��4�?`�vۉX�,���w��H#h �7�
)�$�Y�8���EJ��\���K�!����R�2{�"���	�1���B�6�Ŵ+T	�V������!�LBG2ĥnE��u�A���;B�i֔.y &�,@w9���!bȤ]|�Pʡp� ���<�f�e?���1l��|#r�����`�KR�y�@Ϝ��9�Y�c�p��m7ߡx�09ݣ���g+��+\4�^��l.����tOO�"�G>p�*�]�9�RC��'t�� Y�ȶM	�E$a�_1��6%�PR�?��G5�M��[%�/��y=�ą��j�D��5O$k��Y:���%!��:�<]�r���Kj�`ȉue1��h	-��9���Ҷ�Upk_f�r@]�q��|b<�E@$z{����x��۴8�K;����SS�⦙V��b2	��1F��ĺ�����rD�:�f�4�j���>�A�C���3U�qB��K]�L��8]�ZO����Q�|�[S��"��S4�CV-W ;��U�-����@º����9(1��Z#�޼@�F�}�TF ؇����8u���A^Z30��Β�;�n�Y�j��T�������&�$�pc&�����q���ə/7�	��bMs�&s �z�)�]�D�ڹ]���w]�\l���#�9#_�٘8EC�]V����N�k�����o���#�������˱�H�2%��U�HǸ��͂z�j���F��lf��+�Ώ|�<�4��W��tH��@��U��a��S�"^��Mj�}����'eY��
�P�.v8]Pp'@����'O��^��[���[1JK�@�i������ܖ�=�����8�������6�J�F�##�����4����~�"�Z
��Z�A���68�O�\e�]�2L��#-�� H��Đ��hmBJmȴ[�//���
�8��G"�	l<5J���_l+�ӽy��H��۷>�:��u�P`
�ۿ�����`@�w�1>�n��2[l�	��DG�A~U�dh߹��*蟋rb�b�0/9V����&Z���\�H2S������ q{<o�ְ�𻮾��w� ���	��*�ZI�*p��l9�D���H��y�<z�cB�EV6�����5�^��q>�'X�3��Nh(v�>Y�I`�r��%��5~t�蝹��q�m��ju��Tc���S��Ɛ`#Xց@�YZ�ֲdo4��v�|)XҜ�ƃ>�V�����d������M����t�QTqcѫ��l���0�����K䞟��3�J�� ���� �F�;ֻ�Aì;~��1�Hk
�\�o��$>��?YV-/�C�e4>si���������}K�bC7�����wS�M��Y�,ȸX7��"���8<�}�(jC�P��9wO�x�������a���<�<p�M����*��.�N��!]�$%�ԝ�EN��UP^��i���#��#�h��c�m�e���zk���u[�6sG��a�2��u�J؆͔����Ά�n`lݘBtp�Q-�ig[��������j�  ,"Q)�j����lS䜠��6eXoT(�כ%��\N����0�3X����zs^���x�9?Xp��~�-^�� �^x�NT��7	!p����T��')���у�Fy�ÿ���&x�r�P��T��HѤ-�3��p��W)�_˓Q'�x���u~�Z
.88����2�6�v��%sW���!���:v����Z_���*}|�?CV��_�ݐhl��,�V�������պk*�Oʥc�}���^M��Q�3���ւ#?��.Q���w�$�r�}�3U,�l �<ʂp�}��p��f��zX,)J-����X��-��&c
������#��I�j5E���#��X�yx=�Ζj��,���j��t*�AV���ۃW��#���GuA�p_�)�cR��"�0���i�sS�;=?���JL6#=�Qi]n���v�݌tb���(�n���0�f��\�-�0u��J�5�ei<:گI�'D#����N�/�m$v�һ,�mڟG�zT<,;�c	=&� p���ـYT�͆���9O�\d�iȥ ��J�w���Ε��G8�B=f��Js�\Ҋ>o�.C��RI���'�o29d���C
&:x:7g*�j��A�tk�l���H�nL��R<��؇r��J֑�k鈱�g,��`�4 ���v�mh}�1�~��F��/�H�^?�Pk�=�X�T�+c��ٱ���΢;�nq︽]�4D�J�q�+lhMn,��&������ۮ��*���D���+����#xj[#��-�W� ya��a���8���=g[["�m��2�EN,7���
-�;BNn,�'?�R�Y=�\�> �Fܼܵ����;�oAc���w�]�lB�ɜ�u$Ax^+����V�i��μJ'j�-��{[e�x�б�m����ō�������;2c@�k�f��'�v�7˩W��T#r>�Ϣą��:Zꙹ ;�u`�,�7��K��5��i=�#��1!�%�;�,%�QŸu��i�ݢN}���w��}�h
,��O��}�͌�Bu@���-q�����+q����"�JG�0�Hj�Ӳܖ����Z���v�ӈ��n�xD<�~"`!�]���E@�ߏ���6GЩw���j���k�ú6n|�z��1D>�|78ĶH
έ��#������S9ޚ�s���_�Ÿ���$����G
{3�`A͗���Q+�@��W�w.=<���+mI<� ��~��i�!3��b�����3wk�x>����_Q��5�Vm�����{8q���J��QSX�aP:��!5�?�Mb��s�.��0���^�Q���QuXY@�$�SX��y1�1�b���K������X��[5�U�㨾�/��~"�����&�� ��/am@�Z*�n���}�,���#�?���-'��w��\^�{lyQZ�۸L| J-zb�/N�Ǩ�f��K�x`�M(��E��F�4:K�8�<��1������Ç_$0�#���5�!�������e�Dp�<���h`��"� ��%e�xX���',?�c���%;uX1I��(:
��qq_.���oS<��64� /Tm�t9R�\��?�^�B*k��lD���b�C���k^��ɚE��*���tJ�đ���\�Zmbi8:4ϔ�L�~�~�xK�0"�o���ڭs�'�mᣖ��C�u]&7Kݡ���;��B�}zh��~�.�s�))�"}����t��j�H��NѓRҦE)�h�%sG˧ҝ�#Y������i�B�-����5v?a�U�tQȒF�׻OR� �}�L꾶q�ʴ��<���\��,^e��$˫|b�|��4�\_����T�+���Y2�W^�A�#�*�l8��!��� �Y������P.Zc]���\E��:�k�c7�X�f)�C���J.�r���=F���Um�zQl�����t>#�D��5����I��I�J�p���{����x/[L1���[�rs+a�mO���X>��0���p���Z�>��PdQ�qц��3R��iCR�v4������(�������?II�X���y,�?Ů!Ν��>_�8���g���:5�2�ֽK^�.�������WnӢ��D�%�#B�*�d���r��@�h���+Q��>�̰����M�z�+��;��%�l�`t��6�8�Q�m�������G��eG�k�Ԍ˚|���E�[ʷ��3��N��*5��?\����4C�����~x�O�y�BB�~�b��������5���	�
�
�����C��ص�>P\M%�[�s��r���NB-=��̘~eؐ�#)�����Ɖ#����B�A����K�8�������v�1wqĒ��������Es���z���^�Z��_iUp�����"��I�G(��2C�3�CH���l]�A|:���Z�� �h�!"ڦ�1�;�܏��.��'��k3�t�Y(!wX����o�^��*��,!�@K������L1����QGN�J���*�2�BH�v����� &+�
 ��q��Bt��W��$�x'�JdM̲ژ(�
�)<"#k@L�H���X9�Q1�R�љCC�CD�:F�-C���5������s'h��΢���sOR������nu��:[�zis�5 ��\���a��t|Ō�8E)��.A 6*�D�)�f��UL���e������a^�*Q�F�?����S�UY"�3�����'t@�M^��?��L[0s��E
����g�C��	eR�\_� �P}I�BP���M�˜���m',	�MhӡJ��܎^8�7q�'�|�t�E�CĎ�F���O��}~���D\�h���ә=���n�H��#�98�+
��r�����e԰�S�3�l"���v��Z��&�5���oK�s�`�ҍN0g]�zɉ�Rt�;�'��p���ɹO��iw�b��6�W�* &E�u,��ѕ'w{��[��a�dH�­+6����e����i��v5���4D�u�p��.N\�14P:�r�Zf�1hD|#^�C�\�,���Ж����������4�T����W��.~'A����>�0���:4M��~�o�w�p�Ӷ�o-�M� ��wR��=����i���{o���;7NA�G����K@����V
�c">Ӱ4��}u���	+��Vn��J)�6����t���<�U����pu�H��f�d�q 嗀�c^s������ѧP5s��c���_m�n0 �Z�k�^�����D][-���d�L��0Ҡs�[����ᩧ��<Z6{d��m�֖O�5����ɗ^��gQ&�u��Y�D�m+U�F�����R	�M�e+Q�\}��Q-�K6I`)����C���jf�`�b�g|Ĵ�Þ|��v�4V� ?T�YL[%�� ����RQ͊k �:{�qRn�#�]��\Ç�e��1)67�Pc����bbU��D���!fFp���6V�OWA8���K��&�z;�A�d�xYw,H������ܡ�dt\\�%��})G30g5�L�Ϝ/�����è�f�F�r&u�ȑG�0t�o*�i[�"T�ҍ�..��7��bl?�d�Nt�����Y�9d �
�Hٯ{_�8}U��s�]�I���|�*4�5��4|�j��I�}}�P���$k9C��v՝}�)���p��,'�R��/�v4��x�%��DN��Վ�� �
���u����V��p�Tl�s�h��s�e���,Ҝ
��m��`��?Y"㋯�T��v��֏�mn!�M<�2%&�d�s��u��I���c>(W0mdp�.��'���@�*	�?(d����X��;]z�z�������{��V��<n2�ͪ;�<z����k��k 9N���"�B�m~�E4�a|�c��4֨��E��fa��E��dL�
���8NN5]��Q9;��)V���0�gn�7�m�����I��k6={E�TO�ϒR?
ƫ�6�S!e��҇vbF�ٳ��d~�������O�U��(�ћ n"\�:���Sox�9zo��ܸog��XU���?4����bIF�VXꧬ|$�љc�f!u`^�k}{�}_�X��?/WJ
���S.�j�ʌ(~#��n$�1�y���+n�ֿQ����t���3�.M��x��>�K)�,S��]4�]�j��w9(��O��]Kp�i���|z|Ш
�|��,��kӴ�)�(g�Jq�/�qK��]���9����H��y�����SP���Ch�i���F�)��`LF��{�<�������TY 	���(R�5�7;D��8��/a�ɐ��Kʜ����"�
�ˁ�2`������:��599�4��l��%�>�C��/v۾�k��{c��\�����S�52�Ej��]���'�+Z�A���ӄ�d�l�d�f�vS4u~��'à��K�yc��B����Q�+G.yj 3�u��I9ycF�����!h+�*�J�i�5�c5�N[۸�����ru� qY96��H��6�,�@n���z�V)p�%��Kz��k�c��D���m�Ըh���5�ӐsKC��;S���A˴#���/9:�>~\�^� ے���t�5��y�H�*��j����ĥ�a�j�+�ig��C.8�`F��+K�-�$�'�u�{�u� � V�����=ug=4��O��=�D���Zh0[O�M�z�wĄv�s{�a���g�8��ݗp��|���^�;�}�M�Y�8
���H��=��>�xƑ�n.P�/���l�=Nh�/q�L�Ѐ����b�Y���$���W���-�|��h7����sA�A���k�;k�M���>��F����`�71c�i!C��I�*�ׄ�%�7��L�z��4Ὁ
�h��8;X~��-���V�_��J��f{�t��Ɨ-��·�R_<�U>�Ҫ�Zm�~n��~�H�� ��]i�&���&�����+ ��M�{���}���0fτd���-�<��?DC�/h���e�t��{5��@ 1w4eLP��Q�̽(�aUmQ̸�֖�m6�x�R4�i��/|%��>t���Gu�3��nm̙шWh#�_l����K�7b�u+5��4M	���csVծ��nLHq�w��?Y_XCy-=[������L� ��ty� �7_Ǫ�ӛ��Ql��vN�4^��7�lq���
m��L�a��G�d���� ����)M�H|;��O���ǘM�����0x��v������?Ĥ�d�����F�d�A}�F�_�5P)��t�XQ�	)��^��-��{'�ڃ�Vܻ�;ɂQ/�|���ϗ5c�ɫd��M<j`G-�!QfJ�7���{�0�;��?\Q�	!���IsJ�W?�O�z!�А,7&2�v�N����ɡ�/�x.n>��/X[�Ɠ�^Հ��q�e�5�)2�c�7UF�z��	�<�ʝ��L�9v»��>7���}���ɾoz��f2̀8�k+�_6>�����vY%���uX�H�S[c�5%�:���26�� n�5���g�jA���Y�9���EC����3	�(���ՙI�e2F��=��'�k��a#䝄�Pպf�Hy�5b3+j���A�G��v�� �4�Cz���S�B�ѭjQ�PêӍ��7T���h�\/q���4M�-v�&6�q�K��=�zsg�����V�8B�
�����݃�lU�T����+*�T������� �#ɀ�!�A.��a>�&d��WK>�9�0_�1��0���Ge�3Z��>/+^wZ�v�KG�ܨ���z�ϡ����{�R7�=�'��]].JT+RH|l�"K��ͣ��)E`w�PQy~HsP����TO؝k0�����WN����k�<�pq�L�#w�E��ΐ5)`ұ�:a]]�v�6!�/�c��WsE��!ן|z�M���u/@' ��;��h�'�|��*X�P�F�`�H����$5����������5�ܱ�[� q�|��*;$6��c�ֺ-�nQ�Ԉ�,-/A��U9��ѣ��Z�gA�"���.G1�~��%X���V��9���H� Pyi{_��:�C}�6�Dr������,C
.F5��t��(���:AYCNY�-��\o7�M1q3,� j�������k��������,�v��e�XE8V�F6����v1oV�x��
�G$�Ho��9����їI�5�5�1F&�q?�c�N�|�k�{�;ku�%��> �@��<�4����$4b��C������� �r��j{WcN�0 ��R���:��_���)>���]4Hr8�4��u���;zT6��H����]<ݢ�����W�Kc��B
���=���|��N.k�I�1ڹފ�օF8�r���Gy���,| ^q���A�ԫ���=�)��w��̽�}(������#J{5��;���Ğ���/������2���Fm�#�1�Y���O��[QF��Yp��B���ԟ��:w��>��7�Vt%Z�8m��5�ET��i�k(�%��j L��g�y�vH�6̇���#�
�R
�C��0�|	�2Y�W5� n*~J���e��s'1����:�b��S�Ra���	!�	���K�2e��ICIu��=9�9	k��ܾ�HPW��y�>A��3
��D��r�s�+����5	h'��o����qZ��f5���N�����f�6&۔����L�a��%�����{��;�\�n?9n�$�\�6�Y"z���3���u/�q��`a���t�9�Iꪍusմ��r���Y�d�⹪~fu�X�N�*�P��P�m�	[��XM�.Ϋ1�'��Q|^�t.�U�R4��?����nxeV�1E+S�U�#Z�C)
k�2M��ҋ�5NN�wJ����7C.��#M�J�����G�أ=Q%݋��,~w�:�j��t�27Xd۴-bH4.����m��P܂.�2�jb}&eI���{H�-M��F��k[�K�.d_�ҭ��� �c@�a��(�Z���~���\g&*0ۻ��{�{x<�xL�w�a�$����� ������6��r���b�d�L^p�^z�2������gh}p�7"����=�!������q�Ge7����y��?�GO,�ғ���!������P�<�t��lz�vf�T�u���DX�B�t�5kK����9�ދ:�X�!
��WXИ|�����(��v�I�C	=�8�~�)z�d�X�{Œ[�k`tPl	@�U��o}�$�JT!�� ke������g`�x�/�`��Ҝ������|⢈�D':Zk)�Ԋ��?�^�����e����~G]$<h� �ƇG.���O��,���n"엛�Z{����SFNi������9��¸��)��R�Bi��p�oG�z�9;T���~48RY9�+�V���3��_�^ #C�@�j�� )��4
 B>*��corF'\΁�q|�^�!�O8z���v��?:�@�#���<���;[�)���/l@���_7Ѡ�� �����݂dF �/�8�{Z�Qu�x���C>�'�2Z�����u�{�K�K��=&�[�HN�h9�2"T�Z&����FK�$��d����l��X�̴"Ǧ�D��������0��,PĶ6+I=F����Gš�r�D��dyP"M5YX��b]mYʛ'i�b�Xn�ѤϞ��Q�Cr��e�aY̿���RT)�/�5t �*Y|��Y5Q�=�B67ӏ�æ���&�Z;Q]����@�bglX�ʆ&;�����GSK)Ut�zL�`g�8��Y�<T���h������+�5ϻ.
���R �%���� �2.��\��R��
X+�ˮPْ��HUū��m\~]lKN�)OԈ��p�n4��l���p�ỎĿ�/�q��Y$�ȧ�;P�d$H4ZZ�~<1��p�l��ӝ+�{R�����zɉ
΂9v<q�
ܸ$Q ��U��Q�u�D�JZ%��ӓ ���h͟][kg�q��U��٫ta7	���&�sJ�	��⯂ïSMp,�0��m�� �&�]A���˖U�������A�S�k���>�"T����-?��C t����;�'�x�FL�P�嵇�"x03q��G����zf6�ǭA7�	�1�=2�ԍY˸G�Xҭ���+���Z����27���&Ŧ�xQ�ӛ*kRFp!ը�u��C�Z��̯1*5 ��>�(_~b?qX%��ur;�^��;��.���j�1a���C����֊Pm�!͔c��J��j�5qf?�����.�Q	�(*m������"�صzU4vGʰ&�&竮��r�<�`��	��ݯX�5�(=�Qsl�#�N���"�	�ש/�l�a��?Th���L
�2�]ͧ'+�썏�1U/;��urq}���4l'��� �����T/_�2a�p�am�-1C����� 2��-^�'�%�s����y�di�q\�B���	@�Ll�4d;ċU#u+��$ٕ�,�=k��v�ͺ����H&�3m���S�Wc��&�u�Cg�J�t�s��m�̈́<���P�d_�]�� �7;B^�j��Vo������,���rZg�N�e�e'����[Uh�;��a+.X�8.���^T����>�AӔ8�W0�:5p�*����#ava>ͧ��1�᧰-{���l�����F�]ȟ�����-���h�� �h�
�|<8�[�j�*�@E34�;Τ��,��*�J�@�[����F9�uj��֭�?�z5���B�R z��$��sD�`�Qed���:������U���p��K����lktRM�[�LC�Wo�T����YI�Ñ���2��,j<��*����$7�����7�w0���ڭ]ߚ��>ڎh��k-29�},W0?�9]'�4��!���J���|+a����/�t��G.G���)�R]�]t��'Zb���"qx��]�|w�����]"�Y#�)���
�EN��Ⱦz�^�^����@؈�.(��]G��5�`����"�U�-B!^S}_&h��Sk�k��UdRi�>�J�j�1������Q���'%X�X[aO�J�}���/'�_E�GN"V�b����)�3/C��#�^��`��O��d�RsĈ�C�q�N�v*\�ٛ�}�6� �� �2���K-"jVY-@Ё䝤8e�����"��+1�����D�ְ�f�'��P�>�M�G7ݙ^��!�|�'�����IS��g���R,��>$�y���$�������Y��"u��
��!I�xɸF��oо^��ґ& �r��O$�~9ק�H$�HGؾ���i"�?H�w�~�!Gt��tg�4�����z+��*yQڂz�Ѓ,��O v��yCu�4E�� #U������>�\�p}0����؈1�+iG۶v����]f5�(��V	�T+��F�U8�*\k�NTN`9��#�q/5�
���|�H��f��_�tU��"gQ����|+��c��o�L�����P�jOi�WGJg���:)9�z��aæ�}P��G�4Y��&�b<$��
n�*o�1x���>����M@��u*q��P��T �g���|�00D��<3�R�4z��.*�����Xff���FE购7Eǥv�E�z`X�7Y]Ԧ	i�ֻ�]H�N�s�aE��k:���R���ᓔ֪t9�- ��6u���d���M~�<>��m����U�ˤP��N�%� �8��:��em���C�UV���ҏ@"�1U;W.��!�T��&�]	����}��?��4�$�KT�pq&�/����{%e�,I�A�ʌ@��]�/6��,5�TYſ�*8�ri�s�|��Ȩ�(�Y��[����7�֢����܋q���n3#�n9-������w�BnE�7��g�b�?�&��24�9&�[ �k�[��4�c��ZIV/q�%z�JV�[����$��..l��Lu{��n@�Ek��S�;��'4|y��|�?�?�>�ŚW�LE�⫋����3���%K��1O��6�LwhA��Fnn�=����4�k���Κ�VG����|3M.�xsG�x�m&�;�.V��� ,+74���NU�*t�X-`go�Xff�&(�@ǭq�A�Rl|"�F`y >�������fL/���I�	MC�zտ�(��$��g���]��_�D���,��~k����ԉ�\ZYtJL��鿋�qɜqGa-O/t��r�Kj4���!�>���>_�U9]��=ҳ��,r��ʂ�Mk��X�ǘ��	��8}�;r�J�c�%���W٘�LZ�\�<u��8p�aWp��o+ �N�յ� p9 �K��H+͌P;�2��H�k$~���(!�s��-�����#�N�5�fL��J��`�Dǵ��.D"<���o��?4�3\w1���f
1F�x-�t8﫺��\�K⌶�iUq�G��6��p��&�%蟱�lvENJ��rnU�
酓�4�ߘ�3�S��fP��{N2+ ��U�����i�%+,\��G3+ol�
41DI,�r"}Ԅ�g@E�h|dBf���u!�
�d����E#�S¾���J�SJ�6����y��h.��T�<j<jau������+��)��!� C��7�^����w{��5�~��|��ۅ/��7Qp��fM��	���&��c�Q�Bd|$�t^wOT���^�ר��l��xԟ͸1�3���ŝ!�cK#���)����(s'ޢ�{�; �}r�l���bQ�ʖ�\;ݘ�Sք�c���i8��~�v��ݺ�t��O>��λ�'`-��g�X�*��S�9��%9�a���w�Dk��_�$ ~�/�/�j\�<����[cD$$�V��{�+%�C��&�{/�2��b#<J�8E�</����^2>�{Q�9� .�7'�(u"�t�U�F��y����,��
 ;n/�Oּ�\��0����;�3�Q�U���Y�9�����`��b�b�R�ߣ��">?p�:���N��%'������e\�n���L1B��B!�)p7+e�݄��6�)d�=6jo(�#�zH�����i�|��#	F{f��� J<�i)��!�a�Bٴ���T�L5+�8;z�d��z֔|�~d���ֿ?�V��5n3nB+�R�i���Q���1��O��j˝��� Ƌ��v�½�HA ��8��D\	L�����ת��d��h�u^��Z�%�1%��tx�.�'/�}5�9+�'g�]���	0GO�o[)[�r��h�df��}PMI`&�T�v��#W���.�n.��V�|dj����o�x�9T�{G ؼ{?�|[b��f�i=kvL�0��a��H(<M������8FK?=�%��ue��a�O�����+-�b���.�m�_}dR���!r�Y1N.�Y8��$]㋉N(A����R�΄���;p���7�A���;v(���-+,'�R��X�8����yN�+�Q���e�,��mW�^����L<�/�g~n����j ���g�@h��������ǽ��}|$�㆏c�yM�9BC�Sk�X�$���Ȍz<^[�c�K�V��3�fʘ����3< ��]�LO�N]I�0�ZShf�c�kB\*	��]�M�9��g� �N�A�'��r�o��p���B�L ���E@�|�4�8{���8�c=^U���#�q��T���C2�-��a͘4�P�TE�ѯ������ApdȍѨ�LYE�OP�b>0w �B��|.�ɉ~�Če��zV�=�C��o�8�j�
s���N��I)���.�!=O�y�JM~�"����췥�9������j����S#}:W+��+����Dy��*�`Z��R��;5):�����|�e�a��%���Xg�E�B6j��$f��y��G�\U�����O�l �d�ƃ� ��{C�~IP~TP¶�ݿoS�>���	�1�_�	�0">_6h�g!Ȫ�1�+&#�m�N�Э3�J�4�x�#ު����b��0�Ë~j�P�gñvױN�"3�������D�K	ϮͿf��3E�>����=M�)���_���!��FZ2��� ��Ch�?�=�,������E������0���9߸_��4}�ԥ:8a���#�o��Gl��2�I��e�Mg��{�-U��!�r�ji�~�4�������
�u�avN��XH��";�� "����C0+F�Kk2M��B^B�'ߖ���l�0nS��_e*OEk+�-�KD�LX�|�Y8��!�F�bc;�Ѿ&�A�����Jc}��#�C�`R�G����,V2��2m��x`(ױ�J�:���)�`���7ܢr<�Ĵ��~o� JF���}��o0���*&�F���c,���i�I�"G��[<6�48]�����P�M�]ǐ�.Y��B��DB�qiZ߲�`"���r�|���R%��F�)�Y�^��s~���AG��u4��E����f&�s�wG�!������a���4�Yu����V�
Y:��c��-��M,���zQ���9ɿ�d���Gz��=h�l6��zz�e�>���K3�&�7��/e� 5��A�$�w���PS�����lC�����c3��j��L)�<C�;A����]
Q43t��I��q��C���� z]"O /I��TZVR����,�x�o���A��W}����}�"v�M����L��K�
<A���藀{fiv'G�6���J-���M �7�!���!��'|^����|W�s�XvXB��ݶ�]���MWZ긑��0��o��k���*�<���s� ��P��1���ͥv>���G�o�N6�&���'�CJ\�nS���|��bpϙ% "e��u��H�9� �y*�Gn���;��*���X��(D慜n�C��C����X��Z�0�U��'1y�	}`"EA�	��H�zc��X��-e�>
�޳�f����������~��郁��oS�0�ȳ~p��ZP�{NH�����i�>uU�~��{��<ny~З2�W|�LΠ|��d���5h�h
���[f�+ů��6ed^�h�w뷕៮��g�]�Q�\�n���/�'w�K�6B���b��$Ԅ���o��Ӭ���X�G�6�Bkω�W�!����!���M�U7�������-��^��B�OE���>ZGǻT�Zk�����{��a9�U�?յ!jY��I�(���d����8�A�"�+.dT���[8�b@if����$LS�t7�N�M�\�1Vƙ�-�0dyi�-xB�=ԔʧR46�#�ސҍ���mE~�G��>�.�2�J��^ ?5�8؜,�H��)yfJ
��H͘5ŧ@C�x��i}�yf�o��jHA����/����(��i���Xxa��E��bTPR�G�6�k���( ����ygb���k ��M�̳CX�c�9�27% W1��e�ʣ5D��g'>#ղ�P�D�5��Ț�K�C�8��`�gk��Mx("����dY<�.�+��t�J)8E"��=s��rV^��y�`�C���S���̖�f�F��@G<	���Y�HH(!�^!Q(^	=(�x���G�a#��U
��H��(#�,y�u[X��f��yq+��0(i��	��E�Y�ؾ~��zg�6OD.!���cT)#�qF�,����)�i������Qn�]JM�DTI��ᷪC �5����K�It�w���͒p����#��679�$��K@��`�Fsmէ�S�n�
d&F���iٲu-$���z��'�t]�Jw���t�i��4H�#�i����#��K�,U��c�}�"��@0�b�w�ؠ��7�*���'�����;V��iu�/QD�Iug�˔�:.Up��b�wR��ܭd���l��0�ز��9�ç���7��H%7���$v�����AK͓��p<e���#᫿�����<,�D���)�۝J�Δv����\�ZB��&%��ǇB� �n���!p~���#<$�rJUկ�����Z2�?r+dg.�D���������_J��{��R�>k��ʰm��һd'������~�VO'�@�}��0<�֋F�q�
���;}-���+������N��P�3 ���Ѱ�9U&H�U.RG�!F���F��'A�7���7l��@�@?;�& ����	���3�엮���#�qw��߭v�sɬI`��1w,P���3F�΢�d"C�X�s']�
<�Nlvp�!'X��n���}�4c �ڎ��t({����Œ #NPcP�~�'�HAxC�>?O���sʡ�}��(��w���	~Y�>v��1�)�.�1Fi?t��֜2�phS�ƱE�eA6@ˤ�x�d��J�̓Ac�I�%)�D�:ه��S���,����$f�+���S���!	��b��Dd䠀i�M��겸@�e��H���xY@8�$��	'f��!$�jԲW����?HWq�Z��M*�I�v!(B�YD�e]ط	Q��1M@��w����|`w����Rf'�}\L0u�@N���dH)����>�\B�`!�%�����%��x [i����4�-�+�b��Vҫ����靺��p0W��U����%��ME����/^8Q��׸�ʺ����E�� �)�g�7m�iK��C���и�
�s��=�����s]����K�;���z����S_�	H�l��Fү�+clkr'���\&��`)6Ej��|�>����j��U|�R��EK��U��y'L@;��+!l�8N#���b����bW�/w�l�/8���E�L7���#��]S#�	H����Pj}nd���C��� ��#5���I�o_�|� �C��X�}��8^r�CƮ��_�>
1��Ӧ-��O_�H��uy_è�f-}V%9g�|8C:�j�C$P���=��Ő=�Q
����C����6].�c�:��:�/TJ���ϴ��c����:ݱ*,0�}����b�B�l��k��;a�_O���w5пYr�t�{�l	�@�\�Z��L�V��X�OMA�P�c�P>��I�Q���Õ+̥�9X��'W�#��M�� =H��Jg�0�Sj�7�>3���,�!��s�uh���X�Mw'���N��ϙQ����%�$A�M0]���rެ;���<��)_�R(��\ ��~�m��HM2%�gA-���p�b�ˇ�%�2Ё>L|�B	p ��w�2٭�I�J�`�Got��IZܕlX�x�A�8���K�ayTB�w�(h�]�wy�q���
!o78Q���6Y�������bὊ3kp����|7��1���}�R3�k�R-�4�jHtȰ���1��oU��o���8��G��X�� ��H�7O#Z3�;��9�}��F/k-��@�S"��WZ��y�?E�����NΚ�P:Ҡ�9{��J�w-����1�_�@��w��ZS����#d���#8��iX��Q#@��6��AS��j�� �A������� �+հ���ɬ ���AvH���yV�/i������� d�:���=��D����A����^���6�*5ūs�U�;I"��L�o�S���x��̄r6D2��A!t�,�ލ��E6xX��F	.��sa�6���?tZ��T�+)õ����l@�i���\� �~U'(A��j�b�>k�)�x�B�v�3uj'��S��G������a"��G�'��JU�S� >�u щ�7�B'��l�af�+��=%�;601�:�����G�rMZm��g�NP�yV��n"�Sȶ�k>1����y��m����]�	,�-Җ�a!�����'��2�ڏ�H_ �D���.�R���^U�@������h�R�+LrO�g����k[s�	�(;��� x��i�N������Z+�D��!��Q���`�8J��{��9�c�Go��E����z���>^��.�4{u�hmO�P[�X��}I�!�����FAS�:�=0`�b�۪���;�K\�:�7�(���D7�D�������|��EQ�uzm��n�ZDY����g���R��.P�Аb��W�u;��5q�%�S���E��`��׉ϊ��8��� 82�O,�}�e{>V��y��M$�����⮛�_�;�[k�����Ns���瀋\���I`v&���ֱ�MV�@x(��U�v	�b�(��p"NV�/�ȦxH{��uG|�f-�c�>� Y�f0cI\/j Sɵ=��R��$р��c���d�R+�D�H��*2�7��,�Y���Mo�Ɩ�߉�EQ�ECҚ����~U��gDu�|���F�4�nM;��z�C�25}d�]`RIt9�37����}5��\�1�U�|�ϯEh���:L�
���7��%�������������ad��b&¸��������Z�����B*پ�f�霄pPU}�$S�8o�U�74ԛt��&~�Ο'	����e��B��gG�]B���ڞ�j�0���T�;��� 󡪤�*��S=`��O{�%�6gC�T����@���,3���D�!>(��?�~/����*�,{�OF z/�����E�Z!�HxYS��Pmɒ���EKT�5��j��Cr2�
��{VɅo�Ak �4�%��lh���T�]F$z�ᾀf��l;^��G�x���C�=�u۵�g����8���"$�V:,c�"W�L��IR�^�>|���m��1��������NZ=x-���|����;��<a�x�;'b��zˣ����̘d�����^����I�O6S�!.1N�YƆ�wNH����	��I�a����l1�tI�Ti|x��n=��i���xM�����$N�W��fB�����ؚ�&��< ���!�,��x����T���p�����p���/��I_����w�ĥ���)f�יb�B�OX��f���/�G�W��bUߎ�m^[�ak�ND�񇒹� ,d�0!�(:��-m�5�6s2"j�v��Q��
ߛ���������x�@�;W7H��}��kiZ��-�Z��DΟH\�W' c�g�� ��qr;Va�w�e��)il�sbT&��aܖP|����m�9&Y
���Fg����W���q�w�T���q���
AJF$�a�&4(���蕐Zg�b׾_�}Ȯ\&�	��VA:�DMD��p�15��(�P�
�`�O�Tfg�\ ko�7��'�s��(�'�������慆�W�y�>�q]Kˏdh��{0	K�Y�:�%��'�#h��@��Ga���l!��z��l�D�~s��S�92���W����#�
�N��^�t=�nd������w���kC��ayj̫|�4Vkڪ?�h��мgn��nfg����u�KR` ��.����l���-�Ƅ�x)���\����|��n��/���q
{2l���*���oKo9�Nyx��DK��$��J����=l�B�o�S�ȢKx ��`�4ڎ�1V�����0����8��!_��r�`�;������n�C��P�����b
G��P1"e�	����֪'{׫�g�����������|� ��F���r��C���R�㤟7�L,9}Z)F���\8 *����ЙT��Z�x���r�����6'�g�`U�:3�C��+��T.�ꩵმeP��uJ�?U*��P���"�g�!U���Yl��B�hh�u  Ea6�\��i�j�n�ި�D7�� b�*��\e�Cv�&t����7a��-��"ϋ��<aeHk�[G�bۛw�,N���O�fA�^θ��&�R�I�P�&�o����b��*�òpW�MB�^:*�Y��`薏/��P�	�h��*��62�����id�_�_����z��fkHg]���ٍ�Z��j�
J��W|��q�,b��l��O�����u7	���X����V���gu�@��Y�*J�K�����s	[��bQQH�x��Ԫ�VF,^ꣀ�h�p�^��I~
9��-���ѣ��j/I6l�غ��[�޼�d�~�+ ���W�7�4P�֫����q��~��y;NM%�Ǫv ��&�/^�4�aݮk&1��=��߉�G�Ĺ7d����3	��)-;�x�����1�F-E=��p��;5�g��<lŏ���;ՠ���TM��� ��@�5�اH	��Ň�,�hц �L�z�-�`@U|BB��;�C)(b�Ҫ.��sLzX3��iF�$�85[�Sֳ���QhX���ZK�$�k�Mz�U����u)	㸟 fK&�&���ݬV.v��Ҍp� D
�2�
��fG(��2�˚W@*�?Y�����o��>�Q.��gT���7�a���w;��K5ߖr�н 9��Q[��S�#���p�ϩ�e��e5�6�c�zE�vE87+BŁ�R��$� _v_٢>��Qx�	x@��{ɿMl���)�-�\*��R��x �?���K�$2�~yٽ�����-��o��^G��^�7zUFf�P����oI������ʄ�H�-��ƙ�o}I��g_Vҝ�&�)Ӻ����F��ق����p������J��H��8��udM.�$9��te�[��GSY1���\���6.��'{��I����ĤFg>�Q+>��Yf���b`���s�0[b��n�K�Lb��/����"�e�E���i��Tʪ��Y���Op@��1�Ћ~_.�
"Ցm.fN�S�g�/Z�_61,}G��BmkaJ�Ձ�Z�1�;Y�U��ڡh%�68(ݧOf/0���1V �,�C)�_�#�b[��&N�q��I:뜻���ٍ�t�[�>���/������C����,H%|�g���W��8�������Fz/�� :�zۦ��������R�:�??�B3��í*w��k�I4�Sp[�]���V�𨛠�m�ˮ���6�u#�gB�1җ�w2>z�Oߌ�����~w||
�n���M,�E���uG�C��C~U�,��О�X�>B�������g����,[qg�H���W$��숁{�7*>0�U�2�-�q�TL��L{� l'`7ؘ�����؉"��(���ϷW�Ᾱ��.�_о���)����>��HU� �w�YBk&L4�����	���Jӱ�rvA��H��,�?5s������D�v.�c� �cA���a��3΁���c��:��� ӯ��jS��s>v��F2���ØD��wS���H��M���)�ԋ�
���L����nݼǈ���J˂�
��%�,ĞA�~��ڤ����R@F��ek+bT�y+9��<�2L�����X 	�CUMiZ����=r��M]�3ؤ��;X���Z���Y&�_9�auS��Ҷʳst�D[�%׌�Ai�i���8s4�ݩ^7}1KPv���R����>T����xj�_=��t�����\;o&l5wc� thL���y�z=�����;YK�L�$�*ϡ0s|��J�S�ਐ�-�r-{;K2՚�w2�L��70�� }�L9��c�5�� ̖;4J���U�ޅG�+�=A0���aG5��W�Ҁ�����|y�]�8��ߋ���f�}�w'����� ?�=8R� B=љ{�#���'>NC�6���}.����~�<Bsh�tHocGa�_���M�/%�r�Ԥ�, �~�8��!����\������ˈ�	���V\st�f�9aD��l��PZ�6��=��6D�?��6��
������1�!Fd�:K���XP":C0	l��Xe�d!�n /t�shF�˕p��<R+�i' ����<{�"p�o���ڞUp�Pm��uZ��s{^fN��ρbr7�%�.	��j���Z>��k>ȱ�Zgn�o��� �e��9>Ƹ����ʓӰ����ڧ��ťׅ�L�%�"m�ai�3��~ބ�_{����V��	;���cv�+;��fjX�߮z󀓳�T&s�'i�Y��
�E���;�T�|��@�2���Q����<f�\���Ta&h�~�׫a:�U�g��cOxӎ��`˵��@�Rx�v�7�}v�7��/3�&z�I/o�0�%�1�}�]ZU�|��"��=F��àn�,>�UmAM͘eFA_�> �r�ۻ�0@Ϸ;8	��#��a�g�b�EAى���u��_�ב�	�!+��$E��]HE��s8���������ַrJ�g�?���b�`'t�W�&��A41�%�'⫍�X�b��<NXXz��:\���kU4����3�P���k6�J�X�l���զӠ#[o�6Gp�I�ii�� ����b����vb��9���@.h�q����O�]�H�SSz�jE\~2����M���e/��p�� �\Y�B�$%fǟ�:��ﾍ������'7ߚFsZ��0��O<
;�����2�3�����D��� ����.H��#�\i��- �ծD���5�6f�[í���b����*['}�KBLs�!5�9 
B^@��Un�^�ٵ$�C̕5l�k:kv����2�_���D��)L�s��,Rt�r�-�z%�@zj�J�/v�C�2[My��US�{�s�Om���~�M�������b '&r�>ȉ�����+@�UO��z�Y�μ�=��|��'��vu�~a׵R�7�h���/����h;c�P����Afo>�@W��B�޼��aS���bCJr�9hr㦼\����"�.����}��]y���W�hTD�9�֘!�d�n�!'B�~�S��ni�6���2�_g��LEEs��o��#���(d�ۜ&�C]Ih��;����}X�l�3�N(G4Q�z}B�� �_ӭz���Y8����=� �ڶg�z��&�K(���V�bm��!����~�g��,ڵ{}g�?ƌ���#ơW`����܁���Yx�6�W�#>Ї��=��E�J�&��ZS=(j#~���ey��`)WWk�r��I�d����>6����tP�?�d|TgBN��v=�U��i��qyXk�J!�J��0=m��ɍ�c��G�7׮�=��Ln�H]�u�FF4���1(igpx�s��p�����Jh�..��I&`���6*ĺ�8�r
wĴg�]xa�-�u��,���f�=@�\T�9���l*7��񥵨V�ؒj=̈́c�,4�-�1�،��g�W�}�Շ�HXZ@���x�L#���-?�kL /~�x��1��'�?�Vl4��"�Y�K�I�i��UX���~b�;��3TLj�ι�Z�*y:��wN�9ϮQ�ٴ,��.��+P�P�/}v��V��`����v��wI�"c�*�eW�����d�U4���=��jֆH���s�X����������ū��+�W�b�_�<�$]����o���N�uS�}p���?Mp� �_�@]9I`�"�e�!���b�g=��+��}�N�vY�#)���%N�z�A���pQ�n����l���d�m��9d��W��=_�����rH�ԑ������Ũ�L�r3�y� �V>�a�~7���'�,sj��H�sVA��o�	y����a�G�ƠK�Ԭ�n�9W�j��-���i�B�"���);W�mg`�v�F���/��2�&#�L_�_��g��8s@�s{�pY��
�^>��
�)](I�?ĳ��H��}�Gh$��؁�D��C�M�I�bl�}�p��5�ByÚ����v2v�B��u R��T&���L�;x� ���$��$[��^�Q �ǰE2s}�(�h	�@\��T6���vS����3e���&���3(y1�ɦg�,#��s������|Qm�a� �Ej��8%���~Ax-0����}�%��	^��!9�ܥv���?�U��;���Q2)t�MK�M̮��h:������8ƴ�*�s�R��B��IZ�ޗ1b���ãN8a�8��c>I��sE�B4�69kߪ]z��lH�D�#�Ӭ�����tt�YXW��~N�r'l�I.���(QТJ���RW�ׁO�w܍�^I��b�K�L6Ҍ�Z���͋�݃����Zd� ���휨��G�~H����|���VK��*M�ѝ��M�F8�^�<���=TN\d�φ�z�͓��ʦ�2{qg9�W�}������d߶o�_��(!�O�"B&�c"U�R�w��g�g�ꀑ߻�W�PGVwv:e�,RS�jKխZLq�{n2:�v�kI&������=�vA��4+�>F{��(����o_�b�k"Ī(��{����t������>%G_n/�ҿ��}�f�Kj�U�����8_��fI���L��àv�r#�?�~ �H"?N
�F�=��4��T��\��Bt�#��t�������΃��'\��qt�Q�=	 �xj\�&��a���y�g*Mu����2"�k�u����䨫>�k+I�ӎ7q�)b�CZ�75t�n�J5�U�b$��]�f<����t	�]���m�a(����XD[�ǵ��ٕ���urv�*H��+��$��@��˷�/��$��I1���!�lJ������h�8��E�'6$w��)��9���D�_ၻ#�}��]f�	)%��X����I���ZqE��R��lۘ�f�@煱{�ơ���5��М A;�N���Jm�v2.��mVX�!F�Qj����~Gq�7�(��ſ
�l|U�'�Gw���B�ԤnI-�k�/��F�'�1��!�Pa�����Hs�����>O����]�*'�f���yWӉ�c�/�u�\����hr/F�Έ�6܉0?�ͬ=g�R��������u�N\ ��e����g��� *��1O�T��ɦa�??_�����+��]�Ӛ'	��^��.[��aCڮ�v��(�kg����f�Yts�����t&"7�{�F�x��D}#�?�)7��5#8�A)�0�}a�����R�#�^�Y�x����+��zo�7A{�΃��H��f�[����pK�K5Pr���p�q`�x�q���c�C��{7�nZ���_�<`�r9v�/�4O�����I���,�x�Ai����|YXqx�(�x!����)���[�OC������c�6�e����@3yfY�B65OL�r�����-�=%y�����tZ0u�&�Jd�$b��9�S��T�9��"+oD8��- �\ ڨ#�kA8Y~�(ᘖm��E��a�����Q	�	K�Jw ;h�����$���T$N�c}{Ži�ml4�eC���,V�[���2"�a��[�q�j�g�\ߪx5�.�p}�A��Q�x���W�Ű��߉y?" ���;vH��������}[$�Jn�_6����o!#/�w�5z2cM�I�0�J[��-
���뢪�W�C������M#�F�@�A#�ӡ���X��7�đO'1����b\�I��*?���n��N���#�_IiDM�
����q�4�����	z���""��W��;�Շ]~�ۃI���hE?��AJkv��#:b�z7!�V8F����1�������<Ԁ��B"�����i�m�c�L�����ɂ������Ț��7��@O�!��"#74.@��]�D5�Fx��x^Z��ED�j��g�u'	I?nc��� �y��l?�gGD{Tdz�F�EPn�gtr��P��1Lд��<���4�lu���$bb�ψ3�	Z3(����0�+�Cp:� Y6�Kx�u/{�L6y����jk}�h�ڢ�Kp�ӊ;�P�MDNm�5G?C�<��[��Ԅ��"<_w0> =���YU�3�3-</̠�u�\(آtY*�A�,3/�$���9rh�?P
���?��L|�\?U�@z�R^pSN�#�9�!������+��0i0���EB��h��o3����M&�%FT Uo�D
�o{�`�tJL>;�,�4Y���.AB��*��X{�~�֑���D��w���:dj-��v��A�}�4�_��@ft؂f>vv�3�u{0D������6�&�d��n�WSM}>3p�
r�x}0�d�2Z4��w]=3�+�{t���=]	rg�+	.=�o\���?�F��R��q��Q(g��F�h��|nw�+B�]	��:�s����'��=Gc�z~�F!_��L�0�&<LA�r���(t+�GQ�����F�@��?ʿ3��60��vcs_YZoJUn,�*l�+{ܕ�����c z��m�TIE)��+�+�KƋl������F8�-���_��N�䐻H2eꛭ��ǹ+t�k3UcfGUL�{�O���A2�����$��/�]�8%"�m�-&���`
胆D J��v0�O�Y��n-�4�R]�\`<�w���nv��{
t1�ܲ��N̈́�8>���͞�V��$lU�
����6$K2�6%��?]/��'hҫ�@ �\�Mb���^�s�L�ْT+ q�1�/����X���W�a�*~�v���BZQ(<�3t��������\��'���ZSx\�UtU<��}Sx!*&e�➖����)�z��6 �,��bdU�� >X{*S�
�TU/#|9�ԅ	k���6W��bd`F��cS���V����BӇQTq��Ŧӣ�񕋃�oئТv��,���w�hz ��}�����/׭�pF�b�0sv'�t��p��;��s���6�1��,@��d*̇����?"�30K�Ō�i�D�X"�n����6�;�V)�s�S�0���J.�6A>��pcN����ChҦ�����瑡�&�l�2�/I庄�E��Iv4�X7�K�?~Q���� heCW�6����\�>�w��NU\N���Q�]ʙ�� �Yt�;@�?�@�v)��E1ujn�#����I,\(��[j�������J�w@���b��#��r@��ɟT�R�I�7�7!*.(u>@�%Cz[�^I:+�4�<+�\�\�J�t&��5���*\��֯�.���nJXSC�"���礭v�Y�y�g4	�P ZU���qm/��A��H��'uE
�E��Ё-�r#�k�����lj8�f�_���X�����������*d񄩗�r�|VWSr����T.X�iU�{�\'(I�P��&2�*�{s�F����J������ܢ-��՜�+�bZH�<��$��M���}Z8�m�B.�3����~˷�H���{�ؐ������4k�"�k~��%��(�Ҝ��`Л��Z���G`����6n	'F�X2�$��;��XB!0��-l�U�^��1|�ik=�%{?��앶�i�F�+�19��ϧ��	�^�F�-/jŗA�EH&��c��Zf�aT�E���Qǧ��?�>u�;�$��?|G<�Hh����ڐ��sn]32]���d#Ftiv�.��BY��9j��Em�#f]�8O�0i��+U�U�6�2�T�d���M>^��-�M7�h�Y� ���BQ��t3�r(c"�tK�|�E"(��O'e��>�W5s��Y�rɊ��3�`���K��~����_H��S��]dLB�M�>�uB��ȳ�r",R��lc�?ӯuL[�֒��<���=��5B�'Vm���:�<�����+5!+�T��L�z�S��ʻ�9��o�쬀�^�))�hj��W��W5�t���p����z�js���!�c Y������ذ{jW�kܓۃ��n�Y��c:�����Ak�b]�Ld�і��TI�旁`BTp�t�Cm��CN?��E�S�� �$�Y�ٯX��=�5�ӥ������JYi�[�o f۫��
�6a\ב���;1a&O]�h3օ����_%]��C*Ȝ�ug9$'����i�z��غ�O$���I��I�s��e�9��`pLݭA�ۯK�-� �q@Wwg&�r�I���fE�5�=�i�����yT}:�t�!�V�AuY�~qѽ`wr���[�fu���،Q��kZ�d��ҍ��nt� |��s�z�����ıi�C�0>9F�o�6ef=o�7ۉ�����V<:-�q2�����2֪I���S֋�8���̭�L�?�.Kw��KҸ�G2�j)�끴j�>�Ѫ�+��L��r4��G�jhsw���{_�vq(�a/��Go,H0��R]�eZ����Ɖ�o[�x��
+&����*��c�
Z{;��9��ّ&j�Ҳ�����K�@su���>	;�z�`.V�_����tf1���r�G�V@�+���Cԫ��τˏ@i��
q�z�a���Le���C�񝭔� ���SW�M�#����Q�)���QUPa�>���Ee�޿F��B�L����G�N��yNt݋l�k/@�C�v]�jr�GK���᠌�Du����s����n �PC[cw�u��TP?���C~_3�ӆ��\�g�\n�@�c�	���	�b��N��0_i�B|G�1,1(�����<'?'����d�����`٧��`�yn�;�̠�g�sӲ��is���;\�G��4�l��ė��5v��Ӱv�b�@�E�ȳ�@o�=F����I[NYxh��(:=�^7� et�ya�z]\+�!��X�X�P4ɤ�O���^��ތ.��:��:��|�%4��M�-�fQ~�D0ऀ�ZK��
���)���|������#����U6�$�;␈��5�ރ�ƈ��$���-

�0.�S ��L��ah�l^�%uD�����;�QiC��*)�7sE~�����&�U�#����w��i�>��{�]*��:���-o���������n0�Y��o39"��x��cdM(�u-f�؄�U�*��UHN��`��˄�AzF���m"�PJ0�4;��� N�L�c��vm��T@
�����6��=&�ӬL�7�|�`⭶9&,m��9�k���Cs���0~�����H;�w�h6��s���+�2�'��U] 7NΑA�do��P��$)m�P�=�pڞ��Ф�T
0�!_0o�i���kk��ł�e~1p����i�=nNu$$�;��%X`���,cA�����'�	�<kߡ~5a�Yљ�J㾱LL��0�cr�e����m�)���~�n#��7@K�e#ǈ�>!cZ��b��v,C>Ĳ��m!m�[7s}ʹ�E{�n�>�*�~7�F�[��f��Ij��_T��H/j�t[xT���������s��@n���ܰ�-�U=�Tφ�=��瓢Q,q��]H���ad����7��R7�@�k�2���9�8#�L�a(��
+����8�o�Xڔ����qQE2���g'�x���zU���S��u��|�;E �p�_��?�Z=n�K5y"Q�l;�]U��Mfkf�i�iF�����qD���i��L�N;م ���	.���ߘ8�i<�چ��BRi�@5(�5&t�x#���\R-��Q�bћ�>U����~���U�=:{r�*��&��dX��4y��1��1p/���J�d�z=��_�KF��O\<��4N����P�J�3�XNn>���8�Hj�����Od5FNcV���i6Cg�?w�A�mp������9�=��S��� ��fҚ��l�0F�h����)���*9sK��[L��i���)K�!r�������8�M	.��^�z0Ҧr���8X1�TͽV���<��qQ�!�� >:�����%/t'�����,�{t�b�s�8�BM�����k�1Ij����d>ƭ}a]z���.ĵ�%�+Թ1���v�Y������T�_�VM|xܱ���@ԝ�E(���=)k��ZefL��5/�Y%���fpP��������l<���Q���G%ƚ?�������u8�uE�S_GeR��Seҫ�&���U\��ݵ���r�}�z^i^��&倫�m}ӗ�h�^��u�4}D�ʞ�ς�~_��.b�q	��	��t+�5����^��xV5�3
^3�һ�I�ɼT}��KU���Ch�d@�ՃMg�s��^*[�h����B5u,8� �]/X����L������օĮ��
L�o�J�O/�#p�v�����wW��i���;�͡����Eg¯]�X�ʪ� ײn�CC��,8'bn�l�ܡ�R�K� �ܚ"��1ү23�b�ʿu~	�Ef�0�i��ͥ��N��@݈#\��S�$Q~�t�v�McX�l�7�@=��8����^/��3�$Z<���;J�G�RZ���ZH� �+���d��J�ٚ[A��#L��avV�9��Z	p/sWH����1&O[Z�f�ص��	��6fj·���R�b��v`�沶�륏O�� �~��lp��B�}��Z�~s��x"N���D2�#~��JLW�	n6�/� ���HA V�xm���W1�W���`H��솛��e���}��?:qݕ'�T����2{��A�]e�y���KDx�jY9 ����7:jI�'�0����]Q3 >������r�-��8�Sʁg�}�v�vB�S�IH�F��R��ʦ�V����uGC��*������엏�1��IL�ޥ{�\�Wt�
䈏�r���ϻ�j����	�`�xȅ쌍�(
ja�^��Y�k>�:�h��p�Է·��"*�<%p7AD#��]�ycI����e8��M�1��P�E]un��>`������R(U$�@9 Is�gz��I��`��-�S���zH��Xv��CF{�e|#FLCwK��y;��mN}��yh�n��oT�jPޚK�<�9�
L��==f�k	���tPÚ����J$��A�n=v������S>2u3�[U��R��q+��t�r�6L�J����YD�c@~'p��ry�9,��Z:vJ����1r<j�����Ć�n���"�Z�$���H�c�l墀k]�g������p�r�\ݢ0�%����>n�����Υ��9~$G�F��-�D]�a�W2�Ge;Z%�8�+��g�G���z��?��&�����>��ld��>=v ��T1��vo���+qAG̊�����-��ɯ�X���)-��Gē~$%�$j�2WSA���P:q�nX�(�	q'}��5�RҨǚ���-9��y�m� �^����;۩"CW�H箊Gو�`tэO���-�m.�O#Xu<��I�f}J�@~�9K�7��Y1^�j<ٻ��F7���=}�u���-#�����J�L�X�oh�0���Zz�'Ժ�Tځ��t�[��B�J��ݒ\B�Ԅq��&�)�Pd�󅫖zl���E��p&|�ώd���	�m�<��rD
-�4� �AJ4�ks��	�#s�,�NxQu1��a{ǚ�(�郆Dn���N4*�!�i0�ޅ����V�@sa4��|,NX!{��T�3��1;�Xx�����/6E	~P��j�Z�|�--�d�;��o�b�E�8x�)��7Zt&�PN9��u�D�g���E����{��5H\r��pa��<�Ig���P'��%j����=�'��,I6>E����.>h�:FkLlS�
�t��;{��,�l(��e([4UyV���f��Q�{Ai�{�GR�</�ޱE�h a�Xծ�֛��B���+���_�&m}K��g��AVS�R����^'�`�J��~��P���e���>�d0H���7����;��z�9��m����Fd�6��0�'`��H��r���f�/��|?~i�����Jˌ��*��S������V9�/<0���9�Z1/���

���&�V��T���|�b��[����n@?����M�t��7�*��
����ՠ�&n�)I7�/,~+eH��٩(��GM�d�����-v��d���/>��6�)��n^j�LN�����{[E����	�Dc�Q�`b|���p,��i�����1�,�:��=��=e����]\&�w0�,�{�fC��)��
s{��Sb�L��b�i���i1mi�5]D��BO�M1 ���gÞ!�gL���&%4���u���iSU��O��,����y�ꃣSAٜ�
��`�i���3]6��ەl�н`�t�W�����a�Ub5r'��Z��J x������fR�a�q���>�7*�+���� �Q��,^Z�\G��,
��G��b�D,��i\*G
�K�`V�rU�����pQ�����}m#+��~
mӱ]��(�rt�9�d��y�E6/������ӁK����o���5�x=?o��|�����W�R����|_-TLB`D����R8��F�"���"�ݑ�) �Q��pfط�>�HQ�:y�/ӯ��k��E����[d�Ȟi1�R�)z�=A3٩�~���I�!�h��4z�Wv���I1R �DM�4�Lޅ�%X�}�ڴr�tHR�D��`,坔�'�A�눅8$�2�j�ў�DT�E���ܿTS%0�5En���޷����A�`{���r i@�_E��cZ)�+*��[�� ��jP ���<��u�u��R����H��v�x���/�(!�.R�7O�\s�G�?������9�?Z@P¿���v ������G5�|q�J&��U�[�&{Zu�C�R���Q`~�J���M8�:�~�	֦���6�1�"�ԝ$#��t�P��s;�a�*cYU�G��gm*��#�2h����
|4X�ٴ`��[��jc3����i��8'
1���lW|zj9����蕃f��x���4γ�ߵ�x��ĵ�pm� 1���-��Q�k?��/ؐ�E�(�w�bq�t/��}|D�ý��>����JK.>�Xʶp�:�a-�F��� ������U�5�Kp�v�n��c�d��d.�=�.����`�.��R�_�����ݸ�S�H�p��]�/x:
���T[��A��h��2� ����h�� ��ǡm�bOx*k����+އj�ﳙSL|yh|0F������aª���h'y��J�DL��0?|�%�-l��=i( �򵬶�=���6��}{��'$P�l����aTJ�9���n�m%6�&4%gV��%N�W��.OZ�ϿH��+��=�V��B����-���h��Jn�Z.��c߅��&�f�l�I�>	�� �4��h�h
B�@X\b����*�Av��G\��0tg
e�f>Z��xa�2�D����9�ؔe�C���l��𺟎�Ʉ��N#I�5�8�	(Q��ܥ�T=	�D����u�]��ڴ)�0��-[b[A��+9�О/�+0Q�#��R��ܷ�0�44�yd�y�I�"�&�"�RN���0�s�%�:��j�gҪR��>��^�:}�g.���ubHgæ�k	>,� �J]�1{-�yV�����Z� b�F������E����,�a2Q1�M�ׅջ�]uAo���i#D��]d�I��*��@
�+�cu:wF9obz��;�[�y`�:���}H�kb�
MGH�;�5��\O)��t���|+9�!*�ҽ�:T��b.5VdRܓ������ܭXh+��������B��q�H�Q��Dl�
"/ӕ�0��>>�x]��4M.�mi\��j˨�<��h\��?�VnĮ���nӎф�����^�3��S�Loca����M�v��Fc �zȠg�]}��+s\2�,�;	D!�|�ht_VkCL�d���)���.�U������1�?W5������K�haj�-���rϮ좔�VG)�XA&~܇����j�\�׽R��X�:��,HH.>��tF!�S�����`+�5l�"�I[�b!$sXz��"���ӡ��Pw��!�O?)���CYYL�协��K�l}���ϼUy�,/mv��IK��D��O;�殌d�ÑR��\3����HH�|�07�m��d8�g��l�Y3� /��1db�K[���I�$O]a4�@J�/����� q���F�|�����d�lun���$1�)�Ǉ�[��S+�,q�-uǯ�[~�B�X<`7�GxM'��V�t�6sBh�G�hW
��b�����B� �h�ح}P�Ĵ/OU��ި��� :U�0Bn�)R����VZe�"����r�;����*~���l	+�d�w����_�nc�s?��.�J��t\�pR�R�#�C�zۅ�ZAfv�.�o�K;�'���^=��&�1%�����ڒy7
wR�'��V��!�\�5��k:'ل�c����}L���Сj�C,g���iR�r5dA"(���2
@�)6 c/�u@�إ��yg���Y���M�]���Wy�G������,��_����5�¯�c�έx��8k�l� WsC!}k�/6�!zXW
d�.[�`3,����}Iw߾�a;:�` �FTD�nVxf	�t6cT�Pn��Yڶ.ˇ���������*�U�%���غ�N�A'VCU��W���d]�r��L*�4-��ov��ﶵ�ة�BCO��p�T�-�Xy#�=3q��3iJ%&"�u�pa�K��G+K��MBP�<� 葒�y��Msnv�k�.�>w�[4x�)��9��ڬ��,�,��$��癍=��g9��ʇS3�8����0��;�3�ᰃ�ptG�ROVb�D'�Yh�:����+��j����q�O�t�g۲'q�}pC�~0�'[2\�M�^��ת+�^��f���V�$4�Y��ONg�P��g�`M���<�_����h���Q\>$�f�㼁�$��}]*����:u]���'#rF��d�n��=���	W�m��:�h��Z���{i@�h=T�g_qZΞeYL;?]TZ��Y]�J<�zY��Ls����I��S���!_�:N5;�ƕ]��ܣO�s�Pv�EZX�qQ��nʁk�m4����G�U�ٙ��#y�f�\`'%�V�tV�< ,.��?;��[+
}F�RjO���z%��/�U�,�jM�]����{�ށ��I7��A�%���2���~G荗���[��J�n�g -�����䣟����A���
�P
F()fX#�+�̰o{���}|%މ.	��Ɂo�%��0�D?�s�����`��2�Y�| ;C&�}����W���5�|>3�̶j֟���ⶐ�[Z쮢v�`Dj�kNm�<��U�-�_�.؃m�D13PNl[�q:k^����髤ΚZx�]�3��V�.�Oǎ��*�,Ω�S��������W
����5u��wK>ݦsm����Й*$>�.)��`J�H�[dp���2���>f=O-՟z˙dDa|ZG�؇�2}���#N�� ��s�<�J3-{Z#6���9�"�Oa�l�grYK�_KX���ك|U7!k���Ȍv��csb�u�OU�o����8���S��c���# ��:���z8x����x��9�¿f�>TR��n�z�}Y�lW���]�VYxg�?(
�%ˤ�Km:J�f�ޏ3�7U�҄�����ԟ� ���`��@�O��$ܪ�aWt�@�n��J��/�	H��1X׫�Wje���Z���uL�7B��_��W8>��~�U?�l�s�KQv �VY�{Cnk��U%��fES�i�).���D�T���2Q��[�vF5�f���	1� �}�6��DZ3���������'5_Ǳ��=���`���/7fx͘�ȯ('�� 2&./k��}�Q���!G25q>A)�Q������-�@�g�Io�ju
)��v�a��3��@��
��Uђ�fr7����%ڇ���ꤩ��>�n������3����!IN�Цf]i}��h����E�G 'X�BV����9���w_-�f�_Kx��+Z����C������8����;S|�w�1,��XPO��\�ԑH	�vY�C
9.�B����]gUA#P�$(�x�`�g�K	�7LӒ
�����Z�ݹ�_�H�����ۤ����o�Іp������E���S?N[�dٕi���h�Rd؟�f�=#Y[���Qc踌h��KY�H
0���魎��$G��_`��+>T�z/�^�ɖh��Ƕ?	;�H|^7^������ܽLrA?���#s�'#��J
M�c���\Ŵ㧩�|.��Yq^�-:�.}�/�s˅yZ�˷���PP�~]�%�����L}�6�Qf�S�g�����0S�ȟ�.��JN
�K\��F�c7xK����r"�����˙�a�8�`l�V�Ա(ɶN�q������s��!���L<�=w��E:� ���9w�hD��Вk�?���i�����b֓<ɚ�B��*S�(~Ȍ�B��w����<��k�줾?�)Tu�#/�! n�Y3G�`䓔?Ɣ�ݰ/O}�\����"�������c�e�k}:~��Gu0�� ��s�,0Q!��TK��v��Oᑾ���]#�L�8�mEc{�e6���bzҔ���UV�acJ�s%.������՜���֢�a��2�*�`���J��@Bd�,��H���b����R�u�1*ӊ1 �w͠�r�oC��W��`�K$k\�)�<�<�.�0���ߐF�\f�&��3'�Ǜ�|G����00W
��dv"��ԧ����0N��xH���L@� �u���3el*������} }/�9!fl~�g������ʍ��8̵B��YK�@q\���е��7�5ehf�?����3"$�,�X²DԂ���Çg��=K�8�p�"l�3f$g�w���P"�k��h��L��&=-��m�{��+��+������&I��]��\OC �C/�|�H�7�֚~O*|�33�||�u�j����mVhr�.�*!�5�,��x�񥓪�ͭE�'O�D��]�8�#oh���ڟ8�6E������~"�]I~���93)��E�G@S��P�/�f�w�"8w�3��O�������М~�>��V��h6��и�Ӹz�է||�dUdS�6�����U���!xz�����hM�|�)t;ފrBao���\n��g/�Zy֢h�%�#�Y��)�FK9O�f��4�u��x*��l#��F/j�C��
�	~Bw���T���P���҄s]�'ᠼ��JL�����}p-� M#U1�	��^[�5߰]���3@P��7��=����V�z3>��?�ŗ��z��L��)���3�K���~RA�(�unsRCS����1��Yw�4V�Es���4�[�ӏ����`A�M/��Ԥ2�S������`$zϚ�k#QM�"_2��p�4�P��N�axC�e��LD�֔��*mž�Uf	�٘������~��D~RJL������g�*&�0s'v� �E��j���+����Wo��X�K�A�S��/�-��a�0�����������l���e7�f�~�Ď���.ׅ��������>����	�/�23n�3��������CSG 'mLG�@��9L��zBQRa��DmG2��{'_M>r�3�Qz�E���e���}gƬ� �_�=�����|��N?�J��2��"2����ȨO�F�}<�ˍ�I=!�w�:��u�HV2�B�n7Eն�Dn܄�>l�F�WD���R��3�r��� �k̐t}*I����K\��Ѷ:��Ȯ��5��d�����@MCV���R̍����t���W��dƎ8�rK7k�r�Axk~��[�<�'(�Eԃ+?vP��_ŧ��bN$����=�Ԍ;�����`�0�g�S��e��^��?�S�>�Hm���>���̧ �툊Bj���;p^�p��qP�X_���Y�6*0�wDTs�;��Ѳ� ��8�G�/��I~���q����v��2�����>ճ��8��I%��&��iyn˿�
ӊ:����<�=�_�j���D]�\o�M���"�(i�r�0=�q��(������,_9'J�JF�bQ-%O.̗�KU3�p
�E�;xo����B�`l�#d0aċ����F��ժ/��"�����V��ih��:eœ�8}��o�H'�+j�k�V2�$�#{~en�@�.�E�|,�?����V��_B�?B�p�{�N< �n�nw�/~т�b��8��@��/���ߋ��י힂Ñ�l-o6)I�e�G&	/VO��(�zP��H{tNXm>X���fj��p��c�����5\��=D������w�-�_�xK���EH�ǥ�_��Kny��=������ݐ��h0�8�`���~Zs0>�ۈ:��'|y�c#
��I����rki�+�.j�axTN�ع L�j�$����e�:�3k�Ț����b�#A=����u�c]�����ɩ�Fy0�W߄$b�7uc]��յ���:	��x�~�����/a��`�I_U��OԞ$�q���ˮ����#�Y�n]Z�i���._&>{P�������o��m�O�Lbf��Ē�ED�A�)<��t��
@ �o��?�X��B���^��͇��h��kAau
(�X�H$��~.k���,͛�:��o0Y(�L���]\�������sL��Q^�}��y�ލ^�J�����J�]�҄�=c^n�Xo1K��~
�iA��c���4nJ���s[��+s�z{�F:$O5BNS��G'�z6�xa�rW���9q:��� �$i�4�!�]�0���d,j�Z/��R��!�Q�XL8�0C�=�G��ۿ���
W��"�b�S6�kC�*FWޅ\[�L�~��i�Ơ;���e��AC��fJ�	g҆[�|����eG���O=��N��<G�et�vo2��p��_���H>��!#\?$lQR>���
���y�`�lö�㤜����S��u��!��3Ԥ���G]��y�N(���ȑ��hh?H�5;uc��V����P�}��.��E�̂%��,��v�Y��q�b_RϻtޗV@��Ǳ*���&:Rؼ�NE�h<�Xw��ȷ���M?������L�5U�@xI�*pVk�r�e{�����R�@��~M�x���@*JA�8^�$ia6��p`{���J����,q����S�W�$d� ���Uc������- �en����B �p�@b8���$��a�L[~{S��c6�?���`��xn!!��S�౹x���k{%���-b^��^�����[t���IREE3�'��1Zv� �j��E.ӀY��.��ʪ��������J�/suTG��	�2BF����I��c��	�t4|�Gi�eZ$�D��F!��ǝ�r��~�ɹ�dV`��g��q>87���-�\��<�C��N��~2Ӷ\=@z��;<S����R��=���`K�^ᙚ�����[���(W%GI,q6ff����os���3��x5R!�d8��:tԙ�^��$��(��ͭ�	�hlsij���Z�IͥA��s����/���� z�93��:��A�xf�|D��s��0�q�R����O�Pf�soYa[�����#;ev��,щ�t�G�ȵj�n����X�=;��8���]\"ݣ&��5����=�	���.{D� �]����L�.=�P�;�}Q�)kҖ�h�d�]�EVP��}K���e����a�:y�`_�p�S	L6R�}	�at�id���Sjt�t�L�7�|�bf��|B�˝�9U��8�0��3�y� &�y�v��6E�bn)�*����5@!h]�yDRڄ9�x}~��"�A��d�{���6�C��Po����)2�i�0q��҈ۈ��H�@���mŗJs쌭i+��l��Qj1ݗX?���[L�%��%���x�B����D�iX����O�W����kY+�Q�����ͯ�%���	�;�37ID���膳��E9�ᇂr�}�.�=���/�[-Iz�F���ʃ��vw.���L�_��Sٟ���x����3l5{�55�Q�7� ���}��LB�pT�./�E��]��p�;WK�O��U�r�6�p�/�\�M�w���g���(X���p�1^�S��OA9$��p���|��=����� Fl:/eaH� ^���P�\���e��t8Bt`{zНAZ�&��e���9��&�`�H�#ߪHhm�g|@�[�X]ZL{�L"�~��5i�����E�ڹ�w�tme�=-nB?6 CX���?��/�"��y�{b��l�!��X�A��o��}��0�	��5��Y��3�n?��w5��L|�� �h2����hɍ���(��[n) �;�)����b�DQ���7��fq��bŮk����{���1ݔ����m&�ofb�9�[��rW�V;�G(���_�}T��pX�ߢMK�e�L�J̛d���.xn1\Qj���T����gUV;ۻD�G�|�;��=���LIF>��i gN\4w8E��.�ı=�)��\���tw�o���Ѐ�7���3���f��7aJD2��'2�&�~� ������hT%Gl�]	!��m��cj�'���}?ŹJJ���n���b�~G�����f	�n>�ɍ�>�d��Po��ӿ!Eqzچ�3ln��}�d�i�r��f7刍�Dd�$M9�9�"��B��)&���>�)�p3q#��`kv3a��t,����ѽ��?~�t�f�$��V��B�;z��w"�'�YTΘ�1�����g���P��$'�:�v�R�1�'ӌ�:@��\���� ���p<�g��U����G�"i]l΃]�R����Ջ�����o5.u:c���UX�|���h���1s87��R�y�z|�-�Ъ���̜��\T�(������5�)�������a�3�9�c��A�&���D�Ƴ����-�|L��o.�m���
�d���;��?�'��
�ҿ|8���t�v���B�!s�rA�jUb��. ���ZB"j�);��8��]n��G���H��,��XY�\��
���3p�!T3���R7"����B�KQ�>�'�������xoք�_j�#��A�Q�	$�NY�	2u�������-�v�O�u��xO�Q����{+JW���!�N�'�#ɡ��F�=�b[g�@��Jq8�L���R-r�,��LW�7�QT��7��Y�f~�IV�'����5�3���2�"��j(�N.�BQs�6����Giu�I]i��3Sϟ��v�D�wa��޲��l��������]̞��VY�0��������q��[5��H����D��$oa@�<��5�)�͖A�[�'m$2��-W�31$���Ώ�o�����Y���ґ^�Cn�F��}�=Y6tN[��T���/Y3g���R~�(�h��"�� ��\ WbN�z
�:STzh�ê����z�����?[J�:i�U���M���<;�A�[�YA�ΧL���ޝo(�Q	I��V-~D�rY@%�G�x�ZTF������ >�];3�5%�uD����Z/ǳ��|���rZO������5�ӋD�d{������ɼ���1��G�>�Ԩ�2׍�A7�;4��a)=���xP�aƓ:��4�F�ˁ�V�磦�l�Ӫ�$�o5/�0,��wJ2�v��*֤�]���'\���X���Ֆ�xV��N����R��x�_�i{����ӏ����D[\@�v1��9�Ǝ�-�#A{�4_Nl����L����(�3�uI�}�4QCfoY������暊���%'���er�L�̈h��M�ġ-�O�+�K`B�����x�I �b�~SȾmAF�qO���/;Q�Z�g��<���n����{vћƘ6�u_��r��u�{m{�#�
7�Y��G����x{c{)z�Ȋz	]�`O΢������DT]m/HG���kg+D�V�;ӓo���q�j`�����}��7����SHɧ�n?.�?�1M�j^�.�S��J[x{��l4��G��_U���;C�z�`����������
����#�o_r�Ms��gT�`��8�ȳ��v,���/���C�p���M��y'��y);W�r��gU���FT�p�p�s@�zެV+�b5��e� V���$�����(|�U�T�E�7����0I����w����^����������%A��>f���5=Y��¡����$�zo���i��9B�)d�7�2�"�`X�4
�>����4 �ji��D�yO֪�6LX�a���,����t�h�
�uP�Ǖb|AI����O%vM'��ń�{J`@�Il�H���j�O���n�n���e()۞��w/�x���2��	�I_Hv�<`�"K=l��g��6��Öv��������R;�Hʡ�2�_��&�.\���~"l鎹��ŷf����6ow��>B9{��y���E"�r��L�ĕn
]�$�[�`�w����#w��]�\��m��!|o<��@Y���1����Q�N� RNA	�����nKo؀�+ ��"���b@,��A��@���oO�!\��6[�v�}��T�.�y ^b��A����!lw�?�-����A3t�m�]�������k�N�S=���W��e18�D|�g�ږ�3Q�� 啓��-`\�0%�QPuA$�Y�mx? h��Q���^���+�j* U@%'d�`׎�Q���8D�&H�$.���z�7U�ׄ�Ǒ�+�[Mݵ �NU��E���ϛ�S��B������1����U�-�Z�,5���Å����ۚ!x���澎�yĄ���l>>���甞v�=Z_!�{������3���?1v����O|"�6�R\� ���C�2P9Yx�z.�.z�&Q>�w�<�S̿�Dt�!l�_�Z��Y��h���٠��j��j�Ԉp#�6�͏P��Sx���@'?�j�o� ҕ�°���\\��/$'r�/�ٺ�c��I�9��07��	1f��� Cz���1չa&k�������=v#���T�l/����M��_���?��.�Z��p!>��)�{������w�c��
�,��b�9�K#<Є��I��$Uk�e�f T����c�`V��tN��H�1N�R�#��B F�xP�̾L���';'zj��<�5�+���G|p��ף'�2̕Iq�S	�Ō��nd<�;I�i��������L�9�[z\E8�v���[C���4���(���U�/=�}��\]5�c<ͻɅ��ܯ�K��Br�%����ǰŵv���=�WQ����O�6��Nns>��M[MtI��L"أ���ȓ�;ﴹ+ə:gu����a�ѱr=�$��It��6u�5���Ofv�!l�_H��ٺl�A�	�ֳ)�9�O��� �z���U�gp��_6�ְ�U��o�%�8�|��eHF���,:�w,8�t'��}���)[ ��51�P\��,���O��ᜭ�\.Լ hZ��y�L}�\%�ڐ�Ͳ�_KU_:��R�s8v���B�S���W�%,4 Rw@@�, VD]z��״�@�jE���}�#�Դ3�=$<^1�@C�bAs2Q�)��`����0 ֣��� ��dCt���a�`����GK��}�B��>g"��/$���6�u��a/3�L��\�x.��6s���� �Bw~�،*d�»�:��r�BY�͸"P6�]�By(A��%x]FEG_�B~����h<�m��-HO�@=~W�3*s�{����<HTh_�g��f+���yd��L��J܇��\�Px����Qͭ$�z�_�%��]�<c��7u��[2FIڻ��\?�5�.��W"�Џ���9>~�U/��v�^��Pkgy7i	N�X  ��qs:R��ھg�c�0
���� '�䶬��"�ZD8���>NۖkZ
%-]�Y6�]n�mڨ��L.�D�����A��tc��ꦗ�Z�N���1���ʯ�ʧ��V?�!E�5 �OTz��ϢB)pri���(?�9٩��ѯ�$���a��sn��YXҏ�XQE�I�N�ƾF��8�5���nī9�Fb�j����Ov������L�0S 3��sl��Ƚ>�+'��	�^o@D/����*]�����J��L	�RJ�j����p<4|�F��,g������`8���ONU�G�VS.r���m ����n����]����_m��Iw�Z$c�OpA��L�g>m�~�v�7ȍ�aT�1T��c����C������i�������*=�-��LfBeH�eIVWb��|�$<��4C�a��{iwh�o�ZIa`]�満���M�_6�md�=�4=	��0��y�q'�Q4-Ӏ��J������׉?���ր"�V���q7���|��ܢ2��J�Xm1�K?�oR�S%G]/v�"�X�Ru_���U�2�/�E��B������-�|�z� <�xeph�RW4~��L*pY�w���O-�w"&V�;C��ŵ�J9�踀Bc*�b{����c�O�}Q�0�(�'*O,��k]�IO�d^r �K,k&$��c%����)�g8���'`��`��(�i����`��e�a��W�%��E��U%9�����T�!i��k��Gr�U*��p3�H���96������ޫek���j�_,��:N.Ӂ�{}���{� C'��S�8���d��T2yS߅B^��4>V��֋��i��P�����Iܖ�	u�I\�W2�:>t$� ��Ȍ��)�1���ˑG7�d�I�t���/f�gWU:�pN��g7t��X
��z9�ⷲo��~��b�lO���Q�b1�Ԭ"�y V1�
�a.}x4&]���*sP���t�C�k�?��
�y�#w̰��>_�U�j|^,mH���7<D ��0h��Up�6r�dg�T#�(nz'�N oo[fg���ۆ'�<%cX�=AElj���^�&�.b���u�C��hQ���th�ؕ��[8��n,6�n���ԵԚSc,\靮Z0|�
Ě`���X�l���v�5�5��D����y��Q�y���y!�eB5ν�,]첻��EY7h����\m����uI����!�I�V�5k�Aq�BX_����3�ly��T��7��v�ʦB����g,>��V����&y2��q�����H7%�;.'������{l��xZ��:��K�jێ?���q�vF�S�W���֋F4�R]�?�V;���>��˟I\|'H� .B��>ؒZ����)L�*��������˕]h9�W�Ӏnt}�pVd���x�f[�ui��]8վ1��9�1�A��/��343:+	5M��P���#I
�1�v�'���p������Xϔ�$�Ar�.���}U<�`����^��7�N����Yxi�И��w���CیS�]-�LKY�|�7+�r�S�g�},=9�����l�SQ�Ax=���ɵbCi�����s,�ﳙ󻎩
��z�g[�&"%��h�)��%�McF5	��)���L��^:Xa���QJ��Ixw��U]6��Qnғ��/�QEe�g��6wds�����3�i%8z�qBU����R��30�v��-/j<3���ᾣ���svT~��ABa�"�̦#�4�q��z��|e�8�q��0k1�CAi=j���~�?����Di\�<�HK2ǥ�E-�Y���{�I-�T\~�#��1�ggc��Z���u
x�����]�[&A�~���Gu�LEu�ż�Vw�>>[��k�	ķ^a����	���`��5�wő���t�Aމ���]ϩ�k�!���~�I��ɒM���"C�MB"��l����������3龻��
Z2Zz�e���1=���x���\@��Ř�,!�u?��)uO&�\i��P�C͒$��x^/�D�2O�F]���?�����t���sY����i	���<�vt�n�:�L嘾���h�����X9���۔bw���a��Ұ5�`�Mx+��M6��mW���UHDMbV�d)�l���G �NE��
�ȃ64s���A|��-2	����Ϲ��?;W��R"�(�_�P�:o�IM����D��:��od�C�<@���#h��%�L�U�Y!�9�f�ɒ��:�R�7�3� ��ި��f������� ,}[ޯcb��=hצZY�8�ZpL�̸��&-�����3{y�<�n5keu�G�4�/{��^/e�|�c@Z@e�_䭇3A�3�u��	��|)��O�����9�%�싩Сg�H'fZ�fw�DVu1 ��Rw�<N��v���c��G6�h3���
3�(8��U�?��t{�+6�~!��:���������O��H�}���'�?Nw�nP�ɘ�k�?�`�`�aT��ލ�Vv7�r��߁,�a��%�U��g�u���Ҋ��8��Ⱦ��U20!�>ph�K�Բ�P���r^��=@8����޳����s�2
�n�S���Y[�G���_�|*���4�|��b�K$��)�iI<��U���%�W��\�#N�I�\'~7]:g���b�%�V;io�1L��S��~�����"��d����!� `,�-��T¤ձ�Ys\�����-��B,��<�ZZ�B�[��}���5ٽ?mlv�:
��D�>x�X���4ry���Ǻ���{��
̚"��n�7n�o�X~k"���{�).�I�6I�	�r$x���ƫ���;'����էh��'M�;��z勎=9�����~C�o��jXL*%@�(�%��,)�w3�����i�o*�`7�qca����6�D d%�x�x*�q�v��ݔ�ƽ���m�s2dC��:~�(�=��M��2����
f�_|3C�X.~D��2\L��s�r
���l��c�������ɐKSMYc����*�vc��&�f3��j����E��ެ�����?$�.K�6��wjm��]��s��o�� �{�Z�1���9_��7���w
���N�rh[7*�?F5J~mP:�ALRs�7F����*�EttK�+�K����xw�_���oyh�1v�&,�v��}������3�hO��C# *�{#EXQ�	D�����&�P�t���+1U���|~��L�ui�T3Dϒ5R�;f��Ϧ�l� 8f�ś��ϑ{*)7Dam��ق���7���k��Q��c�j=	��k4�i<��2�/�m�S�?��ػ-���Lg�Y��m���L����Jy M[O:������N]5�+�VG�JӼ!O����*)% j�����y!q����Շ�m@��[`�Ib��$�ŋ�X�d��q�غIR~u�)ʌv�
R��uk,�[6F��&L1�����^W��5Þ�y���N����F�W��J��#���B.x�"�d-�Z7L���U�r=�9e,d�Pd�%�d0�a�i���<syS���!�[���_�y�����?�f�d����!�׬̈P���3|��7 ��P72�4i-^�̽&�/��D�dXJfab���_7��pB̩([l.�'�U:�H����:�&�Q�����'fXt>V-��GF��t���n��靲?���1����%v��6絫q(���3���q*��kۮA�?��:���cމc��9vׯb\�>�@�Nk�`�;������n\�����d����ϔm$�[�3���:������14�6A�����<�$�<����(�9t�8t�un��wXTS�uH�){��U���1zh�`Ԝ��H��d`�t�CA���a����f-�94d�j"���.�U��S��?9��U�O�L��i=���M��V��t'�)e)��
M!����0.o%)|^?�������.;p)O;pr���K�{���xy�ch�g��n��S �j1��c�"�l�`7�o��s�����_G��9�V��,͖+GR�t�À�xڷ���^�C�G�{W2�a���$�p�-� @��óό�i�v���R'�M��w]�	r�H����u��u舴�9�0Kj�W��z��Ẅ�d�q�9N�3f��BRS�ޡ�ioW�]ŗ�����)�w�]Z��ULd�J���`̕l�g��Pܤ����3�}_v硐�s��&}���WLY*
��<|�� �K=�L��us��|�?�I�]kh���T�I�P��oP��;!7��8��r�F���̪��m.�TE.��C��O�" 9��������͊���"_C@��ġ�u�pv�'D�V[Sav��Z��8O�I��Uj��0}�Ϛ?p-���Q��Α*e�9y#����W���8�qsT^�nB��O�`$;��t�����Zj!�x���Շ߫�	�m9��Ɔ��+S�S�4�'��BvE�S&\����*7W��������&�fDdܣ��:G~@a2��N��{@&�W�<@{�m08�tX��H���O��/�7�;�zUe����#y��oV�'GO_7�I����h�F̌�K�ID��q3�8<A���<�{)zÇ2"XEɳ�Ξ,M�#�}t>P�9�ܾ���CQx��}4zz36�T�}�3T��V֮�"S����r���N���eo]�>غ��E b���Ø��<���e�TRM\�6߻~�1��s��#��wLsִn��<�V�����)u{�^�/SC~��z,7�J��O.���CA�В�u>d��;�e���+Ɓ�}�RN'�[�tk)�!�h���"�>	-�{u�P�����j�����$	6\9�E��qO�σ��N�Eeu���=!;U���ԛ�,��{s���9*���l]��"��2Y`�����@2x:l�2�ԗ`!�g��u�"��m$9ҫM��If.�3��Q�3��ŋ�:bt���V��?�$f��T�������2�~8�����?�q&c�6�ߖ���JϖK�x�^��)+�@pa>�Mπ`�N(7��,�o�p`]0~�8��}[��}��`S���%E�8t��̋h��N�����w~0=?����Kԝ�-���������1E(��e���P�c�y9tƅ1��[iD$�{d�oE�0s�y�����wv���ژ��~t��uU�_$�zn�,�������P��e�{ba���{ה�J��sZx���@��{�_�Z�����|p��sۢ����ߓ+E[� ����������.Pk��P4/r��zN�!��~ۗ�O�A�붙='ǣ[�����b��tѳ�s�o����`7�P�AԶ�z���N��*��^�P	�U�2�TG��B�&CU�V:?ڡH�.�A ��`	х�)pO���~�G����6SEo*�])������ļJg*#K��W��å5.X����4��|�-��~���[�ʮ��E��\g�v��C{����<+��F8H��Ѱw���Z�+�&z#ĝ�c��j��o�'�e�<�n��v*nP��kԗBLH��y�H+�e7\B��a#�s@���B��AV�<I��Ah��T$�ԁ65<�T5Jq�zK��>ž�{v#���u��)zQ��D�srfP�$����F
�z&���k P������^k6�w�X��>*�၃BPP>ډ2�mTz�����+�<�Z5,�Q�)�H��t�+S�n��<_Z���5�)��&��#�г��JϓJ4C�=�4��n��*�v��ֽR���H_�|K8.b��v8��x����lh5\ӣ������{h�+�Y�Ӟ�ȴ�琐�8%1c�q���Lg�pS�_��)����KY��~#�"��%�}8��	-Y_���3�S���^��H{y/�&�YԒ������C���z��I�q����Ǜ�һX28[����[��1߈����*�W�0�I�U������v��^"AJ� LF��P��.hi��0��Vq��:?�ֶ��%:��2���ش`#�� �T��F�55��)&�����H1g����#]V�;�ZXv1���gU9�+���H~�!jU���5�{f�����wrj�s�M�+tq�hWP����]�Ï�������_v�S�S�;���I��]zƷkE�{�fFuh�Wɟ�g/�$u���Z%�^cj������8گC��*���8����5)��$�C�~�:�\�@��g�ֵ2n�9<� ���>%a�]��gEy�����,�|�O��+� ����c��<���i�pR	� 
W�f�&V\��=r$-��T��y.���k�<U��ȋj_�Z���B�:&Պq�+���.�4ު" m�'�a�腎	#��FF�Ol�(��s���(0#�"b<6AE�)�/�FZ;z䎅�R΂� S�q���s���C2�V�tE���'N�t��uB�������>�[{2��hWR�6΃b�A`+����_?���p��!U!\��j�ko�D�Xc��fui��hWcft��26$~�8���4֗��g
a1@ԇ�b�\�A�O��q� R6�����5�g��[��awE�q�����c�cQ+%x���4�`��3q�0/�����oZ�?y�R����"��K��D�loVo�������������x�^cIB��1�e�y�!���$�-�M� ��\�U%���#�UF��	���A �h�7�3)��({�	:h��q�y����NB.�M�"��31���ʿ[؞,ݚ���q����@S��%�:�n` hH���GA�j��K�`Z�cvl��ǈ�WL8��&�*��HÑ~Z��}�Y����NG���\�E��c"c˕ZA��Dwi92�Ziz$�Z�Mr-۬i����=QZ�,4?�� ���tj��h}|L��M��6��.��mzГz�#if��I��'T"
8S+��pi=7Kc�˖D��X$T�n MF2��1��YZ���P`���Iw�g���E�C�܅�=���8e��}]
.>HH�4�dv�,�"=�� ��K�3��J��%�'im)�^ż� /�;LeB�5�64ҨI�_�R�n�W#��J6�<�d	ǉ�;�V��� ��U�¸�ȉ��t8��]��_�C�k(���Bt�}��X�4F6.�ʡQ�h*S��^o�!�]a�%2��٠1ט#Zo��s����ݺNj{����}���󑷷��"�1��D�nyQд[l��l�~�Ԏu�?%U	�nC���(�|�;T@�S�c���xk��s�t��9q=�h�j��]�
!x�#�OVp�4Y�AS��ܴZ�2�������i�&�tD�ބ��K�y�;~L>T�t멀�T���GyT��$�$]\��bޏ^9�( 2�E�`�a��`�njJ��_�,�Nc�P�ȷ�L�|r"	��O��xR�\I���h�}A��&�M	su��kݾ������`�M�rn8��R~�4(o�]��0�@JF2co���=7�N��%~�F{���N~��E��O�z˚FC��\l>��tTį�m�5Xo	k�5���Sk�s*��v2��լ�GG�	�\M���\�k������Wc���K*^�ٔ̔>v�:#�U�[''q �K5����`�X	f,oaTu��@2[�^㔨z�~6o����n�3�Bܑ)fٷ:_�DC+�� d�'#o�R��s<�^3�יyu���/?���_w�v6w�=j�I1�ɞN,�h���stJ\wг�<���$U*�:Gן�jg|%C�O^�y����q(�·���{ŭ�a�ĶW&�-k�A`�xD)(+G�ǿ�[CY{CV�^|����LD��i
ڞ%�:5���cQ�+`zl���l��i`���ޕV���8�� �&KJ��c�AR�z,I*b"����w����%����ňH�B��ϖ�@�V>2���vl٤��*X��
���~��z^��X�:d �Ez�M��b���:٠UanH��:�REy���x�$}6K�o�[O�N<�Z8�C�*��4��L��X<F�p{����Ib�tByl�b#����*���%A�c1�~qQ�.�͎�X��m�?�J��PO�y��ZWٓ�t�`��J��a������f�:���+_qt�!��l�~�_u�7|��	���貏���*�2�NqLu1e>;�r���+�\Tpەy�}�8�u��w��~R<@�}
D�������7h�~ѭ���&~?@O�7���n��"ᆓb�W���@$��;�C����2;Fau�g�I�.��0´�G����A0�}�gr3��h�Эx��� |ɎX����M�T[A墷���W0s*1%C�TP|.s��Ó�:�C�|�B���l�.%���YY�;�ZT�w��/�YS��Bxܙ���yW����pզ�J��C�u!C�lV�*MÙZ�д ���N��(@! � ��E��J�g�"Z�uI3�)*��4ĉT�s����4G启d��aq�	^�2J�0�����V=o��[���F�r�����g0RWTqМ��p��]pgl���Cý��ӟ7�5T��l��|�k"�i�
rp�]����%N�����8�C�ޓ��i�E�h�N#"Qc�Pe�05n��~A1*"<���o��q��qp�3�����Yw5�R�y�KP�!E��L�	-[�"�����h���rd �3*��Jt��9%����i�O�F�'t��+�qx,>N�+VZ߭摓�םVr�([��V���>��#@�v���f�9J������=���M�\�ߒ���:�S��� �Xt��HP�5)��<�[W���2��P�׃VT~}����Ν��Y��X#���)t1�Foh*`�=k?(��l���D$�E�Q�E˰��oݟ�㌽�ٺ-�� Q�����d���w�J�H^�M.N$Jw�-�y����%�g�d��\��K&ǫWA�U�7v��@�BFe׎�ϭ�K���H��ڤ}K�����^1LA�ID�� �I8e�(h�v�1��g��������l��Q�|_��[�0�>��Vj��+�.|����R4��S��Bjܪ�}#9>S�otnR�iĿ	��v;�͔�y%�'+����F ��<�e�<�����v�Q~�*��� ����r-�����#[�D�1}ͯ�O��w���FP)�{n����3_��k�^w�O���Qa�Gu�N��qDU�S�Ui溅5}��QJ!=�����Dv�<é�8�'�����`�[o�D�n�3�M@$����~ ��ȍ��F��|S�J��������
�(c���@r>�����a+�*e��p�l�{��$
����IF��h�h e���֛���J���f��K)�	`X�Ŀ�#�U5K�����Q�bA�,j�EÓ$�+:w�T?����{_�0N�ZQ�{��|����^������Yv<�0�� ��#G����k%�Q��b����k�Ȭ�p=�{��MD�և+O�De���6�,���a+/ܒVU(,y�o��r�kQ⼎}r.c�1 Y�w��wX.~��KHy��hʱz����t
y0���s���M=��ʟT*K;���a�:�3l`ѷ4�T_^����OH1���i�p�$���cBa
v$�e,���ЍLLߧ�֜5
iL��sK�H��_0�>`6"2���0�����c7��!6�O@B't�!��ԂQ�X]��)�Z�[��r�͘�@�	�l�J�X�Њ��Ҵ���-_��E�{)�}b��Vd�U!�۞��bB ^v���&��cUzQ�9:�=����!��W�������-��&��pGa�g��*�t|G�
h1��$7�qN/��Tn���Mc?V!�F�>iXT�I�RK��WY�D���^�Q�nF7_+8l.Cʱ.)�[��^4��R�}#-p(Ev�e���%�7����dc�FK��-�@5s(?��fn��Vd�:6k���I�D��"�� �s U9��9Q]b3sɯ�E�i��Gh�9?�{2T�7:pG�%���܎�(î"���yU=�w�����Ny��P�沫l�iˀ4��Їߟ�pͷ���X��о������2��MbG0�-|%��&��Ե���~�r��o���5�Ɏ�ӧpU>��"� wH֜���HY9YT ���o�]m��~�L������ʮ��7݃�J(�z�F@����H�A)e�M2��l���縝�(�����"c5h�`��]׻��fÕ)a�bZ��k�w�:U�ǀ����$�c����AA���*�CT� �$wۍ9����|�֗���*��*���υ-MѤA1�}��Lo�����z]��Sqb7a� �d��	��u���u$m#jD�މGL�k���v�<�e|���U�	�r�;�F�֧���1c�6:���Ɍ�[��y��Qʡ��1��۠��Ct�z�$����m�|�\P�ᑴ+^5��(����Y-�A��{o�:<U+U�t���V88� tamL�h�߶�(>x���o��H:B����V�b��ӕ����뤦#��,#���58^^*���Yj��������թ����|���-�V#!����v�t�\��ˉaPj��#7 �O�q�ьD�&��$t�=��kё�;���7���))���Gôm�[xF_��b�X�(�cM����6%6���M�w�W����2iN`�
C��B�ZJ��W�f���1߿���,���F��'�(�W|v��y��z\��ɤ��lŰ��N��)g`�^w�h�!.�	�@�����ȭ4Vf���Hq��[+é�u[��ۿ��r�\U�6j #���1���n>�l�|�U�1�t��}S}h����W n�b��i�2���g��Y����K1�✘�����ٜ��!���q�$�9�+�����Ȋ�GT؂�a��J^���=���3��}śv����T%��a����6K}�Ҩ�Ų~rLem��z�V���:&.�� ��[�6��t�N⼴���m�K[�b^�S6kppoT�g���kdw��4f+]p�X�A��}���w��@f�\U۳ e��q����,�i�X���i� ��e�}<d#�!mpׯ�J���^L���ū;x���o��Z��˸�l�<odPY�7rO�$�����7�x���P�r�yo��X���`�T�p�� $�� o=�n��2�2�n|;�"!aW��倂��t��%��U�KQv�F�Ƹ�����F��S8dE ���S@�}3��	{d�^�V��;i[�ga�-a��ҳ�R���B!���n��R�n75��S����̵J���m�z�.�ʊ�&���H��4�j<|+�$��v��k�[c�d��<Z'�T?z����ڕ��b��<=ڋ�1[�:� S���GC9��q�V��Y��{`=Wƕ�)N�tZ��}p�̖$��L���;W���F<}k)�)�u���H��*̹0�iEST�p�.�]X��v���؇C��m��"�x������F@��b���b%��{�1r��8�lt�����d��+>�L�f��S�`�Z2��z3آѹ�K���'�x���]LUo�ir��r5���2��`� ��J�)�Z,
�Dq���^���
���>�BN��,^�Ug�����x��3P�(��Xs�������dRy_7����nB��a:��)�jN�=��w�ٟ!���I�,U�p�y�}[?�Z����áiz����@��������6<� �G�gE�!��(�}SS1��F� v�4u�ﱙ���X�&!�gb�p *��Ѣ��ń�
�)9qo�A�d�EI�YNP�C�<�;D�v� �?"9~��d�5��Kq��Y͏�"ۏm$N!4����u8��)6�����3������s��ĺ�٣����61n鏺�Щ\t��h�ᥢp�8 �x;k