��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd��e�A���j��I�뺲z_��T]K�2��lّ��LsVv��ڴ�!>��>���į��e��G~��(����
��*D�"���y/9����̉1��1��s*4���ߌ��� ��=��_BO[N��CO�K�,����b9{�/!d)+c�uG#2�ȉ;>���@E�fEK�D� ���p<"���,NZ'i�C聙�F�FD���?��i���@���6rlN����xFwHw�U��~�<"99�T�����C�J	�@����E!���2cp#i,���e2��Z�/��Gp�C:���.�W�H(_��*�s�
�柙F=���a/K���[�I�1��-|��x�dGmL�K>��B;�/�	g�l�,7�YFk<W�	Q���2���e������:��@�v	GXe����L�L��_���@(��)�\=�����1�X��������U;e���	kA���&��5�$�6f�yK�$O�̀3��gPE������ꅠ����ɥ��w�cvX;�G+��Y�iH1�H�U��&J�w�S��,ۋ�_v6ۦ���V@y�W��uѱ��񶇱d��Đ�P��?0a��<o!���椿3[y5i�]��[�lQho�R5�dMv� .b�mW�ͱ^!aJ�-V~NpL�Q���"��'"MDT����Oq���9���N�T���o��12��~��� ̀����R���{|tnI�Tj
jpE;���<Y{�(;�А���Lh&� ���?C_I�G��ˎ_�JE@i��@9�����:5H��;�&^l�yK�T�m����a`c��C��go&Ay�m�my�I{资����>7�b�h�P����M�6�g��63V���r6v�݉��V�'J���=�f9,��d5�a�<���}�1��q��ɤ�G~h�"k�Y=���K��(��%v�TGK#�HV�:��,쒕e����Vh1GSs�%L:���wM��+Z�[�����7EK#�Bm7 �ź7d��*O���4����r��R@9/�n̜�_g�yo
3��n"�2�]@��P���]E���ȃ
��b��y��kS����}1�w\.9�lq�p
�5�6�Kg�0 7���q������UF��B��Qa����	�,��:e@:j*��JL;X���?���χ��_���0�Y�q�'���e�W����� �����O��iC �����q��tiǊK�dm����~.a�M==�']�˺Q1���,^�$w��*�F �d��uY��l�]��p�v��s��
6a�� )����0,D�͊��qў�Z�d	+�O�0�%Ü�E�ݽ8L���@v�;�a�i�Vz��Z��D\���C���b��Q[{m�	��?Dh�6�c��
9�gQ\��5��6g�����n��/�<MU!��	�L/��T���x��R7�Wh�q
�\={�,�*wN�̮
��n݉ݘ�訊�Wf�_�Z7	�n��P�'{/�f^�]�$1K����|�������B2�(�V
r�7G���׊�
�.,��2�������A�:�ԯ�0�tE���<�rBݑ��D�hķ/��X�M���Nz�c�|�t_~������v��Or;�����ֈ_x�?��,�'�y@F��S�L<��S"��^��TCi��>�C�C����Sg%�?�K�o>9�P�loJJ����̜Z��������l�H��n���9IZ����� �!W��4<w���7p�D]喩*u��=';o��Q��vnN�A����㢋�)�:OԂ��_n�)��.qd$Q3s������"�8L�|�z9�-���=��h���+w�m���y�>׶��|iɏ$@��y�h��z�n�E���2a��
3�l|�?˚���G�Bx�桕3Z�05#�Ѷ`t ���υ"�w%��/L�l-@xJ;�>�A��~[W�%n������s���I+�(`]��4��Uc�ׁ5n��P�<��C�DBx+w:w\h=�(����K^Q�&`x��1��M��L_����&T��g�"���2R�Me�t���z���;ٽ�4��,s~�]¤3 I.(S�0��5�������b3!�.�X~c�1��׊�H�n>�Q ���Ҿ t�I|�O�!��iw�t�C�����T
UM�C�w;ʣ�֔�|��G��*�5�hf�V�o�B��(W����+��3|�IH;%+�~��C�p�=$�ʩ�M�fQ���1	1��ubN!�e�K�ci�G�[�zn�U����4����:Ǒ�k�J�B4"8U)�DB,,\�VU��GY��a�2����%i ���E�����L��Nj�ؤ��MGAy+I�=�4����T��F�᫨�#�I&��B�#L��*��Y�>'� ���>�KDR�]�5����i�����$p(�}�7;��E�Wt{��c�VI���qY��'�}�J:\��^�}<�>o����[g'6����R�qV��u�"B��S	������QRp�����@p=yRyS��l�1��Z��[Y�	�cW�8��-z���S�9��tF��D���G���)��G�񇛭�S.��d��y�k2�Z�n�����H3t���/IOǼ�H��>�ѵ�Z���ɔV»�=�uYX���n���2]��œT���x Y'�m��\qkz���9N�y���(�E��2��u���#�!�:>y튉ܤ�b܀�:�Ko._ƨ�j�.ʬ_�ڪ�6�g�-l�:;l���]x�)�h�`�pQ��|���#�PX�&:_U�����	��5��"d�<B���?O� �-�����9�]c��h�] 9I�@�� |n��K��+����X>[ɝ��+T �F�5�s���7@2���}lQk�y����zh�EW̄�`��^���'y���ʧY��-��~[��nA/��ܔu���U�ө�R��hX��b��a&��5_M���9���/\��Zl<�]�x=��tP��h
=\l��0�fB�u6	'=�!��jߝN$c�������irs�,�k��2�^,hf7#��1_�0Jõ����MZ�>�rsG�ؿD���O%q�*R?V���^��Q��*���(Q{	ML� �n��cİ.>k�,}Pt���,\`m�'F�А�#
�f�;�ȸ�l�w;}�A�Ц�����7
��~L9�k�ѕY �Ww�S�	�`.��R<D����8`I��܁󠮇h'|
9���(3t#�_S���|߿��o�>J�\�=,��&q���O���D�t��EP0���`)�|����/��aS=�oe�9;z܃��ф��}�ֈ_��?v�9`��Q^C|�4o�y°���ˋmnI��\[�q�	3�[- vA6n�3M]ii���'g�Zv\@Y������1���/�� f.=�Cta^����8c���N�����P��ũ�M��m��G�� F�g�&۹�ֽ�S�?v�H{y���݁��X�����g�4L
����/�Q���>�N�J-#di��G�x���5X8E����!��r�c�u0[���E�_�0XS�2u�w����)3	��ǟ@��ڤ�,LN�j�r��ß���{������8}u����$T�1�zf��<�����a%�����&��"�=�f�2�>�2Dp���Sey��M��v������]SY�=��҂�Hz�[7����c?����@���72��'A�g_/�	�n�l׊���tV�IjP;d%���{j�lG��иLX������J�8����>/�}ϥ2|.����>p����XQ��ڠ�,Yኇmh˛د��'1�����#���
��j@Nz�0ν�S���?���Q�A�E���U^xT�Onq�/�t���	��3 �rY�y�5ƶ$0�8~��5a��Q��$����i(��Oۜ�4M�p��ɚ�{���^�fH![t��,4�'t��ɡ�O;s�T��d9�"��ǇvK��i��{�e��Ź��XFDg���Em8���4��+����(R����ɠ:Z�`LT���Ұ?������E�|�
�<*ǀq����s���]�\/�(�a$�}��2��\���a[3��ă���1��
Ȧ#S�I�c��(��@�c��UܠBF��_C�<8>z�♖xW�׽e�|�h6�c/���mC���9���l.���WITЍ-T��ʌ�0��0���7� ��H�Y�
�;����<�0�YF[Y���|���j�h1�4�����$�t�Sm!������c{��'MFv��r�~��q�����s�t`A�:
<ӑ/Z�9_�����3+K L���S����CVn4k��r�ߴ�M!��Z��x�i"��Z�-����X4��7D���J�p�n�z" �#�V#��r�X�\h��t��ϲkJ��&��(~t�j��?���A�����[�/Sk��0б�%�C����2ͼ�)�q����]���+�������tSB@L�5-5�W�`=k���z(k���{�Td����u͝�ϖ��*An�Ô�*!�zt�y"}un���{���4��5�ri�6�j�Z@&�ˮ�_"Қ~@K�?��̆�דlY�\������/*���^� �]&�9섽���F]�TV���ŋ�@z^Jīښ����WW�0���?���6�7
�*����G,��ңW���]�w ���f��'`�6<7�N����s���J^�D��,���G�ap>�o���'>��RF#����Iq����e����{��y����+QH��tz�1ʔZson*<�A���ا?����6"9;�˃���O�!4����M��[W�n��l%���s�*&׾mZ���{��i��b�]-�\�����;��Bs
������eIX�W=�?��kyc:��16 �{,\�	t^B�X��H
"�;L��}ř|�k�(�#gazO�(~�4���B�y�@
˰h���z'%����ڰ��}�Y�qu���� ˎ '�Yk�+�/j̀�t ��zV��}䚼��nz��.fx��Ht!����K�r�M�%�_��")v�5ۈ�{���#	��U�D6����=��H^X�?�T������SP֋c�)�:��w]�v��s�Ta��VO���VZ�m��Sf�d,eQ�8E��'�{�l�,aѮ�W?M����F�ߚ	���
��U�?gB�� �?�-ҳ<*�F�����G蛺=�e�^n��/#^0�[rQ%��?u'$�cW)���6jq>�GT�`�$)}~�H��Q~�CL��vx�1��x{��S�����'g��|��d(��<�|ib�[C�H�5���.�*���U�&��[ P�ӞY4>����e���A����%�u�Ӕ�9Zg���z@����7����"�rլ��},D.��K��O��on �=:��Ēy�छ�����g��=�u�
U�u-q���dT��� V]zv1��G�Y&�7�8�~��%�����KD�����e�i�f�����@L^����[Կ�ۀ���_���o���vR�b�a�Pf�>���&�NF��l|_�}��/}
��3?��Ie�7����#__	=�8������.�Ĵ�>�*xj�v�[���Uj�I��~���SJ�;�u��v�M���N�6_ �+� �%3��XZ�X�H�kP߁��N�m]��j�a�&����v��5!���y�1�+�����qyCv��=1�u�\�*����?��j�봏 GEZ)pl#�`W�ץ�IM���e�3c�V��H�&�t�6�T+=���b�=�U�TU�S�D1���v'OWóm��9/��x��R�7��Pu����'RT$uR�w��8���{�;�z���Ŕ y�m��8�]�>���DN�!���I�I\P�B|hz"�`�����H��:���Y�w=���`�P������:�XT��s9�ϔЂNGp(q�o�-g�W�X�3-��8_�8�7Ύ>Ex��!��[�h�W�2/��.p�.X��r�)�enG��L���h�WP��9��_a{�D4���S{k�T2�UG�H�\�x��F+�*���������ҟؘ�%��W[�|.��
R�>|�]z �����t-���&���G��L@2��?O!���5� �:��Kڴ�S&�����ƹ��L���C�#�-m���
{����x��QGr�+p�1�č�����C�c�ݝ}X��Z�o��TV
�ތQ�m�]�qMF�Rpd��6=s9�4��T ��l�x�\\���e�ý�7���� �[:��C68=�`�e��HqҀ�/�5 �If�;�KbD+�z'��H�7b��[g�������z����PPx�j~���x��+՝��m*��� @��q� mm
�8��ߜx*n�u�{�0������,t(6����
T�5�a���C����q��+4Y��> ��ʥ�/�{�OR��Z\�=b��9ᰇ�$�Dw��ړ� X�X�X��.?�GQ��}録%�>��Xj�������`�7Vv�q~��j�����;M�Ԉ��������	[%��I�`�xjb�!�Z%jE�:J�^=N��Dj;�>@ W��-�cm.*���` �7�T��dM�DU��j�B�YmM�'�~}\�OJ�V}�j�IZ,��h`�n����j>~j��Hc;BIl^xϦP{��O׋[2䛞�|(r�X�SI%=�����H/�Öm��:�H�-���c�}c��g����fKpA��&��T��D�蹴��N��|�k���¹$�Zq�,���j.�z�y���a���`4�����w<lOĘ{�YD�Q�j����ʺ�Y�2���S<O���.��ܡ��Ϡ�-��}� ���²͓$�9=w��G}�$� �ƥ���W��a�o�Mv�լ�Z����|����%����ͽ��k{�w�o}>�㼡jsFsP���'k�&T�IF����p�kg '�&~�(R}"���1�g͑U1s��?]N3 ����kK��y�#�H���x�c��^$-|Ae��N\6�ް!������/SE���&�Y��cᐅ�5�@m ��a�i��:����[�u?ڡBUb�2�?�Rk������'M-!�kI�jؚ�T^� �a�1C����_�0���
������x"γ���ݙ�����j�Hv ��,�9͊K��s��������\�#��!Έ�������c�<��wb�����*�>,��8n_��ON|Ɛ��yMm'��j=�NX���ӵv�L!�Τ��7����y�ҡ� l��ѭ��C�/r48=�`�!�*�q5##���L'mp͂��ۇw���A���hc�F!^��q����g_SjX
Z5 �]|�Q�s�	 h]qW����yL�6��dn�F.Ay$�7�[oU���i�+�On�����p���!�������I �xi�9�!���ܬ"au��7$^����;�h��g�J)� �ۏB�N���fG�	ނ�l<{����fVX����Y{~_�7q�1�Z�Y)�t�t�K�i�M��:M���C���j�9�:�A�7F��M��rʷ<+p����y�_�?��Oo^6�Jt�X>es?���Pr;��6�8m�V������IY�E{4�DL�eV(��? $k#��uP��$�؝�k�^(=�̓£]X�x�0ʦ� F�6�h��Sz�X���h#t��tq��I�C�����O�,-E�B�I���d�B(�T�|\�`�iWv�SN������b���^V������(%B[�h���%����THx��x��N�qG5x��VF��`�hMu8�e��$J����u��8*UX�~է,y�r�eFu�M0�>�Mi%I���-�-\`������)���/�FK�:9_��)��kM�$"!I��źIFCh_� "��A➺�.!f4jF��;�n����z�ɩ��mmR6ɒ�T���o3_ķ<Yimװ�^�](;��Z�&ɯd�9��{��	�S�Eu���S�Q���PR�#Q:�ߔ�jf�p����(��
,bW����JkY��`�*<�i���\E�õlOg_�}��8V�/��Y������
�X�f^�<'&��ԛr Gr�UX%VaIy��&����H�ewk˄!I���#F��^���t���Oo��ye���������'�'tJcdw}p�:�^O�YJ�ɔK⊥t���d��9���t��K������>��ΝQ���}�eu�2x�PZE��i�*����_�_��-�T&1> ��#� ��G2�2ڄ�����>&���kTo�*�:)b�9���{�NJ���� ,��(o�y�e�%ň&�̸)DĵΏ!�!V6q�\�f����N2Xvd�M�|[�u�3��-����Q�h�	�\��� Q��Ù��Ogv+�������rg���LD�<Z>�x�b�Z5��V4�jE[����Zi�jU�ӥ�cB���%<�������]�Ka���!Ү�Cd�їR� �".WیB�i��+O����#��gAm$�T x���Q}��Te_
�/G�ewA1�0|���̪� M%X�����p�=_'O��O���''�g��#fDlg�̳�,��>̰�O��d����+s7�zVK
�o�a
x�I��m���U�11��xl�����	�QV��<3���Qo��T@Dfbx��=�����FN��U��_���C� �g$/��������q�v|����h����*�Fs�SJ��G�d�
!��K�?T#�P�iD/Jܲͥ�$��������+�ǵޯ@Ӈ��퍑�|n�S���