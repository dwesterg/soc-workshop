��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ���<�Y���9~��z�;.u�Iw�݅C`��w��Ԗo��1.��8S����VM�4Y��M!��0���4~�V�zr����J��x1M:G[��dL
��s��q��cV���ˁ|��F%���r�m���t��J� طd��.�'r�k� ��V>��'���:�� ڸ��R��A�G〝���V�b2<R�����4���E�"_^��ʄ{zKn�m�V2_�$�P�c��F*�8P���c#�?��� &.?��X���巺��n)o#��<a��q��ɖF����M0[1F�����㹇�&�����/���5�}$�}0aA��Cz,�3�w i�j�y�E|_��`���}2��aQ��
�1��
�(;�r�.+�Z]��^��(`�v��� <c�g&�sEީp�߈N���ա�P�B�k(�׮!��Vr��Ü_O[u-/E�![��0;�Rt_K���,����#�Z&d�"ʔ�������v9<f�w�93���*��&>��E���e[i+c�S�^'����J�IH<���$6=����̷\vB��,Cy(���	�!G"�+|�jie	�Z�˹���Ԑ�Rmc&٨>y�v��d�Ǻ�^;�<g�LbH��SA�V����$����+U����[�yg9�X%�'��Tŋ�ҁ�����[�E��y��$��+}���\�:�.4 ��\'x��U��}��ג�gb;�`U1�VK�/T4��ڜa#�J�)�������sXpQoߊl9o��:�*�fկ�-u/��&r�EG7�
ie`Ѹp�d(�lJJ���L�TbO,�wU ��[[5�T�~B����P9٬�Ł�=hѓ��Ht��lE�<^�ߠF� �unӪ6���6�9,ذ�^%I٩��b�z�\t��{Kr�cI8�c֑�� D^�ۮ�16x%�n䨚m��V�AH�z�8t��Iy����V
��@�W*��mE��؀�uTgL(J�S��Ħ���t5c�{(~�Yk���pc~�A��F��O�c��Wo�l7�:�;��M�t*ˊ_�-�19/t�y�rU!g��{M�i�W�,K��I�QTN�Z� Eo"�cVL럁'���2�nDUH\R󀥒���v��;v4�8��g��vj%{�����>P��;�8D\U�i� �6Gn�)�?/���L^U���*�b�R����^��!3���y�3ncTx��ȩC�ѹ�X��3ȃ����,v��/�#���"���2Wu���dg:�"<���.hX�Z���a洞e����uS�' �{�:Kki��w�Ů��z���wl��k���4�D�H�W� �8X$1��
e�WK�8���a�,l�L,����p�%/�T\���xP�${�f:}�Q@"��!�+�b�Yg���}�Ǥ�?F�XN�	����?�pry�h>�-�c�R*c��M����J;��A���_����X'�ș ����yl��7(�S	<򚎫��o	�=�t�4ЊGC�g�:!�Ud��jY(�+X���b�("�H��!�8�x�ث�0矨�A&��!y\�#�K�\(������p딯k��9���0f�jL@����W�bD	.W���f�^`�*L�� ��;П�����5J`�2�xv�_�'����h��,!�4%�Hl[� ��X�5S�I^2y�8 B{��v���� �8�,��y�J�����MV�Lo�B4�R��p=[+��$d�w��+��<�h���N�d����:�+Ip�s\�Ae�����'�F��1WʢL��3�9�a����8�t��iN���ܙ+�#���B���8����G��(��kiK�0>�\ �ļx��Q�Cr{�̎���f;����l�n��L<w�gp*�-h��6��gƪ�y5l��+h�:mTf���]?����q X�azq�s�DJ¯��i�'��G;��"H  ��CV;�(�5rb��$m'��\;ǜ?6�����ʷP �\�{�bj�kt�|�lyQ��~9[�d9�ˁ�>�/�$�k��{�Y�z�FF���7j�^���E.,�� |�-W�u]A��5e֐�/MITi�;;��yJx&���SL���i�9�ɌY��|����nGMΆeY�wM8{}1G��l�y�x��zb7n��^*xD�֩T�4�Vf_#�
���)PE�|:#�W��qW�<ǒX��,�0JG��|2xv��ID���.�GN�S�3��A���k6���k�U�G91�k�����u�_)-����3�z���Xp�$�$mH���	B<V���(�����R^���8\]����j�2��m�1��@i��"��O8jD�f~������&�"/$$Λ�:g[fb�=���Q���4��n��}�0���Q��9~����]հ����`V�p
LJ�7���2cǡ ����aZ�/莻I�æ�N�B��5lv4��.ۻ�����*l�K�����L�;����դ�q���;���7��E$ ���6,����!�E���w��1��H��f�v�L���{��k���{x�&���۲g*y��+��qGsdX�^���T���/�%-��o앥�k��QjqwP�n"�O���M�&�&�������ߍMb����C���E.pŎ�3o򵁮�f���H�"cg�;�0�ĭ��E�ȗ��`ǁ���"v��3N�=X�=����\�PLڂ�3(����"�A��/�E���{��>�Q�Q�rp(8r�`�m%�Sza��l(+U��sMtime	o�>�e���o���e���InE����4m�.Q�a��#lF���*����7�d�p �_�Mo��í����=�-���'�