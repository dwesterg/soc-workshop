��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,�9���/���]N��E�]שF����1Z�#ߢ �d��o2����TS���(� ���3N����$�F5l�@
r9|~U����Q�d�ݮ��+�4%��C�Nx"n��<�.�����U��0T��'���w�Q�z�[��q0(w&���|6BP�4=�����ٴ3���t��W	�Aت�� ��a�͌�09�\�<\����� �f�v���%�z�M�7�:A�����k�;W�qNI&�Ǽ���Oj��PuS�ق�ӆ�k�>�N�ɔpe��$�t�1ĺǎkޫ�ΔZ��I�5�u9��D汁w�#h���,e��`���/k���ſï�&Ǎ����tX�.UI)�a���t$(#��"|pv��3�֐KW(���`̿����ݦ��iF�v�\��r��S;��ݡ�����hʧ�&`�
"E<ܲI�hՆ��|�����/4�Plb1��<aa^��@�}�`��:3϶-��Z�!�i|�?�o�h^�W��/�Y�<2�����%%��pO^A{�͉��S$��#U?��$EW>�����j;��F�>Ҍn�=x�?K�x뽿Aڭ�iY U�Ba����A���!��vE6��n��Z��������Uf�`�' Wa.	q�4E�)1A�G�AɆ9��{�oH���( �EDB��I�Դ��|�U�����0��Q�5�{�!F��%�m�p=�[M� o2bG�Z�\����R�jA�q�y�\x�S��	�l�h��3����j�|�b�*�+��X&㟓��iƹ�ۆpޤ�^d�qɔ>���=��K�y6g�u�C�q��:|7�TQ}μ�\i��9gZ,�x�9fsA���-�� ��	a�z{����Y\��#�G]��fs���9M
A(�~ugF�ܟ1ޙ��<auc�1%����Sl�Dϒ����S�_�����/1XeP�]�#�}���IGX*ʹ:��+�����G:�>س1O�[T.>MGG��Us�z�#�g  F�u���[A�\����S��n��lm���&i7Т
�s����g�W`�F*�u�[�(NF3TW��6��s�,N����X���e�/Ә��W�/oS��ߡK�R|W���̘O"�K�v�"�H�^����ȋ�xϪ�>�:P�OѫMw�ז���=L{�r��n+�8�9U�[����>�`~�fi
M:B?F���BMO�ح�YmbA#���[MV[�7%x���d늼�`���۲���;�ic���G�ˌu�!?��k�9T��?�J^x��uM�)�I��`c�!J��.~�=轂�w��g۴�g�}T ��2��u�e:��r#�t8��mc�,�	�觡%�T[״v�Q*��K����ItJ�[oC>��=�P��z8�"�^���hu�m�?4g.�#�f�̅��F�`�"���Nz o��-Ҳ�o����]��o%4 �������g��40��l��Nx8�]?~@(j�h�
����}��
bH����;Ig�g�9Z�y�ǋ�:�3	ï��#�<j2ak�<��\p�R�n�����@ў=�m<�+�)�[��Mva�l��.�{���!�.����˛${N��d�V�F���QU՜n�G���#O�C�xbeo<�@�I��}�0Y	Q�<h����{L��5_�� ����{�Pu�`I�ᰛ4��w��)�B��L�T�Ǵ��V*�-��4"�+z{�[��XV�@!�N�s{�v�8	Σ�ޘ����N��/��Frf��6TB���*	�_�le@�U<�� 4��f�L��l���vbލbV� M�Z�M�ט�>����u�/�E/�:���gz�v'����v�(h�4P���q�[Z�2�F@�x�i�mh�da������.�<
v���{��t7a�/}��^d��ӛ��`b6̀�8#գ�,Z�m�3��V}�Ǉ!��/������X�De�����!)���$��[�R���V���%!��_�J�5���*�M/�KrS>%�%ѹ��(��6r�P�NN.JdX���!�`��v�r�*�B�RU`��hKR<�r�o����X�>t��B1ɏ��-ĶJD�Nfxd�ę����HB.�Mf_#U6�rIʟvK� CF&���0_!&!{<s��'aZ,���|���
*��o��G%�P�S�=G�
�&[2�G�����y�r��Sq�2��~#쳶��b��jX�}u�	e*,�P[��i�@�4}Ճ�
3���^U��OQ-T-`+��y~ϒqg�������/�/��H�̻��[�2W׭tP���E�Ӣz�E
�6F�
;K�m����S��"�m?�X�w�T@8X�Lq�9]5��>�;�j9�~�|eCЕn2��\�	)N���Y}'8��)��Gi>�]#���qv؋e��e��P��ȏ:�)6��,�i�ր�afҚPpļ�O(X���àa��PC�<����!	�Q�vB�%��9u�cY*��>�$	U#�ey�H��K~%ţ��<��/v������X2 ��N4
\Z���=OkT�\�.y�23�C�k�f�nb᱓��/Wp��y�ؖʃS���YړyB�.��b�AY虬�x�0��j�\IA	ޅ�Ё8��X>���u$$���n:mq��W�����Ƚ=�-�@¥
1��)�ȵkl����.&���Z��1���;@:ԃmhɦ/�/�aP1�GH7�?�ݖ�<�8mB���`Y&�X�q����+vP�������,T2�
L�d���C��K����Ug�1��@�aF���O�~W�p)H���`�@�s�%�;���`$�sQ>g�em>3��$���f�D��{�Q�l�'�~�&���g��n�;t������;����h&�h�O��wu|P��m��F@�崍�LBӎ%«��=���$�˙w�x�4�x�����EZA��v�2��ո�ܒ�J���8�������`����2hf�ɓrr�/����z���֭|2ay�?�l�$�h@���ۮ+&ҟ��I�v�@b�n9�F6茖�����b+k�B%r�K���xC��R�A���2��E�̬KW��]%����lÀ�p>_�*ʟǥn��j�_*����,OoL5��O�Y���e��V�[�ޞA�=N���D�=vȻ�Zre�ٟ�_W��خ/��9�>G�e/�#��\��u�����h-R��7�xᒅe�+�ׇ�W��H�P��}#�A��J�AO�m*�?3_���6�X�� ���ɝwV���ތ_��B�,��yf�X��W�N�Q��]̑?��tM�Xr�2eQW�z�s�s>���
�(,���p�]q#��w��`�B8�A�"X��>-�g�1�f�7T���p���Y>
ܛ^0������@����$޴h�(�a����K�BSY���@�b�Rȝ]3!�C��P����xM#�s2�+���-5'���*�Cn��Eމג�R��&~`pΐ�ZS���Ė� ��0,)V��˴|G
�#ػ��:6n�hT�#�>�ׇ]�&����Tt����MKs+�C�!V���7�^DR�]�#��+�[�u�K�D(��9��t�S�ߊt�_���/�;�.��r+~���0���f�˚)塬�bl�'+a����8������b�f���k(���LSw;���ե��`#����{Yb!M��(��µ*�jD���b��G���a�wĎA��C�~<��n~� �h&xyP�}ft[����H�~�z�)aїn�P��3�(�܍��Y�y��n��&�W����7ޒ��۠�."�O�0W]�f�5��IN*1J���6���M���o/�/�f��G<�q_�4�-��]�í�7�N�G���p����z���gt�2���^���e�(=�ʘZg�R]�\TO�y�M��&�- �ڒ�u&Rq	>I�ew��2�8m�:&�7�U���#}�+:���f]t���s�^K�uփ�m�I�Mh2<��b��4�ԊQ3�����SC9Zi4�����*G�.��49#S
�v'[�9'L0�H��s����=���/������iу[�A����iŗ�B�Bڠ]?�A�1�Y����1'�>���٧1P^�|��"��z(��`�Y�w��=,�O��E�����2nG���A��~���P�g@�C/6 ��c�Vs�L��Z$b5�;Eur�:L<��Rpɥ:�O��_i�(u�0�T���������ؾ6���9��AG������`3$��[�h[�4V���6ěn��?�͍�[8�f���aJ�vE�ň�;Gs|t�Z�XS������;C��Z�-9��	a��>��R�(�l�y����|�ֻ{��?[�?nF`$mO�&��ٹ&[=.�+�H	��*|-�ҵ,#�UFĴ�7�έ@�{%�>�v�!�4�y���C0����6*��o��).��r�c�O����
p�]W�_�Ĩ���L���=#��{h1#�!�UQ�pwS7Uy��*4}����rU�ZA�����X3�ʝ[��W�5����Ǹ��M��)��O��&�[�k���e��o�	��M$_��V�A?�u#�n�c��0��6������K0�Pcq�56n��3�|�2sf��h��cr��:�Ҁ��&`EE/� _����Q#7�RI�XG$��Y>��{0s��������k�Y�Ǫ���I.M�ÉN�X����P��7�������h{��^�������B߬���Tu#�x���� ��Ëw0���2�8�������KD�=q�_��˯@���T(�d�h����� ��O�;4z��OnFF�۳~�v^x�bx��Z��I�{� i3����@?�D�~N�X���Ӷ��S<�np��B�簆�?M��<���Ts�\-���T��ϼ��w!en�T�p<yw/�	�[�q���H��|3s����LoF���F�_Z�32;I5�׶���U��	X���j%�Y9mMۘ�] N*�~� �����vV��7�P>��!���QD�sI!��k=J=[���-�}���Uj	^(�N���={%O!X�q ŧ�<W�Fj�|�%`�8]pX5R�CQ�e�4�@'>�� �;�T��}D@o?��@' �j�M���i�M����}��G8P��K_��6q�Qag@EG����!T��fQgt�-�����c[ѧ�ģ��♓�)xl�6�ӹ�CfY��B���e着!��f�n$�Ā:�CE/�
8
_��Me>�Y�t�W�Iڂ�9�p�e��t��V�����0��)
2�Ua�wx!c��.��C�Å�%���²9\�[���|�(2* a���0oG��N�����3�d�������s6 ����L����1������I{�J�k���U����J9eH�5�0�&��?;Y6 NC��$Jh��ٯ�C�ƝN^�t�\kZf6���`\�'�6��&q.e��%ML�j�&p-i���(�C�`iZ��~�s1RUV/�?=O��9�?@�d��^���`�>��b���1��x�y��
�T�	}��w"���1|�����>�X���Կ���K6�S�t��a,n�z
V�[D�����u^��°� �t�����' -�YC�y�q���%H*%�n\j��"G�
�(��*���,h;�� ȍ�nS|3C��w��¡xz�?��m��MR�vkZ�Em��79�/MERX��%�百{U��9Qf�T��`{�pɀS(O���ާ�%̗��W�>�������;I��.�0��e�h2�\4��X�j�<2H7&vu�*3�[�;��K��V��UI��.��S-�� ���!.Fxǖ
#��P�dUȭw�,T��B�z6�f
�D9���>���a�z�F\�kX~<��V�_�qd ��P�+W��F;ٟt��~��(�?�z�)��e̖U��pJ<V'�t��nN�ƾ�O��.ڵ5id�wa(���ۼ���irY�'�5�Ui4Az��'ݛ7���>s�z�lg����6�?��5)��Ip1�?Ϸ�;��D:�k��oV�2"��>-��)&ρ�o��b^�e#S8���v��%!� b�;����s������� 6f����-g�+l���˵�Ʉ�.#_$�G��5!-O�?R��U�����v��Zpk> ۟p��Bz���u���F
���pb�b��ZUixvO�2�e$��P�`��rH$��J�*��m�1.���kv ��i7&����3����1��[�u;�Mc�=UϜ�ع>������|@
���������Pc 旲}���^)�/Tq(�ȵ��#�Gd��i���w�F�o�Pd�s����v���#�r:�������k��X�o�w�e*��[��6��S��ɱ�����6�T��j�7I!:�/!���͚�2@q^����L�[�_z����|5�0a�ա��0i�p���l�$�h��_��� *�=���j��.ԍ#t�MU�SU8#�l
��YQ�}�V�b_�6�2.M��3G̊��!�:�$�k�p �5��Xs��&�h?���w�Tf�E2GS�f	w�U��a�}�L�`��:����D�xt��5w'L��a�f7~�3
ً5^s:E��I�IQ�C���8����|C=d�4����H�=�<m$Eָ�����CWs���P�4*��fK'C�'�3���x,������Ȓ��d��,U�4�����!|h����L���qa�qG�ZJ�$-�X	�8�^.��+��a��>��B�(&�'�|t�p�KZ��M�S�#�
�Kb�ETk��Uc� �D�V�*����,c��N�#H��"��l�~��xO,"��x9��ռ�G̓	���X�4��`�1�(f(P3k�~��fÓ#�	��`�K`t�hpl�����8F��@��aZ��	:����ez�W%��N&�".4�uoY��_�?A������O���W�Yb̡����I����Q�Y�����)!��~o)�����O%��X�^I|���Q��W��.���0�姛�z~��^{+]d[a:WO]GSL��}���N�T�;���)���ꟊ5��yP�AtW'O*A��DQ�\t&�zŐC�����~����e ē�g&�N�m�6�|}�f:�&�=�Y��j�JCn�̤E0_�A���-i��0px�N����Ғ,A���漘�K<t��,o���Q�*�P�5���Y�c��֮��#~�Z��� ����C�eW�a��T�h��r�WⳂ��Fo��zѸΙ�ٝ��#���ь�Ӻ?�J�G#����a>�6P���K�9�K�8�(��-�5x��<�S��� �NI��`��k����m%ASL��9����F�X�?Bu�	� GxL�����Al!��D9>�<5�&R�R�kԱ�`���ԋs���(/E)�}[�H<(�2uXqrDQN��Ψ�9�ޱ�%��NN0�jHר����J�GͪR ����y��ҏ�l�U��4��[@bQ[{lޓ�GDE�A�IUK^���w���]�����~"�[��.qt�-�c��>H���hҏ=EL +�S3%Q�g;�*MX���h��`�^����4�M�6�X\�x�(D���#�o�O�-��&�h�(!f ؼ��i����̴��mEE��L͈*��r�Ѝ+�S3��Q��|i��`�q���jK`�Zl|Wik:gq,O���u8�x�"�]�әΉDE��������K�j��+B����/DL�
Y,97�.�6��9f�2:8"�wh���4�{\[��@[ Y^ZW�F a!�˷�Ȥ��1Lh��OƱ�<�N-L]&u��2��=1�JG,�b��N6J:�x_2rQ"2�^����ݵOv�ǐ����3c�z��86���BA��W�L]���9��ϕb��|1�˦�l#��B��p����<:�r�C�"8��Te��^�(�=�o���ʓf�;���� {)d��e��8[��~.Π�No,��x��2��J��U:�ac�`����p�@"/��ˁ5L��\����|N[��T�v���������.��2���	k钸�L�v6,��w��'���xs�=|�6�״6Y�n���fnz��|�"�k�Ǒ�%�W�[/�@��m��\_(ͻ��)���X2�f!=w�7���B_h�0@���[��Uy�Ft�Sj���)8Ȩ��8>�@'m����U�x��L�98�J�0Ӵ��'��=��e�r������}S�,R�79xdyFە7FK�Eo�ZD��jj'�K��5W4(9��Uz��<�W��a���(u��|f�z��ǳk�6B~��R�	A*/Eh@���9G/���2DR9=B[��څ�VR1o^��AKY���Jv��kXw�VJ�4�4���<dgz���? jp����)��"5$r��/k,9Iq=S`��U��U�ewc���r�ٍ�h�ѹ'K��Cf���LB��T!��j=��P�����C� uAɝ��hݰ�-��W�9������:ڦB����54�{���<#l�/;�
�E�H�m�D�����E�jB�5x����M0����Q-oۆ�y�Yo]�m:��.A1���3o���Ă`�����X9��Z���Q�����X��~� e�^�,ݦ|�.�a�ۡ�[�B>�Q�� ��x����֓�D��r�nlr�q��I�9�M	s�lhvז#UrQ9O�y@ܪ&��z���:��M��U��!��j����/qyޑĹL�o��jy�-�n�Kci4��X���[���ӗkZ�F~t*��	Ҋ��=U�����RPMM�/L1�Ӣ-��"�'����^B�����H�ͭ+��l���:b���a��?��3f�>ڋ�4g����]QR�?�N9�<�6�>'�ω+=�M�CVdZ���{���?�;-�A,\W�� ��<tz$��X���<"�@� Z�������r�֥G"��x�rU��Ҕ��3R�6�V��F{���1T�n���=�����,�FyZ�ۣ}�[[V�O��1��!r#�F �׍�jl�|*��?(�.���6$������!)0)f�0"1�,�[���@f�
܅!�-yҌ�{��fo���:��yB��.���!��5���u���;�A�ٷ_�5���&0��M"�y6����K�`��FX��)qJV�N8t���P�9�u>%�}�f��$g�kf�E;�sf���*53����~�s�#0��Z{��m���W�Fow%4��T��R�?c>��P��w���2�Y��c�3�|W��aT7�ip��x"%��b3zIP��T~����M��V��]���5by���Z*4�k�nX��ܖ�/HY�Jr@O���o�$+hs��C��梺0�1d�D���C�c���m�����զ��Z��V&�b_�h�]Ə�_�H�s	'�5�Bd�8&�8~Q�7勼u�_�,�w�G/a+�������{�C�Dcc�"�I�hE�
� k�E�8��ڊg[h���,�JUӭ���	YBPO���q���5�<���$��:`ى� R��ҋ^n-V(`m5�6�":o��������]Anϛ�ԧ}���n��1yi7�o2N�5��&X��m��~f|���-�n��%�@�8[kת��$�F`��c���K��c�˱��!7�M���@�4@WY樿�0��
�xE��C�3�H����}G�P��Nx���J�YG��`H����&��+�P���w�'g��<Z-�5��+��  {
)A@�#l�sp�E����'.��9�z��v-7l�t�<a*�1�\G�!���\����c��
�	���']��g_� ,iĭj�SN�WH�l(��r�U���+B���r�U����E�O�I�b��z��a��a�bA<rWY?#{��Y��V�A�5�Fa<��%L�>(��`N!#U8ǡ�6�Ü<�,��"�I��$3%�F>���mV�*�L�9�B���+�P���<X[+�ר���8���Tx�JQ��� �3�Ǐ�m'����\FJ��I	:���B�o�(��X�5	��,]&/���3 y=���D�����ڜ��݄>FK%�(0����T�0�9;�eu�e#�bY�C�ݒ�O����F*��k�D�ԕ�S�ٕ*Bb6�z������8�(B�PRU��4p�	Ł�@���W;nYxH����%%etkt�U��i�î(�j@�f�T=�1�e?���S��h�G�����O���ȻA�	LD۫ѽZWdV�`{�t��D�ӆDW��EN����H�(5��k�gF��_hM1���1��A��O$C� �vm��MY�̑x[j�2H<I�E�wCqR�Q	U+j�v�Vj�V���}m���"}�c�Ϝ��0U�9�?3\�Ӑ����*]m=���˷�w��z��f���A�y1.	�F5�)���MH��d_�:�[�Ո��b �z�e`J2��>�ˣ�O�fV'W{���[ϝL�RA�T�Ɍn�%d�i�q��F}G��ó��_�nʊ^v�%��?���}˂6!@�_<���AOnk[#�@��0�#g��ۄ���I4�jfMg����%$9�����F����àlul��pI�d�(��I6�w#��J�4�f��b?Te*���x��&��L`\`��*jP}�9��7D��b"����x�״i�6���(��g	�q��y���1��lV����&��ߺ&(��u�X�t�yb���]
�d?�^�P\l�T��.�/���U��W-�z���bx�/ū��3z�u�׭Z�V#k��� �%Hh��t�5�f��*O�s�!n����\���*�J�-�hӺB���A/0wQ�d��9eҖX{g�#��x���(��^�}%&0N4���UH���s[{g�#]N�*�~b�z<�[<X���ƀ&�2 �2���~'�M�5|���-%�&g^/5�n���k:\�jU{Jכ�AYz�@U�S���:�4_ߍ��ո��8�~l�V��#�j&׮�K�]
�.��=" x���THQ�E
Ef�;H�b0�͋���<�翞�����cH��?mT҇�K��*&Μ�|��i!6�����}T��Hּ��o�9'-�,Q�
���_<8l����k�ַ�܋�R����O���>�H�8rN�b�X�/G -Ay���e��t
̕Xބ�uЂI'�ۦg�[|�}2lI�k�l!�TnT>'��IGQ�zM��#T����Tl��N��#i�|^��.g�����Z��w���Rs�����s�fk�8I�������lT��Jڲ��L1�᧕ԥ��:e6Z��Lc-a>*�2��b"��9ǉ�V�:�H��9�XE��m9�p�?GŁ���7���~�!�$>A.���E4"�Q��cX���FWC� Shn�?�)
��*~]/�{�~��mŻ[�t0L#c�%>r��-��<,�M�'yk�ځS��0T0��50kR�k�v�M���砳��z8�ϸG�h��I����0��/)$v���S^��X9�1���jS�\[R����D���#��hp�z��m������DA�Kh0�)mbF���4��R{��`�3.{��W�v�5l��p��Q�Ζ�? �*
W�W��-��	������v�$;�Hn$rHB�$3����	U$��bH �跉���J�-�T�]�6����Z�0l��`���WlQz_*�ĉA�e��ߴ��ҏ��oP�X��P+�T,�ñ�0�6��9V�IdW������[<�r�� ��m*s�}���?&R���8��m {.����{���;e����C�_m`��잞�\���!��A��K~�Bc5� ���Z�\u��
��c������|���U��v*}�{�%�S�Ej�]C�� $�:�'i���e�b�o�ES��I�N�}&��;^��������+]�� Ν�a|�v(���T9OFBZj.ND�Ӟ�c �9i�ˑ��P�:4�����SER]�Ĝ��$ޓH_�&�ʋ���� ��|Q(�L[}đ�����-���s�V��
[�b�)���p@:Y_��J��E�ߡ�����3�&�����h/:.	�"k^z�]x.^��Z�8,��t'R<f�<���o��.��BRf�/��C&E�Ql��z3�?�j���w��g?ʢ*��@p0�SlڸQ���B�C�`�D�2�1�˝�+��A���<� �p�zf�^�\YZ���x�B�)o�h��e%#T��,�0ts|?��>�m�Y.�"��S~:����	��5XKe�i�h�o��.͔{KT�m�B�*[�"ǋ���W��+3�G��[Q*�=��ԁZ��f�C���}�y�`��ï�+�	�� .��Ȍ�wZ_��3I�O�)#��0�B�t�G�#�+:`�͂���k�n��(X_$z��1;m�DL�P@��m�q5 X~�_{��q?���l��e�f�4V끂#&DYĖ_⟽���=wٖX�K$�LQ����DQbG�0�s�"�Yϭt}4�! G8��YyT\p3�; iM� ��6F����q�`2�B�`		�>[��/���E���g� �r`���[$ʪ�@F�-�C`OC�l@B�Z�_��u�3ƌfK�h�:�mΚw�w�D����F�	>5�Ek��b]R�G��9іd�0q�J�K���-T\+ý*�ϴr\���Dv��'��U��J�a����7snN<��u���p�f_n�$�_ �I$ry��P�XN����}��	��<��9�	_��(�il�Σ1:�H܇~@G�|��ߐ�5�F��T�{���|!�_�u�:o�m�(ҫ�Z,�pn����.V�Џ���&ez.�8k{zf��" 	��M��[>�b *��~Ab4m1�uu3�)fV�+j����5�\7�E���;�[����3<������nXפ�	�����@�X�T��h�������o�X! ���-�*T��C&������9��c~�RE���Y7��yh�Y��O�µ���k�q�Ϋ�@��»�����������35_rڢVN��vϭI q��2<V��x��:�o�]PCܳƚmA����3��x�:ɓ ������_�9/�.%�@ҙ�(�rł�zf9F���i����I�m-�����g;$ݞX��,��U0���ً�.��ϻ^㠰ó;�ʎm�fPB(W'M}�]���wH˺����&�P����,��7@�<�{�hMMQ�rK�Z�	��m|��-z�,)!��`� 	M�ɡ��ǅ�Wz9�<�ۈ�t�foX|���i����-|��g���t��4/.�lt�y-)����4[(8qd[��f�ٳt��*�a�1����n�0���헞J�5HN�s}�Xx�&ۀk]�O!'���9�S�l\�$�ܚ����
G$������^���9�WÕ�{}����D3@ �Jx
o�ɔ����/����ڃhV���/)=�,����_"��u&+�	Y<y�K�ٕa�1~E�[�;�+�����1�8��7yμU˭�:�����;�:/9�HdI�h`�RZ�w�ئ�)�L�u'��{9�T6�� �/�~��	�>d���T[ĸ��@1�OIu�(��-a���z����ܹ� ������Ŀֆh�Y��L<X�P����%�}��jP�ŉ���]�I����B2ɠ�
����}c	s�G�֣���Y�%�f�s�`^x��Ċ#ɦb���H�+�Jn�F.Dwr'CG�LE{͹�������h�c�n��Q��n�DZ��=�>r�~ϤՔ���']��eٲ�������+LU�����]LWq�e�lX�&��VA5�4kV�J��B�J��3�]:��-4��O�*֤��3����{�W^RS��7wn��F�"Fpr�\ห��~�,�D���k�KГ�����2���(�)����}G�DAƑ�6Sl1z��w6�S6%w���z�SX�Agzj����.��ù6/j%MW�og|h���է���-��h ���%�,��a�1�'�rI�3���(G_qR�|�����zc��=u�M���_U-盧�����[��$����V�&A�%�Uض#�'�3^��z[�?��>Ce3�������X<�	S[�\�g�Q��f��(��{0�`�=�A1I��aJ+uT�6KMթ�]��B\�7��$C��!�1Q����]�ڬ�c��| ����T+�s4[,�W����,,��Ǫ�Kr��m<�$�[� ]���y������g�*q�=���q:�%��1Tݜ~%_I�;�q�}�]����^t�N���h��tiJ���n���&�����X�҅�� ��A�������^�5��K$�!伖����S�c��������g��[ߖ3��zv�L)�"D6��
mPI�oL�{P�6v&ޑ�J}*d0�#�\0�	m�G5%3=��Y�S/���<�P)pL��|`OyIfLy|
�ח�c�����	x��W�(ߥ5Ve	��V�\�78.�X�1'�d�RY�!bG�\�ϓE�%���w8uE� ľ��U@dn/AV4��ǉ��kz�3�N�Gߛ�IYë�� ��zI���)���v
�$�W~��̟�8�WYkf���� �K��U�0���[���Rk?֤ӣ	���6-A�8�ņ��(��m+��(:e�����X�M�6�#��}�:)���3s���0�$gD(@1��?��mLO����1�݋�'s&�*B�J6�6��)�q��-4�����V�9(���}垻^�^"���s���+�wU�%M��V��6��K��ٯ�5�: @4�O)<U� �x0����p
o`��">x��עa����_��0��^(P��E�@�a,��cY�{C~��̖��m�Hp#\Bج�r��[�n/Z�`̕����<
�A��J��$=2����3~-Q����8{��a�6����{���.��00Y+����bk��n>:�쓸���A1���,�w��j�v�,�,)c;N*�(�t�1��)�� �$�o<�A7B�?J`��V� �[�
��eb���h�ϳC-�x�o�~�*.���y�[n����k�3otv�`��z 5�1�>Bq��n2,��O���i���L@I��F'����-����ד��5��=�=#Apj��g4�I�� �3x$���_�&�rzڠ��'���SU�S�S�j�~[C�Wyp�u�`|��pπ1{c��Ğ���pfm�\|5�n�n|�����p����0���Yʞ�G�<>g����pBT��(2-�Ӭv�fI|2�	;-�f��#�$2���8� M�p�d�=WR�؏����/1<��KY�=P��Zg���֨�1P����:�N�Pd��MM�dF�t+������~I�,LB�%XwL��|�W��	��Ej%i�A�V�@GL �@gB<����������!l0dau���	.$D�/�н�m~�����H��lj���ٶ:d��=�;�@'�� ��f�Y5�У�DB�-g崍�n��[�:X� L�xߎ�+�u�w�Co2u�����Z��E�M��wDVƳ�@��*�ڹa�U�$Z��84����4��L����IQ9��7���/+�H�(�eΛ���O�2-�b�ʸkS�d���k_�naR�8%� I儰�w"��3�%���� �Z(��{������*�.v��!�j�vpe���m�?8�CcԾ>���Rj�a��)Bka8,�_�R#��JgJ�2�w�9���,��TX�����c Ku���4ǽ�Jf���p ӑ�aO�a7��n���xt��vI�r���Q���7�����uIti���G�y�	�X%k��>(�M�J�	\"�@?�����xM�߈]l]C�F���1p�}{�ĨF�+�V]YW^Wʄc�~JwG�S����h{M�t�r5���f�Ϝ�^�NBA�ž̔H3���ӱA��Ča��mE�@y�e���R�SxU���"v�us���'ڋ�b�{�����5�؂���:0�#y�Ե��߲�9������^�pt���ҼJ�����b �g��"�A$+��'��/X�d[�2��T���%�iލ����y7�}��7t0V������x"�RmU,���CX�ҋ�Ǵ{���ڿ�#�De��v�6�T7v��.��e T�3���;]hP	�_.�RIh�O�d��coF����9�����0v<vU�r1؜V�#����|�����A�Zc�PK���n�\��f#FX��B�3QPc�w��
��@����"��0X�Im�N�T҃˶3�Ʃ4�I�僶zU)���i�y�%_�7M�ח��S���³�	��PJ� ���U����2�X�Ԩ:M��fs�YUJ���7�|��4���$:��	�gQێ��=�ә�Һ���D1�^.�&cn_ �ާ�	���q���$T�-VB;*Q�#7��S��ˁ{�/F�7$�q1�U����b�b��5S���R��~��#��$ ���-��ߥ� �F-S��<��֊2^�z7��ܜ�a�Vڈn�sЗ
`\~d��	p����SQ��W�P��_�Խ7��yD�MU��3ڜ��2'�B�*1CSc�l+��4hܮ(�~n5��&�I�� �֝?6�֏��ƀ���3PVUP�,k�3N�/��J�*�(�G��p�+`���0:��&h�i/�Tg�۠�N���/[��~Z�21��X!����մ���}jK��JU�kX���P��=���`y�ŕ�c��4ڐ�-�V[bυS�5P>���O�2�ӪE�d��j�M�	�̸g����Z���5��[�!�)%'�.���ب+�6�C2 z.��w�rM�:fV?h/�����/��G�;��z@uRa+U���G�8.�B���M�:N����?��y�6�y��� �c�RԬ��SCy��+��=�V�܈'��Rp��X�y/�-�T/H��v�&a�ט�b])>J���H$O��@P��A��*���l?,@82���֢	�1����K3�C��X�����4W6�Pw)
����k=��.�@:��̿c�j��8ȹ�T9��:��:Q-Gk��6Ǔ���!h��� X�)�,�Zd!k>�<��KP�av�w	���"^qln�J_̎�?7;lΡXw���'R� �vk�w���6�<��ז��
SE}�65Fl(E�	Az!��"�r��
�Ƈ�D���XE��Z���Q�w����%v/9�࿎adܦ�	�2qMP䯴���ދy�V����
c��B�Ho�]��I2��X���w�U�n�C����;f�X��Ϗll���?tF�	�\�Q�Y��%5uٍ�F	��n�kbz@�:��	ń3�uz(���N��LV���7�����d8 w64�1=H�i�_-"?�qd��k�ĒC�
�@�Y'��M���+�6y��a!�v	Z쿅T� !nÏY&�jN�s,�l��sP#xˈt!��[���!��Wxi�'��z���q��T�D��EPإ#��`{w#��"2p� |���v�se�V5۹��S�[}9�	Zޝ���xZ>"u����
��%G]wWJ=M���g<$zy�d��- ���t��%e� �;D��K��m֔X�W����M[�TF�w��;�����4D����d�A��g��Ŗ�3����A@���v����DG�*�/�,�'4�$���d%�X��s���|N-Ei�M����4�׬jl�f���j)�opcKjn����J6uP�r���*�ی����L���W����=����ġ����-%)X�{Np�����񎢈��)�r+���E�w�F�V���������ch�+�5�P*�����0�^��b�F\%�*�-�[�W�-��U8BQO|�����l���tw0�z|QY�Zf�c`.�|�'�4���1�� �뼬�ιL;��nH�2�����`C���x�	ԔCG^�W�'�?ɂ���lR���@/�9X9/��/� ��\W�-�B���8���ǪMFւOҩ����Ɉ�j�p�vX�Ω��n���x���R=#;1K���A;�[:2��.ӵ�|��&|��u�����Y�\��<����`-.�)`�&�`e��6�7�x����z��'��x����,;|�!���)Ùrs%���?Ю~��O�}�a���a�k��0��$�3Q�xj��p �12�K38��9�	̓������̝>����zӱ��&�C�U01���e7]������ao��T@"t)(��Ke��nѽ毢C�hެ��fSEG��V��@�3�pU/.i]ځ���v�'V6��.l8*CC��;]���q8�+��3s��Ŵ`]��Ԑ!Vt	S�e�Yh����,�RJ .���ǕUaO��,��޵W����w�)o됾�3#{[XF��\3���r�?b�G�?j�xrӚv�<���g7��܆��͇��<.2&�)av����|��޲7�Ϝ���ﳎV��،�-��ϓ�:�v��<#ܻ�����82�}�.�(�ڹ܄j:��4o��2t��d�}�<	���{D��oC�KN,�z����s9�u|�4�1_�g�1��=�ʳem���i��.*dmp�"I�O�kB81 ��kwM�$�xi:�Wy�i�b�KƄѫ�����N�O�b8��(Ig�J,�g�3?��zD���D�oV�/���%"U�D�����u6�k�g�3Z�Qm�-�Xo׸��n�o���a��y��A���R��"�����|� ��Rx�g����b8��Q�;6�ם9�����[�v�7S�%�r?Lq���-]�K$�:�^F/��r�<�f�;�=�'�b�:�VCmN����g������<<�SmoY|��Q�C86e���^��j���ٸ��.��0[abx���*k"��F!	���O����QH6���z� w�!$E�nI�H�괷��\�A ;���	��q���I�����U/��%0' D��C��LZwK]6��k����4#|7��@�����RV���-���:��.���A��3=��ì0�/[eB�U�L::��x)H��y���ak�'D�M������<0JZ���@�Ϋ&��'��6b��1���͓iWօfF�Y��Z��5�4�1����+�٧��)�m��9��}%�]~���Z�o�%ULя�	4�������2>���q�h���b�D鴧^;����d���i��(�ө�S�D�0Ɔ���Ҡ�⺾#KRmؾ��2_7X��F���l�-}[h���e��gh��~�;��D���T�]�V��NA� C֜A���0=��h��l
o3�riA{�?�}K���&�]�l��������?��Y�LZa�;�k� ��I�D��k����蛅E�C�py��<B����{+�s�����8"^!_5�34���=8�	KU��]�A����,Ps�TM�'@��+���SW���m�ey���r�«e�2���0�W]IO��i���������R�#��`�߆��J��S���
g�oa��ur]5@�*� v|�?�����-!�g^$�#�C��aL,��Sߎ �.�-=�^1|�<MA�c������\�e���\��W���Y,-X�Bl:a��Lp~-{<e����P�.'����x<�@&��J�S��
� ����3�j��b�HEL�Y�9w%P�G/XL����>[�~�]@�Ԋ܏��ن�9��S /�|�u=�͕ۄv>��r���Df�6b��Ě�"��/���J۸�8`�7(�ʶ����(��y�C˫�u�?�e�:{@�aȎ�g7*��
��[����"�]�E�G�Od��u�1_/$x�[@]fܕQ�s��c�`�g+�����v^T�"����̢��L�h�
Va�:�Wle���$�� Vl���|��ˮ����^��fzM�r�[��X!���>M�6�?c�DY��O���̘�n�����K��Rl�8W�*g	M@겓�'�{��i��� ��E7���ՑQ�<SNNR�6�⩿���4' �2�շG�SH�FF薓�xu��HΔr}�hk��JԽCfOr$Pwى�D(�+�>��ć�����)��R��.*0֤��()9Z�:����0%�S��qP\> ����x�՗�lC��2!���	>BX��"-�U@f��O�?kJ��N�A"@ ��C#�cw*r.�8њ��!�Nz�K��A$
C~:�u=���j�7���I�U�*�?�����RV���t
��-�ՠ?]�U���LI���_��{ج���>n�Ї�#�7�ޜ�tgƨbĕ4�E������9$l8دb�7���N�MM��h0M�I���X�ĵ��7���cu��:���@��3�.v��TB�Mb8d�&�p2��w�=ΡbK[�f�q�^��z�9�wC-�Pe�6+ ��d쐾``��)d�˒d�0��z�U����P��>�J@���`[@� 4�1�Gf��)u���|���4Y�l�	?�D���}2u^D������Y�o��(tʙ�7��~��W�̎a���@i���|���h����O���U�H��b_��sd�%>Sdo��qH��*��Wb
ct��0Ò^�+��MH��w���B�]Q+}̟��h����n��q���ၽ�c���P��jӗ�
Q/G}��UᘔW�cY�[��j��\}Kw��؅�|7 ���>��tu����j<f�x!i���8�Z�!D��H�iM�8�7q^�{��^�� d\��`ld�V\A�X�.����3������#�%;���
�3_��>{_����s��o�E?�rހ��~�тl��x
ߢ�I���z+,�H�F)�~�j��bٳ4�:��9�j%�����[4�c���)�\��|"!����v�4�<�w�d����ބ��,J'g"]�iy�<M���V�>��(1P$t��n#F�6���!Ҥ��1$m�[�:���L��^@�q������{�]��g�	�~���7/u5pW�7�u�v{s�~C��Ot�$<�	w��H@$�8�c�FIj��� [g�BM��	��_i�(�G�}c|~������@������~������Z㽪0"�:{8;Os�g�I���6-�
z�j�/�8�_3e�n �t���d�1������g%k`恺YJ����&��p�"�<�'6�^�����.A��KH���r2w�<�,� e �����,
��������3�B�����0&�rt��׿67Q�p� S� ����'b/����lt��k-�x�3[9C\�����]豻kp�I3��C6��	V�G���q� *�Ͳ�6�F�nu��aA�4REC���9�mJ���8�����*�*I,�=�������tWOUׯ�#و]��j�VO\��l���/r��@�]�@�hI�Yq=yUd���S�y!>*��Lw(%G�]B���fMT�!�(,�͞�UqWH���9_��Dó����K �[Y��� ;�g�SY�&mĈ�d����K����9��&��-�3�����d� 6;'��rѹ�\Գ�e��^�� ˖�P'� ج1UB5�o�"���싃e{�8�5&��Ư�`�(Ī�+V��M��FHk����3������&��H�O/�N��31��z�mzo�M��(7x�����	x=�6�9����/[��S���Sbn�v
10[�1����Q��l��!�Z޸҆wR������B�Z�3�<�k�;����[Yg��%-n�{�Ho��C�&;�$Z|��r*���2&��K����Tt���[Bl4Em���׻|%��.���F�{�g=�=u������P��&�ײ�ܰ4�@�(��$dvh�OY�����W#	������,.��x�H��K�~QFh�dZ�٣�Yk+��"���[ ���)]�f�T4��
��rg�#��6E�D�B�w�4���L���OVzCe�	��L>�pȝ�{��MDrh�(�;��ji�c+�#� �U��σ�t5+����1W������r��Af�Q&���eA�Ϩ؄,��a��o�l�װ���F�iw�p�ߙ3����s��J
��aR���v�\���u~���ӧ������6�Ʌ���ܘ1�`y_�ۼ������Xw��K�j���d�!j�O����gFJc��ٕ�b�#���E����t�$���_��T@�D�W�l��Y��=��Vk��mW@��״Y* f	��Q��:Af���f��Q^9>�ޟf1�rt�c_��>��]42!��6_C��ļ�%���Wѫ�d��3S-2�H1)����p�UG=�漩��a��O�c˲>����|�I�Q�@�	�.g��N��vʮv
�9t����L�7��ˣ�r\�$�$uD46ch��%kHտթ��
�5^~�3o��{��������irfg���c����Z��N���V �v��2�,��$�b�����p
w5���vM�FA�2��oH��B�W�/���!������	�:T�يB�̻p����ceQ�=[MrvS-]8=��6����"���=c�C�*�g �=3�eC�GV�v
��y�,ѩ:���@��F��~G��F��h��l�>����ǝU�K��m��v�"��*�B�11&�z�m`�+�V{��E����R����Y�d#rKW�G@�n2C���.�P� !�f��2��g�������5��QJ�"�[{O�U�e�Ç�^Q �� ���	��n���7-,b�$����L3���h~����B�F�r�X��x����ƫ9��O,_gH��ה�u��ti?B�("�$�a���, ��M��_�)3-�� )@w��C�snk�^�����6P�3?���+ll�F �E���{�wa�(�WK*gdPǆ�=K��`u�o���k���o�Q���A�-�m� ���X�5(Z:����[l���� bGU�V�\ɒ�.�`I҈��2� S8Ĉ��������k4�e���P�}d�ʍ�{6�8ǚ;ɛ�P�C�2~��?q�n�\J���I(x��b'(�擉2���U��z����y��Ԕ���7v̖>ﬡ�\y������2���K�u�q������们S> q|���Ҁ��
�I��l�� kwVШxJ��� �C!{�?�_�=wn��ʚ�-�n&0��X�20���W�jb׎MU#������˹�]%�������:��do8�J;�6SA"��\�M��C�S�b����-Ěm+Y�M��4%�&��.�eO��>���o��Pݩ��x���J��ro��mpYdQmP'�]W�Y;��2��+�kp���Bw"�n��Ym����6�L�
V��7e�U�6W~Wck��h�dȂ�迓[ZF���	$���=&��0Nnփ�o[��^��'b��0G�RːE�wqC��$�BO.z��#&�>�+�-&�������c#���b����o_���J��ǔܒ�;MF*�TKB:�	A�l}�$��aR�Щ�C�`5V�Y��L��n�O@
7�B�´�%:][�H����;�w�8&�����0{�6��9��.A�P��ޞr�~-{��nV}}�Xw���C�?��35k�X�[c����)x������Z��h;OIZ��r:p^�Y��|7_=v�y�6^lwza)�?�l+ѷDMD��ퟍ/.	���g'o0�)�eKN�v��}��V�@e�Wx�mmE���f�c�f�0jE�����@�6R��L=��Y���kl�R]XPߠ��3*
N*�t�z�Ŏ�g��"�8y�	 �	08�B9��j����}$Q��/GL�<���
;:O�3�CGDwz��
����D����=n�b�;jɂ��6Rz΅_������X=z���>�P���n}�dE�
Ѝ?���uO�;�`I����lJ�GJ� �_��bt��_�|:���
�KP��/8�JHː坠L(-�/��5w�ϗз��jG�5%����W4��
a,)���s:"����"�͵��Δ���R��c/�s� �6&���u�S4�n�B�(5��S�t�D(⸖������_l��v��?��@ӵ-�r�uⵗ�����Ԩx���ђ,�<=��LM((��S�����#01��{)
������2��$���
�a�}dz_ރg�m��iy{���J�H�{[K�����Z�x?^=#�y��Tu����*� �ך�	cD�ᳩ\���?�����s�+���Wϋe��W4Uw���l"Jߣ�]�q��u�d�7����D��_e��<�F� +�&��	����.��|y���^ٜ���H�(b�A������	�)����+�]S�ń��]�m�3�fEØ�)�	�ĻXQ5Ir��=�X���)kcb|U"�J��n����7q� U
GY��T.`�bs�6���p9g���W�8��AL>����0��	Y�� S��`�k�mv�ȯ:2d�oIQ&���G�B��y�>:�f/V��_,4E���Q��T�PF��+P�<�S��bZ��h�T��8�!��Y�ęv�dBง�ћ��T��.!���3L�s�7Z.(ژF�r��Y��M�ET�+ypT��H��|�$7�%L�\���$����LdAg�,�_8�E��������w�3ﯻ���d���͑�O�S7@��ϵ�^�͟y�qUn�����������,�_!7�5�C�m>�P���c���ZnXh񕍀UO	��rЉ��)��o�o�^r�.�Wh��ů���-�5����u9�O$��(��R����Owcz�)2�/�p�?i�1���7k�H03��W:
(H!�l�j�ڍ�F1�-�jt��6��ē��M�9�3�t2D@)�V��l={0(��4�
	5��P��is�Sz�#G'c��+aA#�%L�lCU�P�6�/Q
����#ȣ�5�-=�D�/t*A�i�އ�Ȕ�E(�Y� ��+Bva\y����b��
�	-�Tv��oK�A^�y����vP��?<��"��5�5�%���b��n�_H�,O�n�5�%ހx�H���m,�^�?Ch6�4p�����G�l��2woH�Y���Q\pb��g�����@���|��K-yJ?�]��A^}	�D��;tN݌l�����7�N�*��j�|�,����=߽�2U*
��e�����xsJd�z<����^����XBU"�r�
*���k��M?��Nv�`��e|T.*�8�������&!~�lϩ��z�|�o���������,�J�ɦ���ǆ�\��CP�K0�#��n_oɀ���ww^*���x[�Ap!�m��2gb*��=��^8�3���ӯʫn��4�OF0>H���F��B��4K(aDO�V}y7Ǹ7I{!"�0N*��9D�ŋjB����@G���6��y��U��z����{�}��2�]k&�ȳf�L�-1�?�1HPO��~�WYN�|yO�{������@#���K���;[g�s���m�Q�Y��Ӗ�]�@������a�&�I6Y��:q�^�4р�!�=~.)�on�[��e�z7�	�O����VK�������,����)�0<�dk꿉�g��qRI��v}T[	&��IZ(��e�|���Ow�0>�822�X<n����o+�(Bߛ*=�@jfS��㒉e���)SQg�uJ�O;pľg^9�Rm��wUjW�oX��|�Aͧ���b�X�_�}J�R*��`S�f�1�)���h�Hv�T/��/���_g�� �]_Q�򊯗��!��d����~�a9���OL����5��Z��y6���Pv"5d_I�����G�nm���T|���xƂdں����YW���`p���W����r�G��3joM��x"�XS0^ޒf��rޖ�����;_@1�ڨ]��W�!�PeWY��`df6����ԃ�u(*�A�^2�W�}{w�eόw�D�n���嬆�F��D?��W�[�U}֮��
t_ӫE�JW6^E�͊���-M"�0�d%��b���B�We����p��N�k�cs�@�{Y͌Ǘ�S�����}k]Vȑ_7+�C�֨SNr6��bmr��؂m�f`sc��N3Ov�����|du�$����o�1� �Ѡ=쭏D�/��S<�n��ן�Էf��m!�R�/��3�n�/�&>�꜈�|i����ѵΩy�R�l�7cT����q�#��S �1r�Ψ�m����ϭ�����%1�Aɒo�,h�<?�/�D��oo��b�#ߥDƧ�Bi{>�S̿�H�R���2t���aOʏ���}#�����'�#¢�9j���c9��~ij�ב�/��p������@5$Z��6��)���.�@�����"T����0�n����Ƣ��K�b3���`C8��NKhcA��୪Su�8����\J���"��5.��{ /aڣ(1;x�l�r6����� ��W<�(����$O ��)�P���Ƿ����z��$;Y*��]B�^/��� ԏw���%Hs�O�b0�O��&a�B������OOg�9C�)	�ء��XQ����R���՜�V�,J�6A-sR�l�O#rV���mϹ�?<�&��ǊAD*csh. ��R��� h˵�fO�9�;�M�瓚���62G���| }�\;b�[�<Rq��Km�������~�)��:�/&�Q��1����ߐ�#"��wI�
��D�_*?�䝐 �_@������mZ���/:�VU��hyt�������r{�Z�kԷ��_�����������T���f]��O U���G	ʰ��t�Ϫ,i�%' 8[֣.�x�ˋaR�|!g���T��X�C@�C:(X�|�����1��`6�-	�����kz�n�{EL�ᒇ�3�S���r�R&�3w�5y��ivYwhi��^�1dU��*a%]����G~0�$�Hk���h��.A���{�v�>3�0&���|��_6��\	gϷ�Wu�b�t"KJ6f��G�P��˲��h�+�+��K�M��&�΅�9������s�X`S�#�� k��3l
l�d��!���2ȂG�����>!?��GB�ȫ৓̰F�7����]8,{��r�v^��ů1t`D}4�~71왏0��ƻ�v�/��խ|���?D{�5��jO���rQc!~B�FBE�+9 �| p�T��'�S,��ໞE�|�J���n��:w�j��N���W��~�'O	��#���5F��zVd�緾x�c���b$�o@����	n�%RtD߄�8#�f������>}�L���^V���^�����D�y���o$Q|�
��R�A�R�Ͷ��SxE��=����Q�g%$b�-������F`C���O�P�C�!mZ	�j�t���A�C�Y���Ҵ���K*��X�9y�A-^���C4~���@ �P9�V�!�Ys+�An�V0��u����Z��k���F"�Ҕ_�#��ZC�|�%��v��|��$r��E.u���_��-�n⾨�ʜ��B/���� p{W~)ְ�@?��g�$u�L�p�q�>^n��X�V�|�.����(�g���'��P<b��$�2H���y��`�劲#~��!�T��`�\&��t�s#�y6�~����a��tC����X}U?�֞��_T�wnz1��?
*���͛
Xx0XCו~���P�ʋM���"�k��&���K�o�bOV�kg���L�3|�\H�7�(�]`^���η߷{�CXJ}���45��j�#�5�|tT��J��jI����e�CqCg#X���iX~'�e`��������%ٯ��'�@K���R�nx���N�����ͬ��w�-��I�;Z�,9����9(�!��3�|�N�yԚ<}�2�ߙG�ua+T���kڽbg��}@.�+��u���W�Tr��^��"L��Ne���L��V?�0ѻg�����>���*`H���i|�}.�6� 1�u����%-�<�;�M�70��0�գ��v׻�M���o����l��N�/B����ΕC��������u
�u)�D���`Ï4k�s�[�{,�4���9*3jۣވ.�¡����-ū�WB�tFpm��
3��KsiE�{�|b>H*��NҸ�'F�.&��ɳu���J��أT=��^��J	���Eľ���,*@z�.<oC�<�Po�>�$�c��:��QRVC�,�[1� ���c�i���k8�'��>��`��[�[q��/X2�L��r�
[^o�q�5��h��h˔�D�\��)����CWYl�r�:���6�3�C��4d���{H�Q6��D���E?v�V,Cp��q��-�Z��߿��� �݈5n甘�x<�m�]�߰�S��)��ֶ�˵�Ŝ��k�/��
��]��E�-�����L�7�J�>��5�u{��/�&+<�n�F1I,*Zũ� H�z6sy��Hӓ�ҒV8�v����˸�A+!����+xS��g+{���&�k��j|��w9)����)��E�Α�TAg�	X({@za�Z�fj�7|�#DX( O6��s�8�h$%� �r�����h���(��/.�U^�e w:l�A�pR���!U�[&��Ӱ2�"�R>4}�x�U�ݥ+qgc\�hO���c駤��RȱBqj4<:��͂�!{�/�@^(�v�<z74n�%P�������hn2Z�¨@���Fs+�C������F���N�C��0�q�d���<㥧6	zl,�VJ�`�vJ|6Z0E�4�weq��cNqz�x�x���aE,#uZL��b�	!��ANS�G"�eQJ�����rIW*�0�+���0u�IE�qƐ�8Iy����J	(�j5��6��N���x�e�;<(ȡ;MS�ޭR��x�OjL,�׻�;o�7+�a��Ɠ����X.e��Pڹ ,>_� wT����S^� ���]����L�DC�ϧ�۷�<�oݼz��d���A='+(��m����Cd����2���%Z�m氭癚�e*��s8��9'M����e U{���"NX��z��AT�����C�}���y@�f��ɶ\�L`1�Nnm��7y��{D�c��N���O֗b.4��ǧ�$x��P����Je#�>�%(�j�a�#���>���B�C�Z��5����M���D�;�p�BUǳ���T��jo��M`k��>�7&��u��t��q��*P�5�xF�0`��:�m��b�e��cÌ ��0E���U(��_��z���j!OE�^Z�1l��^H�=d�!l�4"Ji���f�b�h�X[2�n2�rʶT��j3(��U���X����^.�b����b�h�8V�Y&�����p�@�%�����R��nI0�l�ʹ��ٿ��ڄ�v�}H�c�^�`ɒ'�vp�������z�q����A�]��;����L�y%�-����|�3M��F8?��H7h`;T���AE$L	�}������g��UF��V�����D��_�;�g���y���^~I��c��?>����n��h�T�C�g�Ҙ�6��R�8H�T��eK��m�Z�D�(/;�{�A�[4Ŧ��6���t>bZ�+?2���,�ǖ4
�?�����R=9,mH���X�@ ~�?��Pu�kzY5���4몦��i͈rF�X�\��I��f�OC3U�'��o���l�
�k��k��}	������=��
���=�6z(�ˍ[��Դ������$�MB��m�8q�y9�ƺB~K�D�F�H�do�h�~F���Zϖ!�ȟ��E����I:�(st��U笰} �=-�!�6�I��v�{��}��������t�ȥ��}j^�M�����ފ�XC�g%�~O�&��ސ���1���W����T"��q5n��-6`����ж�uuc��̒M�!�0_����W)�l:V�E��>S��Lg�Q� �n$L����
N� E� s#W;X�����% ��7�T�3�H��.
���������'S/�Y��-�?x���:f��tt����-uE��n�3@ѫƋ�q����F�C3�n.U�|��v��ӗO�v��a��t�؜��&���xdB�,y������ժ��7q�0	y��4+��ƃ�#��I�|�_���❺�(7xށ�s�����S,�H��,y��4��{mm�7F�L��+�8����H�Q��p<��r-]j�[��Mvo����]_~;��I�Y�<L�I[l;��F�^sŋ�I׻��n<�k�S�@n{��@�p��k�����X>�A�o)
7]�1#Dm>\�������'�G��ծ�IQs+��ļ���=�@���&�@|Qn��� �'T�/*aqRH�#Ј���Z�L7Ȇ.ڂ0��H�f��]IQ/!���؆����僼�c���je�x`+0�\'O|�ӼK(�j�߄qO�7U�cԄ�������E�]���5�g5!�H�p�h�"�L*АmA�NE�2P諒ি]|��֘�V�Cl�k����O���'�i��?����_�P�	�9�k������Ҝ��<�����afcl��ȁ؄<i)�� ��+��n�$��Wi)���8�dAQ��ެvӅuI2���&g��e�m��\�;Q����p� ���4R,?�7]�l$s�n}�{r�J`v�;��hh�b)���1+g8��A!�!j&���7��NxG�BsF�`�3�}A\T�J'Iq�P?K$0Ak�Cnum�s�ci#en��up�?���L�κ��0��t$&�pI�^�83�@�_Ƅ�","l�ۼ�Cf�x�L��{�u�2@���:팮�˿s"a<����	���D�"=��֘��v�z�K�����[ -�'�g�_>9<��#��8o�Q_�5����/kM=��M��U?��JF�ސ(�4�_�̭8/O�I�\X���뚃LP�d]�Eۡ�聘5��||��}� ��
�����t����9A�15��W�J��<������Z����.%Q��J�f�:��	���%�4#��)��Q_A&���r�Gfwd���i��-������>�V�����q���~�}��pm*�ې7Ɯ�`*�^d�6o��YI�pS�֟Y���ŕPmGP����~ɘ|_K\Bh��l�9��\����fy^8���Z�>������`��,>�!�'*d����?���n��rDWG���΢֓��H��rj�79R�P�*��~)�(au�X�-2iLT�����ʖ��Y|��1��ݚi�p��w�����s�$
���o���"V�+u�����.�x�k9
Jgݮ���Т'��A�;��M��tץ:�K�:�#0�\P��u��6,+�:�IA�fF�@v�f.RCt�G�"��ơ�ފ��n}X�J �}�<cW�.���ƶ�V��goҰ��ZD%V�!�����(�S�]`w!�ň������������8�N*�4��u���N�v��~�aR��\|�;f��ƣ�_�n;T�da?y��~o<;�?�'������	�*XÜ�����$��$g(񴠆W�~*��^�Ǿ	 l$694&��l��m����a�e������?d�t}/X
�����Z��E�=�_��5*�|Apiʄ��$�����9���ߦ�F����Y#1F.�%}�A�|�Sڊ���奴]rcJ7�]1�d��lj�R�uC]�:�P��L�����rg�ȢVv�|P}��st��A(�=G��x�v�6��seiF�P���cp����L��ࡢ�L0�XU�+I�Ȏ��[�� �d&��Ao��f��"V��o{�>vd"4�c�1�! y�r�C�t��lQ2�t��7�������H�f���o��d�'�\f��7������é^.
yK 7J�A�N+���y��))J}�	�
Cf�*�a�X���ܚ���~���À)_����: dIR�F��Z��������b%�Ye|A7(_�K �O��<t!��H�<l~���1+՞["����P^�&4�Xj���xR�,NsC�m�c���+x�{W�n��!\�#�T�&AJ��~i/!Q!�F8�.���)���6�A��F��M��2]P{�&���s���ފ�"�.�5�$�͆J���;8��;�5Zu!��n/��b9�R���d(�x�f�d1׹�tXļ��I�_��\��j�`<�C&����l�Ý�=`���xz�k���P��P�t��%���Gl������,���rBow��0��,;���-�b�W's��&��7V�&�s�"�鍥����N��P��!����\�J�yz_���'y3>�ͮ��L�x�ܘX΢��P��.Y����Z��Efߤ���Dp8ǧ߀�5���c��U�]d!�N]�X���X�YaD�S~�p
��4o�dv�I;�KU�}xE�5;[����U
�+d-���74�/��S����y�9b�\���y�E����.
(c���y	�6�K�rſ�9�K�H+"�������F>�p;�`���tN�Ax��um���Mٿ���DA��X�H�T`���<��x&^���]ųC�T��XXl���~�P�?�WW��xLQдw�$�,��'�q�0�v63 f�j��A���b��]��F�ሆ��'Q&���֡��05oNI��]�����
\�"l�5���]�����F�-�p�m���ĵ�;ȵ��<��� �g�l�L@�Hf7�c!#y4#}9�'->���hDWy��-��i�H�[��Gs]��_}����?
\��w���V!�����EB{F�֥�%�!u�*����&Ε3yrMk:��R���SyU����`��W%�4o���q�Ք���p��]�9�bMrbr��s���cX
pZ`�3���w�ʐ��.2!�s=�N#�'���T��Tu�\��?������YZ�|��jQP����ǽ��g+��>wd��<@���_Buql���u6=���=�����~�B�I�W���f5{/`̙��q����]�[�q5#�|aC�O�%Z�ZM1��$�j�WG� ��R+���+�?	�CЏ�a��,����^~�����0AC�HAc��C���	��-h�l�=.����!n�> d���@.m��:/��jj�xv<�n�jl�cf~�ۅ����}�7yÒ��9�Y:�aj��23���䑄/4����4���i|u]k�=C!�z�=V��*�=���ZM�:P��mQ�!�@�]Hij<篛𛌦"�6�GW2�b����Q�g�������<�:���{7����#�sׯ46��q沥џ��y`��õ�:�+np�����Rk����7RY�Jì>�,(�	!�~��\�cۄ?����C��Ǳ�.N
�lJ�.5g�) Ww'x^���y�����Q��5Ol��.FC�A.=���E��h#,(r�z��d��1���a��c*ɶ�
�t�<�}0;��4$A�	�z�D'��@����'��4���LUTç�v7�6X�����`�|�Jm �� �'��5�\bI0u�G��B��ٷ��VU_������U�X���Rl���~����M�2��1W�`)��[��8��G�d�87N�^�y(�ȼ�]��g�G��#�Γ�<���mf�Dɝ;��?�(zb@ǈpKm~oI�.��7o#Ɲ���iӗr��\:����)9A�����35��F7je�b��lw��y��b�u;�����R�1'�jm�1�c�:������65?~e>NJK"]չ~��IKǀa���F�q�r�����ͰQ�׹,��!?�]���8�D�2d��Yr �[w� tV�Rb~;%̻S�`
�(��v���U�Mt%c^�V�T��ߙ1z��^j����!hO�������?�S�B�8�0_/�_I�ayf�^�۩u_ǲ@7�����x���M�Z�Hm����ř�$"�È�ZL�]&Y��I�R_�:9ў䯋OL�"�ѻo~��6~�B���V�N'��2��~fp&�(����k�� ���y��J�Bc����(OX��נT١E\'�4
�2�����u)�G��؇�`�S(�>������d!�5OZb������EvZ�&��^i���@'�(�
v,\�C���0áAչ�-�����&�[��NB��t-�*�3MC,��W��D��b#t�ʭ�<]j��;8��&�NńO��$%�Nu%3��]�q�[�-Vc�i��ѓOO%��IIxZi*SՌ��ر)��6��e�r<X�GT�x�������x <���J�𲻘��*i�����E�eF����#�*����JPΑ�����o�x^`�Щ�|�(���$f	kM~�֗�'�Ԩ�5��x����R��b��&%�����!!�u:�Bϒ����2���"6��$?ĸ<�>O�ð�1��ϝ�lN��b���]C^q�iO}_��]�gJ�
4�Ӻs���>I���7�^Q
n';r�s-�34��-,f4Ѫ��c���t�v�	[S�n�d	�3�B�k�ZL"���!��4̘��̄慙Qwl�1=�_�ֱ��o�絕WR�"�W�6y����sv�b��IK���Fp��r^�\r�3�f�)I0�J��^h��������{��;���`�����l��]y��T�fq�j��D΂WK��֛X��V�
3p��yT�-�P�P�@M�;j�	Vu��vV��{��k���?o���j�a����;qq(<I���A������\�L������C:���Q>/��&��\�Lv�o�0Ҥ��3��o���D�5�<|�}�Uف{CG@>'�B:��,O5c\�J���_:ʲl�L�x��̦����$]~��%$���R��t�З�#�H��qF�<��/k�Gp�ȔV��sW�؋���t[-������'�|B�!�Ah��8H��dr^�U	�)d�d�9�񾝡� _�hsUI�����#iY��k��ר�}ӱ�~�'��}^���s���}�-a2���Љ*��py����9!�<���hd�Oj�	�|#�ED͹u�	�EW��`9�6�ᵥ�g���Y�e��V�h.�@�ٜש
{�=���m��t�f��	 nO��R���z�L����O�Ã,�r98[5�#���VB+vi[:X;�`���I�!����/]E�����W�.t��U6���ҾI���)���ڛ�uozX�$A�}g=�s�'`�y��G��zd�P<|�xZ)tM�:��`!��6�߲�:J Pv��AR�ɋO$�`����i��sU�K�_��'��N�������Z��MƳR'Do8F�Z��8��ԃRl����W>RbMc��U���KrXS�t�P#�70)�O����D��F�'�,��I8�k�PS��p�C ����Z)�`Vw"!�X$,<!��WA������dE���L8ro�:L�Y[H��y�A"i�SdG������oy1xsp��:>�=w*S؏A��ٹהj$l��u���BhI$��+��>��zg\P_+���(�A}�"]eZ/e�=�z���jʠ��Rg8���ܖ�>�^H�<�v	�U��ә߼�����ܣO
�\YU�j�'�Q�k� �z��8Ƚ��v�$BP=�&/E��Ccĭ��F��Lf���=l�km����[��tO�O��y�_�œ�%@&�����[��FeuK!��@r��j>�!����v�Ə� �%��q#[��@�����i;�g�˙��R��\l�s)겮�_M�=N�z���g�D&0���ƍ��$�w�����A�\�!�Z�9e$蚼��e��
5RE\?�:]���?��Cwn���8	�{r>@�[K�S7S�����7�4 ǋ<C��S&9�8y8�.�(ّ������f���RS���fa7t�k����ی\I��F^��ݭ4L�nE�f'�j4����7����Ug"C��� u���E�4'%NBj����ر���M���fŃ��d��ھ���a6Od9O���C�j��#�&ݵ�)����tc�%����rg�/6�!l�������6d�Ӆ�4a!˩���n�D�Is@\���h��m�W�ttT��I��Ɓ	�b2R���.��9�;ĸ�񄀐���)�m�=�mg0�.��GHBUL�-���B'���i�(�/L4�l�QE��1?��E��[Ah0Hm��a��7Ĩ���)�:��L�*F�
�V�("���5�%����܈�C����	�X�Jb��ޱ}D����2�P�X|擝+P�;5-Oӣ�q�g��"̭��V9`��]�����&z�O��7M#>]K�*(��,%/�I��7��
�y4�g@q6-�}�V�k�	|< |[����v��,A}�
+��>T_��T��/B�vQ=����F�ci�n�/�.�t32;󵐟0k}��$�~��Nxe'�>Ɲd�4wC����3āE�1����e�7<��[@e5c�+-gEf�R��t�r��i��j�@^���7��k��F�hA��8�S��E`�ct`"�|>|��Q�;��l�!]���k[;=���j��^WS�<o��t?����0
B��
is�c"��U'�r/FY�`��A[ �=�͉�s�
����tpU�p�ԛ9?rqt��o\�Y��\ݓ���5�SO��lZѭ4��jY#K0�D����2������r��s�Ѫ�����$�xz.�`�1da%�l�y>��Ԋ��-��z�ݥ�U�N�Kp0��?�v��C|Vݍ�L����FU^���/ױM��1��h��������!�,�=�[�p���xOD�+�v�J�!ה���Sw���UTsy���ܳ�T���Xw>��ڙ~y�P�N���s����8���i�]�(8be#Q�|o���դ�;"�و��c���wlX+�[+���s�=%E�~�S�Ei�-lM��Yq�'R�[["�~�?���9KJY�)�ҡ:OP��Ԇ�#��'�^6ͻrT�pǒק�}8ϭЈ��0��i��?/ɪ���UPt����U�1�M_l�o�G�-�#B)��m,zKi�/m��#!Z;�.W��u�l16��"U8�^	���}l��	���}d�y<�ճ�J�辦l�+h'�{6�<���|9��WA��z�ݴm�uY����[f|����k�1������$��\5[�	ʙwͣD�� �� qe���#e��f����v�2�7eᔋU�Y�W��D���P��Q��{��}sh;���h�"
���Gjd�&�ڍP�!�xE,������h�I
��>jc2��B�>����0���;ɠm5��{�|�<7����+�&c_����o�)��a�{��톗W��g��-��אF�+�/�dD��@�)�j����D,U1����=Ö_ս��?�|E�P|��2��֚�
&���N����2ۇ�~ׂ�Zݻ��+��E�LcP'�	�Ԯtw.�X�4�E�]�Z1��yQ���Z�>������il��_Pԣ�MV��>��p�*�]�l�G��2�_�[�}�'��c�Y�}��+�Z_�ߏ�7��wu�@��`�J�?�Q�D���BBnH���h�a����3������*nsn3.���D�#���5�{�@��#�u�������F�d�� ;��0,)^2��,���=A�47pp=6P�`zZ�.��Y՟�g|�0��R2h�c{n��gJ�X���>�NI*�/�`� s���XV��%�]�cy�a���+�ڥiyx}�e��ݡLȑ� ���cD��C�D$��-��$����	}Q!L� m]��|"^�v�
�'��aDY��(%�}�ç`�oyl����K�؁���Te]���q�]:a���b� CK�}%���{�Ģ��RmR�M��?Mؘ�o�N�sO�j�W�u�4�j-o (l]����Qqx�Y�,����Qf�my�n	��]���d�}�e��ޒTjn+��8Z�/�Ճ]M�y��)���khY�E=���, 8gM3$敯��d�+ w|Y��q�qxLf��v-�PA%����A8x=c�LK�����n[����T����2���J��]~�[%�2m��w�GVJK!�N��	������9����=�EL�C��NA���=���a�ʾ��>�"l2<���(��2�[�R�,9b���bC��e�>ݮ��ӭ���=D�Yk�#ܝ���!��I��+9z�Cڎu� l�i���M5��@b=Gj�{����wD��Y����u%���Hb��߃ :��#�+*O�me�fi�d�JG�sn�SNk.��@Q�TK�ZW���DC&��?0������|��1�_�-	���ا�͈_��1f�7��PT�̫sr�xq�x��k$�B��(�����#&���x����C��|�%Y�#�6:F��u�0}��Jur`'~(׶��^���c�J�kq��u���ȭ�O�M+���pӔ�v	�����ޫ�X�}fE�׈�Q��l�j���O8�8�����;[���8�<�tf���=�C4��S�t]M��W�@���<�k�iϖ�J���L�c�0�_�0�i֋2�Mg��4J�;vۘ�_�߅њI9��_`���Oݓ�8�����ȑ�{���y�[�5�GXܰ`_Gg������t�;7�䔻�bLݞ��"�YN�7����>�����VUc�
��0Y��ױq�3�gQ���ϰ������<��O|�j'���6���P���"o;A�[�c.��u�=�J�";�}�#x�ǘ��4������½���p�I4Ǡa"z�E	:i��_.���j���y�DB���D:������_Lma$-I�=6j#�-{���N��ي�;�\ۅ�Cy2�$�{��5��%�8M��~^����r��C?��и=[�٠v��BSBW�q�e�JK�%@S�
�D[I�1��	�d�q��]�i��\c4 㛗N� �������M�as#�r�}���H�t������7�)��)�Ad���58��H;��")��U� W��c��y��箕�T�t�(\���16�J/K>�악�[�������[�?�҉x8��0�hX� 0�yW�i���D:���dJqs�������ʶ�('�� ��J_�	�X�3x��<�o����_6�_n�iB�_R�7�}��ܨ����8q�#���x<��m�E|�����I�A���G%ЬyH8u�6
s�t2�cgp8��nz^��Lpݚ5�c__p7����j�S����-�m�x����	k2a7��!S�'��_i�����rڙyu��Σ~���aX���fA  ��wA���$�b�r$2k��A=��f�ë1��k�v�@ꈀ��{��N�y��&;�W.�M�����1���Ý��:b�*��= ���+>UEK�Ҳ@�����ޚ�C��چ7}�$=��TwAܶ�S	��y��&� �������mc:Q�c��B��(�e71�Ј�߈���ȡ���,�9g����j�s*�\���i��zâk�!���;�7��J/{�~,A�!�m�*��b~s��'9���gw�>T�x!5@�a@�3Hg<枼$̈i_�E=7ke���)"�d�����J��c� �?������j}���`�)��잽��@��3=�n��"�w;S��
���uaU8:;q}5T]ﺹ\��E,�cf��%ʱ)h�T"����J4�d��`�G� P�Qڢzz���а���.�
\K�В����/��*�Ds��S���{B�t�q6F��8�k�E�(�������Ꮘ=�ȹc1���h��9��K�P���0�&��>b����5���o��`�@�X&�������KI?��
/��o0ԕi���{��}��Q:�[����;�[ᠷ���L���U�(���X�J��kh5W��un�R?�"*�V�6R0xl����{3 ��B"��at��ɀۗQp"r���+.�1��q(��A t{ѝ����j��K��m]bE,���a�A���E4;��� �AJX7������Pr��Q�ri�O.x�oH��]���(�#���e��5�`z�N�[��{���-2���5R���u�2VK�W"xH�*a�zy�}�!6<�k�R��:PqBX�T�ܔ��Z��i��1��՟tp|�����4��kPo}J�Ѕ}/�+I5����)�@�ҏŏ�χ��%J��	ڴ�)2��C�T�������lp$�X3���]��)D< ���ܧ0� ���*��\�e^ը���.�_G�Ha�E�Z��D �cӡ#�� ��B��-ZP�5>Gt4r�숥a�7���(�K<Eb��X�������VKQ���M|mu�qྪ�c��h���r������&I�Si��"�)�f��@�Az/<C+r3��l���a}{>1X���ןk��'r\�����z��>ď�)_�d����xa��**����աg�����zZ��SyJ��Q�-�[�> jN��D��vL(M�ڍ(��;������-��l��0p헽�$ٰ�A���Ng������:*w��D�dG��G*{��m�a�����L��G�_D�	���j[8^ #�b � G�/R����#!�S����fG(+Ɂ&ؕ�Iw�ꀶ����M������IG�y:u�����k��R?Ӧ�e��;kcQ@(_f������n{�&R��T6���;R(v�^��"�u��ی��1���\�sV'�ބ8\��'u��M��4�����P&]Y��%_��0�^>��P�\�̵��)7����e}>x్�me�S3��suE2���q�H�̊�d���:@��R�0A�֧	Q�M�g4}�߃Yc�Y�Y~�w�ٿꖳ��ARڛ���1�Tj��fCwWܐ?��-9�o5J}����wu[�ۅ�ՙ����J1ݺo��!F�W����/�������c�j4��ɒf��Rp2�~>��M��_k�L�=��S%����؝�������.��L^<�a��o:��t@�J�ֈr�r���e�^�yդCx1��@��w�r�/��w���z����m������֏�%%$8���|�ޠ��d�&��f�2��~&�>;���T�GQ2��7�ƫ)���8�nYrH�����f2��1�a�~1ʑ'�G���?�ʜ�Sj�Ш�`5�������\���@�~����@i�
X�z�A��0i�O��A[���=��ҪW\�7����a����l�5�R�L���e[ù��Ol��d�(���A<Q�CtL��=�4TמּW��<�x��'�-@��C_ϴ��6�I>a=��8��.|���R�Å�z���G�"��Dl�qp������VZ^��cB�4�t��3�����7f禤�Q�|��ӱ�by�����"�xF4>�FR� DE�Sa��w���8=g� �^>�#�
��	�¸_�� �N��3�[�2�Ű����<� '��)x�)ET�ٖ�Ł����ϣ��aaD-G��8���!����N���6�P8]�?���\��wY������NӜ�N���w�
:��j�2��S=�k'EYj���/�5�q���(֠���� �i#Z��'C�6?�.�r��7�Q�[.�v7�,�V�}�5���X�*`cq� #ي���גԕP�n�G5:����:�=.^h &���8d�t{�'@q�e/�f�+�F�H�>�\P�&�j�q� �]G�r��y�*s�4��Z���OK�.���g_u���%R{����ڈ�h����U?D�y>����g�uW� ��AlΠ?,�fnok'v�{^	T��[�����&'CٙĞ�@a��.C��j���+��K��ɾ��)Z��O���O-�<���b�v}O[�	3<�.-W1O-�%8`�v��B�]@����$↪!7l�VFc��9�w��t}f�O'?�	M�?�+_ɊcDһ�k��;2�2@�2��鱏���Sm����� �9��
}<�	�R��J-����v��a�;���u���O	�{�GDC����[�� Ũّgv�%H0ޒ�'��O�t���F���5^��S�x��@�9��(�]�b�0j�.T��U��9w�Uѹ[�K�,
�����P���H�$�,��Pٶ�X�%�������%�[�zV�
V�s}�8�W{�-^JAѴv_�n<p�lp�fk�����v��t�M�=��"Z�M�$i��^����ï��U��&���uS��ctq�2ϣJOأ��p��j���O/��9L�1���/��H��ڮȺ.�<0K֜4_c��*�.�x����:鳘�׽)���2IM��\�i�K���Si��mC��,�h�Q]�wz�!tV���W������ti팭,z�|`J�ѿ�H@�,	�!&W�f�u/��۞��]m��ܹ��$�\�aQ��(J��Gþ8���fI�T�bY�]�Yb�.8�`6�Ɣ�1����ʜ�yH��L�/�.�=4�ʂ�+sU��ύdĚr���cŖ6�����={	6(�7������y�y���ޢ�D#BN��YU��,��,'_��"=2�s���.�;�\�W���pb�$�cڊ� �V���;,��-u�	Oŀ����d+�� �Y+�Ǝ�Pf���[�}y���Q�,\�H��37��o��c�2p��< ^|m�.��C�`�z��K����pY�er �4���9C�wU×�R;�{�(�H��:��Jq������ޅ�ų�e]u�<��<@�[�>��l��;Ț�@�����6�(k�� j�gHr�ar�b0����qԵ���7�,����-����>�Z ��C��A�`{�R����Q'Q�ٰ)�-DlH(��XEh]PKt�w�B���1{6��۴}�E�/ٞ��Tw���#��R��w;���<ˠ�t�D�bHG<0Dg��MK�H?3��4�쎮��N�+@�A-l삊��(L�._�(j]�[�����\�BiB�%��X�B&p�z�  ΅� �K!{5�+B���~���{lw�4e�l!y<���:%R�3A�bzI�����L����bMp�����M��)ưqG�,~� �fi���ݟYzi�R/�ԩɐ���ۉ?g1�K6�H�6���u�y�X���p� ��~ڮn��|�{a[���6�xD֮�_.
��-��-��mr��� �氼�sW!Ձ@�$z,����h.��	��r�̈́ֱ��Z!U \|T~��Bx�er�.�S#�p�v�<�
���j�]�`�0>{�a�b}$4Y����p��Q�D�<��LIҚO�M:&|���Z�j��WFNEZ��0�l���8�]�T��S�~�mhBv�;�b���c�IF�>^E!F��ab�iH�U���)D���7 Rp�{��`�\L��j��h�"��v�����L��߀�f���)�V���	��d5-Q�{�"����t۟Bx��\�O��!�A�	�ϊ�@!��3[k�Re���Wp�x�	JOAԔ�x%��!/j��%�U#w#?:sL,���J�.'
C����j����U\�fI� 杼@�m�^�E�1��-���s#O�J�O�d<~Zi�ȿ���T d|=�6�{�9�Z[���`p5f����<���?m����fǨ�}� �[�+�y�)k%����ve�B�z(n�i��B����r�Ɲri~KE�(J`����ɵ�v�Nʞ?Z�L��&G������Wg��آ�	��sg�N���!���v�FCv.U�=��lo�I�t^iG5�;T�ns��/�E��3�B�Ȩ����½��BVH1D�������v�)O'B`F��xZ_,�;���/�:��?x.<�����6�<Ttk�]�.�^m<��Z�����a��xɊ�~O'�D6�+�5"S�l�4���q���M!OO	i�����/��u�ܦ�K�h��