��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�`�Hӧ��W��u�?a7��D�7Pbɲ8H���%�k�W"q:��A�'��{��Wq9�ѝǥ{0����H�8y/����dl��L��-<hwn�E�P�9��M?$<������*�����͟ZP���r����֗���Y�0��>�7�Il��[\#y�0)�`�!����0,}�(�I�2�P���	5�U��m~�g����9S��"���� ^��153/���j*7��:RW!��
o?��Da��)��"��ҍE�ǆ�.mx����m��t\r(����e�u��z4CHQ��B:@O+;�uyO�3�G����\�̀���;����7� �gz7���jR��(B ��h�jlwXP�C-F"E+z�Ԗ��倸IS"G$�Y.	�Rc%��]���j@����U"I�#E_��9C?�[��US����<�3�0Z��m,��? ut1���l�Q$H��x>@`iy�R��ζx*
���j�}�{�pэJ��a�����3J%Rz��{�|BZ�z����`s���XZ=���d�~��w�5���-/nf=��pj�Fż(QLKڳ�]8çy��dc�;DN�S��X3�Q��L����B�9}[&��Hz�%���e%�ό�c���=1�.~*E��\{���OG�k���W�&�� ���ug@#ɪڃ�{��^����~�Q�м#?����l>3O��_�dnm�N�����8��XbOV�M���W��:�
R���6��蠢5nQ�g/b�;۝�N�@�/��%���*s:��t���P>��b�[�&a-}��6Z�1��GH>�y�P%��B7�z��7���XW�Ϭn�oy��0��60�9�+��fw����I]X*���N޴;�d��YB��W�g�P���c���i5�,��J�����<͒����
߲��4Uӽ�IC�𻷰�mC�=F�#�v��o�Ų[��܀.o�-a�ܵ=��ƥвonk����p>��$�+ɝ�'C8uhZ]�L��p9�:�����gLXi�S�*����j?6� ��/@q�����XIl�e��*��K�cPy�.$�j-��VP���؏$X(�Cm
vX1q��*�Ȍ��1�k�t��	�_���@��10Ϣ�&U#CS"�x�\�h$����k�%pN�7��I=��:���1~���u:��R�'��	y`nrn~��"K��x���z
�����!���,u�}ĥ�P����о[P�'�b��D��c�r�\̊���Z��A�� �W�N�:��J��@��r=�c0�z�~���� !hi��ګo�%��~Uԓ�$IN+�>�諟Գ�Ͷ�P6��^R��j����I��Dk��}䖵�Quv<��iKIN��"q?��6A����\'ߙ��s��J�1ǈH�.5�w�G��kĆ|}� 3�q@dr�G�g��0����q�6iN]���q�h�'\������gS]@i�06�P�0��:��3Į&�c��B>��d��n���D�5zͶڕy{����HqݖC?��0~�$�4�w�[=�R/\��f"��NUkĿ���=4�D�b�*7����V�����+�'�~&<�E��9� �,�֤��^��P"e��ힹ.�^����da�_	IK�F��⃚}�`>,�
R�*.7��2#�R�"��:
b[L�e/�W9�U�9 ��ݿ'pg��@y倁h�t[��������5zG�#p�~���J�%<�-{�L�c��x�\�I m�ݳ���(���.�8₣�hKx��^��0�{�;�@�?�GA�u�n@Y�[��@A�V,x�F:g���n׃��G+#�7��kR�a�tG���;N,&AN=���m�J���t
��9�=��{�nf-$>��ߔ�i�����|��W�������f�>o��} �����Ynx#,å))1u����%j�sϗN�[�s+#�>+��Ɖt�f��HЊ〕������������mj�����ٮJ�L��bb�� �)b ��[g��X��	���b��e�:���}U��A��������YI�
�nd����N��:�	����6
z�l���_z�05��?�H��K���}��D�(ߐ�A�0��c���*{8m�C�HWO����dt��iÍ���� D��>�e��2&^�+���Zo���V3����c�~��RkU-������.����)��4uK�@�[��Ɖ���U#8�b�<��"��,���Ya�H�&q:�	U��8��b%Ik���:��F$8��vZ���f�l�C/�!j�fu'�Mȑ�G"*�429Ir����Y�v�>*�O������?���k8��@�@dV�݂�;�T6�ʶ�!p�2*Cd��I�F{���^tj�#���Ԓ��r鳤�=ϣ���B|�~t�h,p���Y���"�t�U�)뙍�9�'E0�z��4M�kbf��
%���]����ohCS8����kJA!����]�w���a��A6���������8u����l�T���&]�\B|4fI�[z��?�c��A��O��v̋�J��徲��u�Y�j��qV�i�G���z��.K�&�� ��X$�2��[�\7�!�>u������]ao�u������������9�'�^:���f �G�q_N���J�s� �����MF�K���ց7�R� n4�-�GR�f+�*�J�5����i0Ԅ�Ƒ�r�Y������9���Vd�
��'�$7���9�>2e��9��I0!����S�g��R �C#�����&��y��y��Qԣc-�g�)��,#����6��;�u7���gg:��q�yX��E���
C?���A-���ۿ����5��!�8�o��B�G�-xud|''�DV9�������Or�Zq��K�M�u���,�ۜs������5K�[����M6�i&��7�Χ�ޭ���V�%�TS� FC�����uH�7H��M��J���٭Ye�
b���/�C��)6�m�C��F\�F�3��3W�u���lv#G���И�Q4���L��9�Mh��g;9
[t>����%�������;�f2έ�O�:/�K>����SW;�����y�|k/���ߣ��j1�In��t���H�`�9�ݨ�׶�}-.r �f��!�s� ET�
���G8�Q���ໆ��#�r��_q��f7�|�z�:�����]���l���� 5�%�W���?ɞ^I���GC��=�dT4��y����	o��T�zy���S�{q#8�{+{;1Е:/�b���EsyV ý�G$ ������\���a�LQ����dRk=V�����V��QX[�K�9�`�bR��ߵ�Ý,�t_-_���Ʀ�TO���^p���x�tw�#N��-�u-,gZC���l}�;%%�'-�oPF�4�M�c���y���"����u��2���V��V��� |��ʾO�I[�.�>j�}�]��Hyp|���K�,G���Q�\����}�s<�G͢�U�p�����6;�����E�z�*V�,�t0_��FO���6�b�Yv��dBa��E�~���bC\M�ɸ�q+���@TNFے��"��IՁ���3A }�+f�ߌ�c�T�H����5���v�P�tJvJ^��o]�t�x!��h��|y��i�
�P N�$Y/��nh��x1�>O��)+�Zm�3�]�˨����ma�_�>X�A�]9j�K��v�?�2��Z�����[���ֈ�K��uФ;�f)�&���l���g)&��%q���kP���>�H6��Y��t��wkH���sm�c��I�������yo!�پ1���M;��K�*P���_�h�2�-vi���#p"4���G�wi��s�DF���g�2��ÛX"��;bI&�u@�\���ەm ��DmV�ɦ��O��=is%pށ��2�5��v�5L�&F����k6п[i�u�<�� �~�,�q� ��j/ˈ���}[D�����ݎ$3�77xO~�?(��g��f�4?�7�q��d��a���{gz:����dW՞{���}c���;@��٠=�`5�[O��&ֶN������+F�Ag�g�9f�®��_X�#�#ʢ���-�$.���!�7k�܊E(�r���NiYk+_�n�����Jb4�I���|��i�|� ����CStw���[�%���]�$��l&zn����	C=[���yӧ��ɝ!n�:�A� L5<���e^�E�R);9�xù�W�%{�}�Ĩ��_8� �YR}\Ha(�f?�D�&'i�}G�R@���_;-��P����g�	��!���&�/Y�~�q�f��AA��o09�2�6����"= �?MNE�2 ��ީ����cgIz��+&I+�e���>��ֹ�u�'?���!�y���OT�+�f���f���
1xu�#}b�3k6�QM�[��}dg<���(�_<+���V�q���Z~�/֧1�x�؂�->�y҈;�o�o�:(Vrd!7�>��:ḳQ2�hN8�i���!=\/�7��ĝ�P���- ?E�U�1"U�7�G�%?����f.u��Pظ�M~����!�H��S�����&d�AA�4*�v�X�d���Ć��B�Nx��-p�=F4�?s�d_ӲJ�2H���z8c0$$�NJʮl����g&�t"�
�/%=���&6�ʙA$��+&�����A��Q21Vw�*9�13I�.�B(��aNm��)2�����/��ښa�:r/=5Ƚ��'.�g��-�.�����g�RF�H_.��Z���C Vu*���@5�Vġ�ݫ7�Z��dR��3l�9�
�R�H�����%�?o]�̎j��V^�ȗ)]�[ReAgֲ ����J��y�1,=����W�0���p���q���Ó��hD	~u�r
J����\���㇨�?Mb�%x+�w��#m��+���¨���X��%�z{鄾R
�}8���9I�;@�h�*��y�t���I\Y��?�Z��AL��,f������>j�.���6�f���o�z����CCM @��:���V��ݩVMw��A!��z���/m��a{����Hɠ�\����4�p�#�t��!�Ls �\Q�x�H{���{��WD��7Rn���&`l��ιy����Tq+�:�S��@1���П���><��Jo�Cr�e#C�s�����z6(To\"�\tL�[���B��<y�}e�A�9&,��=_j����0�54�}帮�)�5�d:�0���.Q�R�� kY���0O�U5���:&,߻_��k�m7i�S�q"v�ZQp�!%|�\i`#C����X��p�<��r��9�M��Dl\�e}�g`���������ǌ��#�E��TR�Ŀ��\d��& z��Yf�E���#򣜺�o��~����B�L��;;j��>��Pl.ܧ,o����Խ�;;Ҽ��/à@��p��A�$+�O&�t���W�Qn;�'��5�X��M�NI|!p��y�2	F����b�gG-f!X=S���Q6�+:*~	����B1�I�[4�' &ےV�G��
�����^�N}��W���N��J��~F�����k=A�[?Ŀ$��{������1�����%�������*ТW�.`�JyG�-����s�ve2�v�*P�zU"l_'7$��~��}/�/��N�a�,P�U�X����v_�T`�@"�K�����Ɨ�Y`���!�0������J>�&�D�G�8Nze {vE���j�s���`2]�q���$����4#�H}˭��/��T��?���1��c�_�������3Յ���Ќ2p�٪TWD���S�u/m�tؒ	S�����[����H�����`�� �V0"���|���4��h�b=+D����ۊh��O����5�,�t�`֙�Q1��߳����b�-����e���������>�!�Mh�z7\OH�RQ�ٹ�_s�/O�ś�0�`�j4�֯�p�3���#�셡�L%�qf�؝��s�s�$�*;>Z��s����OD�CL�N�kj���\��-���\��AZ�|��3�B&�|�d���9�W�k�a���R���N�,L����
uv�ύ��s���w����o9 HZ�g��uA�z.x��׎w�k���'C���}`�c��`�)5[4��Bл��>	�9Y�n��k���:��
�{G�&���1�{�9�z���m;�.-������੗@��� A��G0���9�,�?��1��	C߅f���'-Bm�M�v0��K�y@�]A�(dB�	��)qa�i�
�� �9^��1(�|9���vmp��eX�Ph�NG�$�,@3te#��wq�G{�-��U��Sϫ[�O�^<��Q;a��7Z!U������tL6>}��n���X��$�o%���"�y7�\�Màq�]C�yu��d+%lH����<��3^D�Ze�j��i�L�e���E�۠��/�¥�s��-(8@W���z�L.D߸9p*���yT��8���#C|�Sb��ѱ9��xC���*J>�1ns		kVP��\���W�;��Ds�2&��DQ���  ��y����b��lӵ�/_2mL2���Bq�v�"ʥo��v��o&m���,�a�b��H��"A����q��ӠIiǍ�� E;H��~L"`ܥzj�!��u��f���-�$����Tq5�BP�xr�ǂ~j�R��<��vm؟��Fɵv��L����O1�O���:!��F���+N�����ϐʹ�� ��kd�dvUE��˵��d�͏�dx�
_@�"���Ś�cZ�C�����}�<됍�.E��/YxN>���%��y�=Xy�A�o����b���N�	�P����HӾ�x��_�F�^d�Ƕ�A��fd�#�ܻ�6޼���zK�*�D6�A�s�#,�Bؠ�̊��p݋�%��6�G����=�8ɐ����:�6�(TȬ+:N&7`�r{�>oyP����D�cB��9�J̅�E�[�e�:�<td�s�K��绫
��1�����-�a�caR�؜g|�w��@��=˟%�_�ѐ��&���'M�(P�wu�/lk_�-�;{�F��-��:K�=��C�s��J�#�?5V;�Im�Nu_�:�Jj9*�xd�&�O��^��.��0�6anUܠ��ܢ#n�~�uG���,e��:`�������Io�C}���{�>�2�B�R(������5o��zJ�t����W�B�D����l�2�X�K����H�h;O9c�p֜?U�I A����id�?�� ڪ���X%���S�|���k���k����`
�x�!�_��/��k������Ϟ$2��j��h�?�r�2rN>���?ŷ�Q��:�-"ѫ��g]49�=���F��C�7/[6>Lgu�
�F�&a�����lTc�y�x#v���}���� ,w%fD�4����|�T�F	�*�1��21�h*���.ğ�<�X�A�Lf=z�����xz7Y.�x�U��LQ��g���ne�qzeg$�!�2V\zش5�K�qd����ژ��ǯ������!���R�+U44N;4l���3�:�r��I-3֏^2�%��ؚ\���������]�A:M���j�E��j�χQm7b�^ڴPY��<�f����]�ֹ�1�C+nM�Py��j�\�ۋ�mW���^�Њk���X�_�+�?T՛;�֛��>��;�7��I�<��xy]�+�o
V6W��h�w�u�	XJ�R?�<���-K~c�J��iQ�HZ�R�?������ީ��+�@4zt0 C�V�C�,��q���z	-a6Y���#/�-I�r?k��;c�+�З�H�-:��Gn��ۘ�y���؏~�W\5�#�{7VF�|���"v��	�I������(տ �H{�K?�ư2$"i�eW]�[�z~�z�g�vS]p<e��"��*����0�ɣ���`�"e>�QO����+;6�?M�+�`o��O���J�Ey��p�
��3��/ة����Y+a�i.�On='��J��>0��%�ꤒ���>�(�ehl��?�g��J�ϗ�R8���u1�x�Kb�x���O��C'�'�O�ޕ��2��@0�D�d��[���4� �2�����Cu�O�Q'_�h����9'�_��خ�2}�~��
׾=�DA���	�p7��o4�7�g��bg�%)Umϻ��Ɨ�:�M��ha��aR�9��a��H�6���V	h\�-���|&6͡§�<��y���ߖ����m��C�^U<m��g��������l���j9N�ݷ���D�)I2�ܫޡ���
ƭ�N�����ΰ�}�n�a�e{&)���	��-������`�(*���綛�!�	�)vX}��M�9+2�F.�W3	��b�TS��{E�2�6m,��3X�ݛ+��D�K�3����PH���w���S��H�w�e�zt�ɯ�P}��(΄��.IM,�L44���n��D�"�7#A�=:]��?�"{k\���ԨL�i�h��nWNpK!
y���b��^& Fx)�D[�=R�B/ǲ^<�a�G�5ר.����J��$�+�0��P�^��>^�e'b��(�J���8��Ӳ����`��Ddq.h��4�H�wp�	͒4pܥ́���[,W~Jo�;Q������2rm��䳰����V^mBE�#����u0�C$.]�a&N���,�q'T@H����`v�l`�MP	+�Z������� �dPmd�;�ר4a)�ɱI���T.ɂ&��n�Rw�C�P���D���[����<8��A� C];��hƨl8=%���|�hiJN�{�z��Ð������@�{���[+W&��	�}Q��~4`O^?��9VyC��ސ�t"�Ϡ@�2�,|z�7Z`��U�A��lk�������+U���,v��{PY*޿��c?��eG�����ʼ�.�!�ڟ���r η��D�]gHd�<|�h1�Zb[���㯮+���pr,8ޚ��!�4[�d���1����p3EP�Y�1���e�S�[H��r�� �!I<��37�J��0���k��u�[VP'y%�F�ca�F�>�|����.�6dξ�����S����D_i�	(���;nF�qX�[�bXsQ`zC��V�w�V(11�����'�펟(i�����P0�8`04K��׃��sQ��=���ҝ眾q�`��P������� �� ��Q�k��ڍh����)k���;!z9�b�2����3|�iq
�d�9�5SU_@�Z]U �a���@�뜝I��ǋU+� .BT�*�D��-|�1�?+o��m�<+n1ч�4��OvAi8����Oo�OW�s��p �ݴN�S��I��Ad��	���f���hF���@�����f��˶sZ0+���T ں�P��ר����0p��q�+[�1S�?�)�֍iu���l�2O��l�ocZ5
��Z
�l���G�2I:��"[���̹{[5�/��C�hb�
���=ԏ�� .\���"�(�������N�(̖�
u.�=��?�e��� #�����a���l�gU�J-G��.�!�n��uD����5q���.y��.�Wd����^�v&�ъ
�L�����n\��Ɨ}Y�p��:F��H˝ �vm�������~��s�8yҠ=�:�����Q�sv�]���h�}a��t�����J =������qAQɇL��w8�y���Cz��'� �n�$J|;�Ӄq#0���5��Z��e�@�T�.�Ӹ�|û�԰f�:�3:rU��+�lֻ��	�*�v>����I6N�'���@�j�2+mL����8����*�t%�zM�I<�� �N���!�Β�D'
���Ƨ��ꃙ�"�&S.iYE���b$qnu�-Z��Ĵ3"�0�O6%kۍ5�
8SS��;H�啻u� � �!]~�ޠ�Ci�f4n���c�ƍ#�!��s���C_Cӓ;+�8�����7P35Q��6��($�{�1�1�,��0��Յ�r����I�u)Ǣ�J2/�Ň[�>�۝|�>UCV���ɬF+�g3�G���� ���,.�7b�Re�5��zmA���EI+���\������!�3�d�1�#oR�R��x�6?��h�rp�{羮7�U �
��QJ��q=u��ʵ��+��G�af<�	��@4J]=�2��E�&̇!�RA���}0��VH��� u��([���?�v�h?;��e-#<e6�P�����l�l���97�
��8䇢�,Uܔ�6����N!�k�E��ZF���Q8��k���E�5�A��;wlL�-/B�d��a�aRIiK���e��E����s�=d�.� n�үi{$����t�=ۑH�g�,�9����N:��z�=a�.Z�z�,W�5AQav4��y� s�c��`�ꢆH���_�ɇ�=�@�,Fb�? c"ȓ �ݢ@1V���l���� J�u�鱗�*�A��<a<���[��H�FE�wbV�1aٔ����!Nt�abN�l���rrW�7���q\�_�k�N�̮��2�;���O}1hX�Fq�	�/$f2]a�Oʹ��E7'���}R�I5+�"�ؔ��������B�WxX�����`M��T�mk��I��y�zz�����z
�М�KY~)��G��������@%���O0(!q�.@`i@� X <\���|b����3aĖ���̄�ZXx���ۭ���@��@��G��������Q�!
) �[����9��,M $ ��#sFw����zw.�ɐZ�@ܼ]��p�0%Ҋ���?Sr=s�,�Z����a��Q8׫���ۡ!�����[]HY���?c�����i΂%K��tf
ޣϦ�]{�Ì(?��L�ή�;)^�_���Z����L}����Z=e�j�0���4��ī�:����!�� ����ت�ph���f��:��НUR��T�+,Ɯ���i�l����������C0Q���	��*˲��e�?uO�3�-���M�@4G~��EA_��L���?�Moh�_�u���jK��Ɨ YU{9ڸ�����C��f�:�]�1Ɯޝ:�@�l���2����Q� .�u�	}�9��K������Z �S�����pCO6�Z:r9�o�<�WE����łu�����@\(Px�p�ǕohY~���pu ��A��\���8y�qPD%j,i��({Y�{"�CAES!�d�C�c#�A�@�37�����4==F�}�[b����-��@XM���x yI�F/A1Ѥ�������]#�1@�7��C�t���p6V�$���!���{�z�	"hԛ=}��� ��ޫ�7���~����
����A*͚�nol�}��b嚐��ػ#No9ˣ3I�/�Vm{F|\?�(��<G��V\���?��p4�b�S�o�nL�����rN3ay�"�j��C#4ZB���gdP�Й�ǜ�8�t
[!\F�kI>�.�`�U �	�\��k2��͡I̆���B��`׷��������i@��
�nҍ�����>�6Cq�Ӹ� e��|�l��⸗C�<j<��U�������(SAeh��?��3�t���ߠ�j��ijށ��0'gl ?�g�X�n(p�I����-gd��<�fa--[X�z���;���-�^=k��U���4쀊9A�1hU�0<��2��tڨ�B`�ZA����^B�������Q�.�>�L�Իy���ô0�cE_�d���Ѱ������<*q2yf^z����]�u�.N3�|B���j�Fh#�/�g֣�tN�c Cs���<p�8L`~��D�=X�!��-���n�B� ��n^��,����D��ڸ+��P7|�iD `Sm����mPN�?�'�l(x�"��?�*�Y���O�O_uҙ��ΙحM�~9F!}R���\�vQb-���4�	6�k���YrqAg'�F��������B��<-D�܌����Ԡ̮��m�������_)\��\Z�P)���ހ��̗Gb���.<���_��SH���!����Q"ӑ�%N����S��?��
-%&'�pa���d��8:r��}"�c��������ʧ�ŉ�l�h�����'��>۠�n��ߦeI]r�z���)��?d)�/ԋR��V~�ѿK\/B�W�F�`.;��N6�-9���b����}�H�����
J+"���mn]}2�e~�^ٶ�h ���ȱG@��5�KCX��a�(w�TCo�ޝ~m�u�hG5���t��Nt���%l��FV�W���+�r���p��t�*�����x��X`P��s;�s׾>rv�{#p�!r�Wb�H&G��m9س��!���3HP�&+4�z
4(���ZJV�r7^��ڷ�cV�-��O!H�.v���V�㢬*����k�hlIb��:�8��qڳf��ut4m9T�@��TY�
4�׊� ��2�0ә�ڏ _�3�(csg	�ih��vFuV$�D��j���M]z�K���m��_�ۓ��R��u*���9TuW$<s:����^5��r�W�'�
2jQqQ��h�0�F'[r2�\���dxJ9DoB�6��a��ϋ&p������ۼ�/�E)���#9W����ib�Ʀ�Y�T]�9Q���+ꌔT&�U�&����-�~[�.zEx*.@@߻���I��r'O�hk5j�������*�@�l�ME�p)�ܾ�TC JB4��r�u��MsPFʺ<s���ߊz3$����v��~U�����e犩�
s���pD���S�1 K'))f؛�6���M[X���U�:x��� Vh�@���(}�^x~�[ceТ@)�{��N�:���xT~��sN�T�.Y�%H�i|�M�����t���}N��[�]u	L�I�#��8�'�ne�=�-U�+E� ��98;ļݸv�씠�R}��{��p��x�ɢ��:��:�{	�=��Ϣڪ9�<�h�wg��<��9 Gڧ&��nv�6py�b�5]`�*�J6�Yy�f�.�A�����\��R)"���V\��H�w�"XA������<]\�o����LK)�����v؝ٳGTj��_&�su�ׇç�U��#C�9Ikk$k�rւ�!�w���5�Dmre��z.�ϝt��H�[4ݏFUi�r&��@��|)8�mn|i	pl�8������P���Sn��NU��
%����Y��Y�yi�︄���`�2�;l�y}j�ˇ�
Oj6´
R�d%{�Jw��.�(��#.��T&d�oMQj���.��J���ڔ4O&��M�?����|�>R�}==�P|�A�g.w���2��6O
���l줶�ڥ8�N`���KB������Z�E� ?e�b��(���8*�tg�s]�W�+����SI��Z��~�p׿�$mnZ�L�Ĩ~�I��41�*٤�kA��ă.��v�v��y8K�a��O��`J�k��H�M_���'���̌ �⦯M�+*6D���W���լ>�gc�yU���^��a�NjF���꿥P�[I/���@�޶.�ɇv�oo���[/9�X�7������.�P�6�p��&��P�)�Ăpz,FsF|��Pff >�ElWl�K��X�J�TёT��/�E����S[�3���R��_X�5��3�Ϗ[t�0P:m/W-<_!�v�e�I����c���cÚ���ݫ���Tn��/f�q���_��a�o��߅3eQ�9���*HaV��)X��{��RSw��XU&��s�P2*~%F;6����w�!=���[�<~��z�U�tX�_�e����#F� b�3��>7��*��tgZ�[^�*V�Ν�I�B���<,�@�k�����;���%I��T��V纍t��ՀjM�+���X8g}9	H���M�hͮt��E^̄裂���`��X
�B%V�<��G1�`8�����W)e�3
$ �T��~�Hm���鍬���k��ֵ$H.5�8U�t�T!�G��������H��.�V�R��(漖O�ຩ������$�;�5>v��E�k|`,�*�t��m<�L)�ـ�^o�Hv5?@w[47
�f��.�t��w���'�nY��ᖢ����/���"�M+33�csk�+�(����9j`�b�#���SP2�$.��z�)��'�л�(3\���*u�����!&���� U��.e����
��4��f���]�?i��<�&�ƹE>�%N(ɅQJ��K�6��.छ���焄��-�I��b��ϖ恺�1���l]SK�b%��م�ǐ����3J�f�n��H$� �b���P�;�8?p�h�=��@G�EߗE�.H����;�,�_�^�~:��"����1�Q�a��F����o��n����l|�Q��P:U��Mmܸ�;�0���m�@O�cy��@q�����V]�n������bBD'�Tx!J�)�X��D~�;�D"Bڙ�`75�R(�{��ir�߮���w�~�6�V�q� ;>F�j�en�$����!ޝ"��DnL�J�0�H�/[V^Δ�7��]6�=(����נ2H�R�D�j�~k�X?l?TDv�zD����U����zc��+�8K$Y���������iT{�G�"�v�5�^˖�6��z�2!����^˙�lg�c���14����j��kz5�����NB���S�2@���ގ�M*�����x��3�.�	ũ*�9r"O�M0�lCZͽ�z/��;$�� �����v�m��zὰ����B&¹{j�&��.H�5��pJ�w�&�p{ED�my|��:!~��AL� `Ʋ��f��S
H/�u�g�Ʋy]a�2OI?Λ�N��`JO���^6L���OY�a�Z���ѷ/���L] "Ie.[���~3�.�r�Z�˴Hj]���j����L�x�V�~,}�����p����7��8%�q�r(�T@Y�xVT��a��򴱆��� 3@���$4!I4�Kj	�	oe妶"����q�&=����"�m���{=ɺt����0P���Ow3��E����P�\!B�y��BD�CU[��Iye�W��Yd��[�R��w�m+�I�V&�AC�G��� �6��*�R<��X�Uq�z�P����cz}��4�wĸS2G��Q.b'��n�Ҁs�' �M`�����nX�2��	� F�ElV1��&�h��#{��MN;@��
��?A�P��@�[�l�.����y�T��7\wAQd�ݽ4���l��q�K�=F$��=31��k��u.��.(�e`�'�c��^��ߙ? ��f�el��8����D(�ܰ04�a�_�B��H��H�-��;'
�x8�&�JZ�B¯%#*�{~���m_����=$�<mT�2k����H&���g�UAI_K���:��C!<A�Nw������qz�M���Pm+�ڕ�롚9��G3O��v�A�<r}aqd����#�'����3�E��K��ʕ��bc�t�ϷT@3+�|	|k���+���P	���3��w������;��
�
[�w��H��Ơ"�1Un�� 7Ihy�e�m�ug�{-1�����Q&�n�er�/���/�mCe蝦��'�zv�ufg?��ƞ�Y�j���Vr�0�<N�V|�9^�u��|��Q��E�(ql�.��0;�HI�M%��mCCQTћ^�u�\��ǔqxg�Z���r�������Z�⹍;^��ZT�HV�Y���\6���<(�ُ����w�U����/�P���v��Ӳ�L��Uac��)TO�6W���ŵ��4(��5i�c����>��(U���v�+*��Gl�Wֲ~��@0%��/J��G��&�vr3�-}Wgr����b��er���?��"Wj���b-�1���9��`}3-1.��5~�ےҐ]33�2Yz�C!	��pG��;&���C#]����Ik��}��=JW�F�6i�EӇ���7Z �ʕ9r^W�~���Ē��ZP�~uÃ�:X��]����=\��E�$�i�n弗b�h�������'O��\��k�㪝Hy��l��Y�,�:�-�c�D���w=�E�a���u}��Zb��Ʃ=U0�P�8�DaRM2�%�EyQ�Bjq�5����=]����(P�7��F]oo�;6�f73�ˤ$�;�i&��~�F�b����y��,�0g����/��^$5Yg ��m;�2
6�%�h�SX�f��o^���д���2Z����m�|������l�r����i�$�j�{�b_���4|Q�V��ryk�l$v�TgS������=64>�Ɓ�=MwBeW��:�x���Ќ���&D�+�GD[[Q*�qN��hg���H��~����z��Bw��턇�i#�<+���L���N�u�C#4ڲD�O�n��X?���Rc�#�S�IT�swTq�B+9Ti�@��"#U�|��4z���%𧮰��i�-<�ԝol��<9����i\�؝`��+�b�m�q[pT��h�ˆ�TѵS��6'pv��H0Uj����'��A��+h��왒>��y�N�������5��r�J�81�i����|y�ţ����&�L�����Q��	��?ՍB���`�3,��i�\ �}�܎bzM�aP�H,\tq�y�a�P���+`<�=���tJ&"������آ���ȕ�x����\d�E�5����j}!k6���Ы���h�!tM�ܯ�`�-��f��h�)���3d�B�G�@�S�O�Vj8]�9�����X�f�0q��(��sKH��d�|�����ZYq�!����j-t�EPv�JGV[��(�{oH�4PMR<点��_����;a�lm*���p�@���O(�v\\��*�ϧoAn����~w�F���}�誡��!5<K�N���N��r�%ŦJ2��@�i�S&K��x�O��Gm���	|����9:���hz�#�C	��������N��|��.a�Kv8�e[����1����L%#��k�3��`,���4�=��q�.Ūa̧�4�RHdwnn�~2@nǒ	9�(���%ȗ�q���H�7�V���D+T+��;Q��+v�_}���aL��E�y����?�b7�����̝M�p1���n�E�o#�֍���J�������N�]Ev�Q��"�^r�rhh�9�7a�e����}1b�I����l�:��I��8��q^K�TL �@D�x"~�NC����`c6﹃�������:ϕ.xq�
e)��ԋ��W��e�̹��M����A�<Z "5hG��6MV՛�Ҁ�y%�RjH�NkF0u�[�HH�O
��V�5RY���q�$�@�3�8�P�� (�MZ���`D�y{��EVSy� �ӔC.t��(��� ������}ն���a��b���B{�Y��L|�Wj�@\�0Tꦦ��%�)�z�w�
����̞�d]t�e��{����@M�g��b��ʡ�k)Y'�X����8P�ajZa���;���D	�!�A�K�Tx�ZF�`����ƼQ��I���ص�,]g��2�q |2��ͷ�gH���(b��-�~'���?p2���m��\�4�uܹ�r�k��"��P��?H��S�A& ��Ǫ�ڊ�zT��D\*��(������${���t�[��b��)����:�4�A�&��;�Y��'��^�ec��0z܊Fmw�m�dҸ�7��,�Р@ �������P6Z����3�S������ �êV5ȗ>��u4�x���7�3ߡ��FB��j%r~�}@"�`�U�O�BԪB.�⤴����2��*w|D4>���sb���2��5�2��b#�EE�%��I�j.t��X������}��ڔ" J���Atn�#��Au�g,x9�o�4)�Ƿ?����&�_�!��|Kؑ}�JFi�ww�5������(&��f��&	��س]a�`��_�f��Z����� ٚ۫��8�P��W�;N�g*��M��h2v������ţ-s�*�(�'�l���T�v=�Z"R={ҙ����0��<��`:F��_�1#n/�"[�ʶ���n&�r\G/��I _H�ꁝ���x�C���T8l�x���^��O4���`������M�-߸���H����_ε}�2��q��|�Ǌ?f��b**��M:%���F�T{]��_�1�1���սPȂM5d^/��]�Q�ʝ������c�`I�RBE�/ndC�"�ٖ&wd-�{@��zW���w�_�זk���>0{>���H\@�	�i?�o���U:�y���J��OZ"��Jbsr�2҅��6o��V=<�N�e�@\Q����-4�K�V��¿�H`bɋs	`��f�w��=ZO�dh�A�yM��R8^��û����jӕ�x���B������+���8���w�u��$���kH8�|��( ] �-%�Jy���*�J{�=#
c��D˽���ōeeX̲6�I��/��r��V��}�� ��ʤ4���V9�W�~=h.���vx'�0}���wJ\��Qy+�#�p�RHU(�&�&���z���e�ӌl�A{�.(�?	�/��6�j7��5�� �O's\�&��bG��w�ƯԌH��wbz� �xe��M��;&����N�U����1�g�WW�sȪ�[C5]Zw_گRZ��OG?$9n��Ű��qaF�[�9�o|>�n� ��+����cJ�os�z���r��y�]����R��6�(҉.2�;Xg��3U!ҕ�wRx��44=��.�p2z�n,{��8O�I��{�m�h�Q�߷�'�@���81z���}���?6g�\��v������\;�f��
�^"��aF� �f�B�?���2'�~{*�ζ�iz{�Lo�x��g�C����/�rLq�֊��Qg�MVh��~�K����`,C���3c,���oa!�)��haQ���>?�9Wթ�I�>��dl�D�̢��%�Hh百�t,N[�ߍ���NUj]m-qeW��X���_�>�-I��O�=�1H�,��^k���2��p|���R�X�]�����PG�_�Β'�v�\���,|,���I�`���
�����C�y���y���V?�}#�����l��7�8�⥝ߺ �|��O�wԉ�\=p�ax I�'J�e������o�������1��[�E	8�9�B�t��]��P��fs @�.QU<��M?vم��)a�S���wJ��'G�K��b8=H!F�Zכ�G<V6�o�#��������ȇ�y�����-C���w����)�D7�Iw�Lp�l�~�@��0��-	pK�����0����Zd�1����_i	_�Ą}!u���`<�����D�~��Ǵ�����E]*�x�Qw�z]�R.S�'2О�7��QG�=0\���`�WX�C�1X�0ߙٙ��Wsr�婋��R8��nW9����d�1SZ���cc�/���%a��̺�W<�L��][4�e1OhΣ�c,��m%S@;@�ϡ���t��k ��~�K򠩶#��\"����(IV)s�<(>��Z#����FTN��Pe=u�H;��M:���K�MZ�ê5��?��_�#Yݔ4�p���*�}o\�G� <sl?6�o��4�~�����`8N�\�T��x��-�	Mq]�>�u�������[]ns�n�� ����}���?�����P˶��N�5!�@ܟAw�m�o�V�tw�<w�XEA�9lI���4u ]��Ƿ����}�R��m�{�ӏ�e�M���҆"�ݜ��\S=�z	<]˅И���6���;W>E���³T��"X^�Ž���qS��u���D�c�k�y'{,����Q�QG5�:L��
�{!�0vg1���71砙�z��L3���˗�5"7��r��i�EH~��,<K���o��h�ni�4�g�M���;2�܋z� ��~�3���Ӂc��*�Q�^�nm��}��#4�j��Dăk�X��%,G,z7$i���z�6�;xV������V�6�TJ�!��4��#�i@�g'{�����_T19�[װ����Ր�u�Dnk	�3B����I|��
�_�E 2��y��2��἗�Q��C5�O�������w ��&3���MB�bO	���r=h���V���:�>����M$�rR���#����m��`�q��s�N����Y�P]h�ܥ��Fbg$>����V��,e����Ȩ�n�|N�k�����_ø�G��u/�$��N�5���^D����[�aIr"w��0�M����s�e�4��E�Q]��5��d�����j�cO�X���eR])r&��)�U�ЧGL7��]3*}Y|Ԩ)sق�lB�'�_X|`�o酌�CK� Ax+:�;�'�����ۖ�k �`S����`}�,XZP|h:y��=*�t�c��(e����e^�M�b���[�r��T~*k���`�AȾ���Gtך:;��w�I�W��!}Bvθ%X�:��Rי�����~f����E ���|�+@7�;�c���>D�\�8D^�37 e58.Ժ�~**1��~�Mq��|W�]{�H�I*�)Z�M/�
�bd�T�叜+�2�L��ԕ?�J�(��<��@e�a�Bv����ZKWBq�O-=4��W;�׍�Ue����ܾYDWVI ٳ�ψ�-/��*@���+H��"��G"���m�J����Ye
4�P]Za/U�ƿnHoŋUN/9�&�(ξk��ѫ`��*X�����\��q�B���hR�S����=�����ѫ���Lkr(@Kk�D��Pѝ�%���\J9�%��������N�n=$GU���9��aJ�D�@��s�aQ{F[�/�*����sE���^�2�m�(�Fd(V5&�6���sum��`E��xa��yd��%��C�VB<]?��4./Dc
㑐<��Ҕ��}�c���|��%��Ew��ǂ@nJs@\.�Jw]LW�	0W>Ҭ�r lN\-�s U��^��I|���:��=:B�V"��o�[!E�((��mg����:��Pf���ﵴ����-�l�Ӡ�����<�1�w�a6��g��Q��\�0����46����^
��"^F:p�U�0�'�Ol�!���jɣ�^�|�		�X�P-��5�#"F��XN߳t���b[���q&��ݷ0�ߋ��G*�:WQzq 3�pye��U�-w˞~�_�1R�<g�������w�#k?�bQT�#��u�ne�|��"؊�+�&��������zt�.{��i������B���6H�4ôթ���!у�� 7@Ax���`C�ʃ�8�����dO�Z�h�v��sT�t��u3:*��O^�(p;!)�a�VW�~���-,͢�xCI3�;��20Lּ�Am&�����5�oM7 7��{�z���[����:��8T�-Z��^��#�.�.<e�pón'���Xflvo�[}^���t,�	�9V;��=�c��{����8�7|����(D�ǿw5v���- 0��
V�G#�>(�M�^�y	F�q	�/��C�_��@�&�7�@eiw[A��B<�V���H�Toίq�˅�f������z>�LJ��F���6?-̿pf0���w<(�.���xx ��V�SBy�}t��gg��y�f�}/-�e�����z*_��WSoO��v�� ����i����C#>�(\_ޯsJ� ��+�:x!I�
�i�Ӌ�.c_�K8'��W �ih��B^l]���6�l�J��@Z�y���f]Q&Eo*G#��Z:�Db�@D.����fKY`��b�:z�}�i���Z��y^��~����N$��g�h��[�N�v����ܛָ��Y1K�c��f� ���;�� ��v��܊Xq��