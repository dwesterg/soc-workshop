��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�dj�x���W�9b	ߩ3��b�K���(��.(�8��5��a�f��Ҍ_����9.��;�Y{R�]5���2��3[�yՋ�iJ6-�^6�Q�u 3\|HC(� ��j�r{:���\�:�<T�	��4b;Π+�I���8�"��r(����$��T�f�~�rm=��S��� ����0��h�[�� �hu<���ˌ6�@��1�x�DP�Ga¯�ZwK<�]���FkM*�	�K�Px�?s��M�����~~<�s�HLD��(6�_�0�0�`@-o�^Y�j��<o��hs-o/=v
���8z���DK���i/R�z��5&�rS�HCZ2e��O��-Cs;��S��B`�0��a����/yȯ&0��-�����-"�t[�I5C�s,}� ����W�Q�~�]Uۓc���{�E�D=�A�I��=U:V6�+V�(7��>�k�ې[}^d�������Z,�Xh�|�M�\(՝�X���.�AZIk%�J"}�@j����(�̹�|�%QR9vT=��;\2����x������WZ ����"�T|�XPl�|�~7x��
nQ��M49oAD�q����y>/�.и�Y<1r�S�:��� a����M?�쳕Y����ׂg��<��@�ͩ�D�6�'(Ϙ��Pe�W��4��O�Xf���&A�8��q�ͅ�7�[�)[1e��{Kr~P?����ꯗ�U�A.�U^G��	e��:�䕎�����؎�`t�]�\~�4�ձ�g�tr�����kg(XT~�e�q�J r�>q|�"�]@�K�Lw{~�����N�ejdvW 
i킓C��tw��垂xA�0����m��V�$X�C�����}M�>�-��K�G�M��*~<��)��`XVZ;M����dt֠z<�zo} ۫[�=�x�yr����9@�#�{!*�eV	�;���\nL���2L���ኡ�����Es{�G�O�'y�8%���d�����`. C��cq���|��7T���o���:����iT�cSt��#zl��Ϡ���C�V�'�|.ސz���B����`��2����m&�:�v͝�ޟm�L�E?~�N�+M���B.&�����iBⶔ8�9��Z9.�Ì>[�\sښ1(�УP��]�$߉��Uo�l j��gW���SO8-]4�FA�}�t+�<�+zfY��U��l����J0�ڒw|oV����ɣ=+����n�R�M鞚:��s��Z��G��j�x��#��
PBk��dm_ͤO��u˰��j_R)��Z�ৃ��$~�>���ë\��o҈��TZ��';[�lU/�d��%՝��Ȫ���I��Y�E�f��S��ͱ�Bi�Ԅ[X��5ߣ+$�P�)Hl[����;]�_�{��\��g"z��X�wf��;&�4���IA��O}4;H}M�c�M(�!�6g�n�L6�xg\��.v�ƦR�|��#�����-��T��?>7�J���#&;c�j��=~�m�n�HY�6
�r��(0)�ns�)`�5װ~����� �#�m���'�	�ҵm��#�z���ey�1���z�*.�C��T
�����\�Eb�*�;���:s�P�_,F<��Z�v61�	E<f�l�d����k+��G���d�!����٨.a)����]K���n�
�P��ֱ�z��5�8n �߀��j>c�P��6C�n�:�~�����M��D��n�����F\�P�K�",�����V��blͧh]_�I�� ���e}!�W�J=������*R���=�I�B�DI�;�L1T���������;��2�I�p��Rp�Դ��ռ@�ǐy��K�W��j"�BE\g�,��6����FU���A�D'R���
���}�
�?��4YU����߉�d�/��OQ�-��%�&8�w� 1A����7���/�_�ؿ|M,��#�c_���c�BŌ�sD#.�jL�o)��D앑,��7�6��y�zUL6QҡF����p�k9o�S'��je�Pf�����G��eD١�*�#�u�f�����M"PEN�#�.	}�7���3�i}��5�ŷ�q��g��rQv��ܬm�ծ��Hx�8�Z8�g_W���m�Z׳����lMݠzB�}����kZL�b���_�~���v�������X����55$︱Ez&�r	��Y�!�#�s�7���k��	�px�I���#�(�p�c�4��n�����Q�u(0��OHC�g�4c��^?<���~��Ҏ$j��ķ�ћ�?�):����.�.�#���J���f�^d6XeO���nueHg�YM�fZ��+(`�4Z���8�{DP;�Sm�������Ӫ�0�!���妥.@��c���F*�⇇�H� ��BOFY�x]S{'O�E`.�׌Z�Z�"`N��ݙ��f"r��f"�,|��$�cUP� ���o��!��'� �5O�䋚?y��+qW��풜�FԈ��'|�=�$�f]i�7dƏQ����wo�OMdj�J�`�xk�t�#���h(G�Dl�~�ȶ�D�H�;glO@5N�AWs�o^�}��u#�=�L�b�?�&>3H-!�w������X��1�L]m��7�Nд_AԗXl���`���c�H�$۝�q ��Ǳ��Bt� N�@�ؙ�Kp$�(#���*6���9u�T��U����7���;Y ���"e�N�*;�|���Q�!�}H=�o ���Q�cf�����k���u��U���g7L >�'K����&�&��-i���}�����ѳ�w=R�6�4D\��X�_�]�䄘��E�W`��)(�9�v�3A5ʖ�[}r�G�I�s+��m����6vfŴ�d�r�gFh�j�ZF�T�XG6@�@�H��(��[��=�ʢ~�p��-}O��4o��R�_�H~ЯJ/��ݱ��Q��q��N�Ex� �b��}�h��j&T�'L^�QQ�daϧ#�i�
������a�p/%�u�?�[T�����՘�����'���:�ڀ��NR"I��:�O�R#SΏr�QJ�a�	�/��o�l�1\_%o��Hh$Qk&�zk�F���Iç4&�s��@~KBY����Rn ��7��ݒ�����Ta������Xu]��Ek��~K�]��L��E��~�j9��|�r�q�������4��w����F�)�e�쭳��\I�
7)jխ6L�3p�y�	��T�%�c�!������)������1�?��V�bJ�H����F�~+=���i:A,��4w0�'�3�������pq� }^�7T߈�,N��v8�������`sl�s�Jb�Z=��c^!�In޺���2CKzW���ʁ!#��:�tf���A�&��g�Z�#�� bCKW�Ź������+�&��W�l����]��^7?�����FF���o����s�8~ˇS!,&����bܿ�l%YLh<:�ڤ�L:e͘l�������s�хo��
��m|O�.Z�iѝ�Õ,(�"� N��z���8�m��c�(	Bu���]0DIZ����챠����ey�U*�4�%nEz��1�oQ�3���$n�����Wk�X ͙�j2(GQ����G��7S�Ls���';��<��_����f^H�>.���w��xB�߃�w�g�h��|����z�|>�I鴡 �{�4�G�߯���`��@�rL�`�lĩ9z�����d��^��í �"��z��6f6$�8o�Y������v��ߨ�n���Pr+��J?X�������]jqw���׸�;�J�#��72c�ZNoy� �"��vg�[ n���g��N}}�kHe�n�r��w��16��
��"����nK>����׍ł�S��k�֮��e�)tT&��I���T/H�s����FkdY]zJ�W�Z�Ѓ��t������!8�}����#о�����_N�R/�[l|�,v�w�߄��Jm�PI펋�zI!w�ʱ\��>�����0�����}*7�#�E|լ?<��S�)��O�j=o$�����CB�E_kƑx5�e�#5���j��]����V�k�xps�l�58(wں�eK���Ż^�bD�Yke	�,_��g߃ /�����T�&�E�
�3��LZ~��c��=擙�bڿ��H�uO��z�ʧ$��䋧8HSS���$;�5�D����j��X�q1n��K����~n{a8�;.����h{09Z3��Ⱥf]���V[�{��XM�/��đ!�WKs'i�_�]׹K�*B��?8�? ʭu5;`;?=;ޮ�M?�i�F�y=֘㋳x�Q��Ә�i�T�L�� �P�*H5��n)�B��_f.Ԗ+��ƅI9+�s29>ӗ�����n���
G|: �+?=UtX�5x���DM��ʦ$=�#��Q��,T�y<�D���zL��slU�C��>FO>(��z:ߴ��ϰo�!gqրefDX&��+i\���؛�UBf����B��T�v<�'�(��@�g���k���A��1�ޒ�e%�?E��rD-�o#�_�!�E�*�\��<Q��B{����Oi4�R�wE����hu`<�+!'���'�����-��%���+YXyF�A5a�#.�kS���A��G`vnK�j�<(�:��K�CGFq69p�XXPpb�℟C�3t!�c�#-�����{"&
�c��L�1�ԗ��m�ǘYC�t#^*�{�SL���|��7�0D�����n)i��A��CG;��aܴ�|�uz��"˰h�D�"7w�.v��tq"m��
�+����!��mWw�� \MD�7��"`�p���5�J~������r�A��_� '[Io�\h,�l;�f
����޾K�L�,E}��XX�kN��fE>��q�[�L��Iw��>:���E|^u켂�c�X�$��կ]��?i���W�A:%��t��i���P_���t�^�a��a\�{��iD(�PF���܁�`R�ٷ-���[��F�G7T~7:s
G��nK��CI��q�69��v�o=b<�Fki\���/�&|2�
 i��#AS��(M&�'�@CɴT�����x�B���@��T��j%��-�X�5a�.hN�O�P>���jzj[|c��ki���YG�F�