��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�,(ۍY�����޴2�bT�y�pAQ{A�}`*q�6�ʘ���[�s�ͼm��!מ�_�=��͸�p��Χ�Q�9��3����MŮ��S�>\ '�Z*ɼk\��.�+L��w#��T�ґ�����,��x�zKO.���uV�UwsRn3p����a����xcț#���7�C�:V_q�*�̾{�8�f؆#�hQ����O�Y��5j��yIt����{w4������T{��XmN'�L�@/i�}���]�:�S�7�U�j�o��d����t&�6KT҅~q\�K�uB@���(:SZ-:�S���{?<�!�s*�EO�NP#���V�9H������_�u�nxn7N���S������=j�m ZU{_u�]Å;�:�؋	��F�*�'7�dNTܤ�k��{�� \���ָ�'F!DW��Ƴ^@6�+< �o�ύ����&J��!���du�(��!����yJ�=#zg�;��m�������� tR�!���1좧���Ԗ��]��ȋy�=H���b��E�S��J��v��9K��)��c��� �c1�h_��$�Fp@�fQ�|i,�ux4�P/�ҷ�'24�@f���@Dn*VhW�|C��#L�W�d�L�y+%���o_|�Ԝ6`�Բ�۽nud��^2�3$��<��b�˺yEȿ�U�p� ȼ]+�#�
�?��4T�R���:��=���� g�<5ҕK�r�B�Bhp��1<4F�!nQ5��?�8C��)��JH�?�dSs��>M�.�Bo:�E��$K����d��\/��q=*Fj�\�fg�$GP6%��x$��7h��l�{����g�̇�u�gp:�����\!�I�]�&��`ۜc?� ���)��`wh�v�E'��xM�I�FƆ~�\����';��;�z�97. ��P��L�g�d1�P������s|� /��c��  H��3hQ0)r��2�k��ij6:n��(C�a4��VL�a�
ۗ[�j(㭌��c��>X��t�{?���%�������Q6�Jئ�#rv�Fb ��Z��f�`�U9�K��Vr5`�㪿�cb�C)��+Y��8_/��C_
�m&���Y��3�@M@n�#����RP����s�A��bu൨�}]~�Ga7I�L|�RV��M�z�'#����-1a�QŦw9>j�z��> ��j�5�`��w�c�Z�ؠkIY��Ӯ�N>xL�A׾ВItI��������ɚܮ��C��|���]?�&�պ��L��ͻh�3{�5�}����d����K�u	:3O݌����'�Vs���o�7*>�[�g?�8!�R����C[2���?�)�t������Ѓ�%�^ ��ٍ������.j�Y �]8/1&��R�f֊7Ti}~��{�؇�Α(>�Hg��=.W��d-c�R~�@VK7y��_��q�`|�@ٝB�ӫ������˻o-`��yr��É^F�/q5KV@n���O�[��x!06�5������AV���2.�5�)�-e'wL���cK.�6�����,?���eN�+;`+�<KN�^&];5!�F������	�ˀ�{'�~y_�2�1��G�as�mۆ��z+e����I-(�T��Ψʔ��|-hv��7E��D�����g#�o�
�&`��G���Î,��<(�Md�yk����2	� ��&��uƃLq�����z�Tp�J���w���~��{�
�M�=��v�}��E��VX4�R3��K�m��V��(eɤ��{���PX��ٺE�U�Z���so�:��%Nɓ)s/��|���-L���V)���$Ia��VG���*)k���y,S8�����B��� �#�//���=`���P'ONV��3�Ae���
�VR�&��^���7�R7)��2�17؟�-��i�gr�w���Xzܽ��:Eg6p��*ј���7g�0�aJ�x��g���D��S�m-K��
_�	�d����2&+���K��۠�w�ݷ&X����6jE<�Dn���&�un]M���x�!6�z��v�ퟹ���{���X�i��@0�MM�qp)��<� �;O`] 0.h*�ن��ѝ��L�OT����Cy���c��n?���O|^���2��, �3f�q���lx��3�%��])A�;��ǒ;�����׳Z�	���~��9�ڄ2�*�Y�A�Qnɯ�b���zw���X�HSt�XR�1�ab
���i�D� ��d�ۮ_��[�y^�c�qpN��FUa������uM�¿��h�00v�
H�J�m�y�⧐��IF�e��������N�yqF3OB �[ݕ8�<w ?��)�|5LC��i�{m�J <��6��%��Q&�
&���V�$lnКLJt	�_^���qZ����1_��O�:f��!(b.�lv���xv�܉�o�yY!ډ�K�#*Zێ��� y�-�"	F}����s��w��8G��*�GqT1��.M���q ZL��ˎq���,q���t+Z�f��&��� ��?���vL����qDM172G%�dE�z֙�1�I�O	����S6(�s�F�TM�E<%������ѧ����x���ި�=ƥa�Թ��>vcO��P_w�Q9I�S�ڗ'X��n��Y�ґ��9;��t�[���ɠb||JB�qԺ�)�ZM;�?6�_	�VC2�
?�XF��a�
���Y4�	���_c1�gK+re �JtnZWx�l��2�;�ƃ.��'\���d^o��.�R��ߒ|�0i=k�z�y�u5h�Qp!�J�ه_)��xL��]����A�_����w��g-���U�h|��1�!!h.b��PJv<E�"!T�4{٦,�q$�|���{J�1�z��ld=��Q��8V�:h���`���7`;H�_�0ɉ���	��1¾'��.Qku�0�BPAsC�湚���D��es�u���$�e<�=�&����E���h��&z���I�q<7l����]���M��+���D�21Yt�[��^t(�}cd����y�]�AF푫���Y�>Z���=�&,�V���܉���^WL�n�d5D#<���]/+l��0��ڃ�c�F����m��-�R ^}�%ƣ��͙;	��퐹9|�T1uaX	?1P���d�(��Kr�����[�<<�W�َ�@�V��ѥ�m�@a��yyr�A�s�Q����鏂rf_���P�pD�}'�A�w�X��ӂ�boOp����|�يޫ�g5�TE�Rc7�0��S�0^8���/�b�n"0K�e|*j\�R&G���;���	_��IX��)���y��*�'�y�E8C���vC�ʂ����#0�����z}���D���Ϲ�4�EEJ�(�u���ca��$O`�υ}�?x6�B#�?���h�F~�?P�V",���d^�ӌFXI:���6v�^q��?~�F��h����N��ʫ��{��G%\ ?�u٥�{M����Q����W�2���
����U�Sp�l<�J5�83�~"@OL'!������y���_d�J��z���x\�Z�]�%����đr�ZV@�iF�GO��LH&���i<w|��n�2�JR�������,w�1f
/����H����Ǐ"��d����&����f��g�L2�2�<��AD�j�/�f�����O,Ζ1q��ݯ���B�24����G��&����޽n��`2k����
�\��SE��qå8���^P#�'2����>*Ϯw���vKTН�<���?R�]�_�����v�S#f���UbA����N$��-��j)^9"%ӿ\�"H����I�ￛ�[�[
`�P�]OR�y"���P�SC�a�U���D.�'3&)/��>�BR�`B_�P����	��w;�1�(F����-\%F#�Y��m�Ձ!��R$��|�T��K�J^t���D 	���q�\:3���i!��� �XM2�0��z�&�8_��9!�&��*�. �N-�du���$R�BI�o�>I���g�Nߕ�����M�^�X5�ü��`2��4�<"�u'\�f�B���l�y\ck		�d'cf��,۸�H砌�T ��Z�gu9�9�ɾ79̯}k}9svПqx��h��aS/ %���P̐�K��
o./
j	LW����"�݈� ����Z>* W71��8�	J��MQM�L��zayM_�*��fW��������ƯKy�I�=�ګ��fG'�h��N�U�knlI�����\�x�����AXU���ไT�6�i�z�|��Z�țJG����ⓙ���tO���k����^�6��A��M���Т�k����m$���-���`�5�����֭���ō-[2tj��ϩ�5�2�:�'��J�c��d����+��U$�M�X�s��؆� 3׈
�3�")7�hR��.�1ДI{�˽����fHK��:�)��N��ݎ�+^4�^�+W=��� 1�F۫��ә���hh�	&��ۉ�x!p���O�G�)a�=�q�H�E��U$X��B�=�r����3�_�Ĳ�q�e���yyJ��6��l�L�
�i ]-�2$��tX�	y�2H�Ŵi���i�}�����_�_�x@��/	Oy�:a�����^�w�"�
	�V����ї�ۦk��0`mg�q0��C���*��LݡN@3����s�^|D�ӡ�H��3咉1>��~paI$�m��DyY���������
wo��Q���X����D� L�*LL��7Tr��"(�j�l����6��=z�딈��o�}�O���	��\���#�	ڼH�4�U3�p�VV
�?��K[]qH��xEГ[����s�_��S��M��d���#�&MS>����6��vi���p�U��e$�F�X�Y��曢�P��m�4�Ŗ���zU�g��A훝�3��V����G#��EJ�ݬ3d"d*A�$5/O:u���T��M5z;��{�����jy�E3��l5����:Z�_�&��D���{O�4�r㿦���Y	��w��	3��E,�����	e|]��|��C^q�ܱ���0E+�35	��� �_ T)(���{��;�V.��s,��S�~$�ϒ��$�5.�І�,p��FR"cù?lb[�p�Ѽ�²�T���<��Q�-�?��I�cS-�"�'r���3h�#�u{��SB٘R3LP�}���8��k�÷��� C��m�9Ҿ"2{J��	c�͑k!��w9��&���Ɲi9UvHF��J��5tg�����2���Y�2��.��EQ�g�BC��:��z�k��$#�[�j�I3�[F�n����0C愤F������"��V۴�T��X�_͜��)�l@OpMmm�s�߸�҆�cEdΤ3�#U��wD�Æd�[��(a�P&�t�3@�2��������dK/�ܷ�Y1��z.
⪟�a4�0�hcC��ʂu�1��1������-�z4��C�@���`�Q����I �m�����H�0f�GC38JD�U�h5L7g$#:fG�B$
��n�	�_�㎠Õ�I8��/�G�]������q��2�/�@�o�P�zlb�S�(���]��t�õc~ǒ|�h.�/����a��6��́+�{�F��F(X�پ�B
+�(Z�#��_i��&܁No�q��լ�ϓ��ڎ���=�&E�e������x�7FzJ�����O��k�A*E�56�8�Oq�
���X�5z8�h{Q�o�d��D��t�4��H�'�x�ӭR���{��������P�·LX�z��_E-HG.��4�w!������]aip��a�`�����{�|�~��m1���]��Mo��#��ޅwe�����z�H�o�˔ʈ(눆��j	��&��fk��1�lT��мt]���j�\���mQ��g��S���-�q��;>���jm����N�aՕ��L�۴��.�ͻPt�<����*��f��8�\� �惺�V#v�c-8(�%��
��L�PC��U�,1�K�RN K(��1�e� �꺫RB�8�7g1��G��(b��!ಀ`$Zr� F�eN�F81�U�ź�_	����J����mc(`,��A�@Tk2�(���F����^ퟆ01��8���Q��K��jC,P.��1�I�
p�j��kT�5n����)E�Ӈ�C Ra���y"����L�kn�j�?��eQc_!`�׍T�_���S%��lP���o3��9�C6���+zfV~k�[7����)\�ZW��(-ȸ��h˭1�:����8a}��ɋmYL�И����P�Z2[T�ʅx�y�)��E�(ɷˉq�n/
�ϖ}#�g݉i�ws~��>a�.f���q�V���<��C�+�Â�m������%}�Q��Nk ��`��?��q�9�Z�皋��E�4������a����]�\�m�"Q/��=R��g��GS]+��daݒ���Bm��i��i3sC��4���r=�U%�DQ�Z��w�܄�XI�,P��D�;`�@'EM,�gEX?U�X0"�T3F��8�8��t�n_�m�qя�g�.�/�p�R�N��Jw�,c��,:P#��1N\t�����WGtf{�Oj��]%i�&��,��tU��G.� �ƞp +�\~��=��*՚�ԫP��9�·)���!!ԉ�'no���>�tU�K��y״�2In�ӣ+��yˑ1
��S�cwf�e�-'o���� ���WM�}���853����Ԑ-&�.u�k�j��U�z³���Lފ��'���1�-5�SbzeЗ��b���n���A���&�����V
z�0���æ���Qeb�g{���7�"�gZ��oR7/�<��e�	Ж��������%/A�����\m���~�����}��)��e~����IRY�QW�;ms!�+�m�Q|q�;g�,@� ���?��>r(C(�B�m>h���Zc!�29����a�D8,��u�]�*d��>�E3��m�%������&3�߰�@F�8��Ѹ�2�ђ��B	x���f�a1�W`nk#>�?�Ey��e�E-]͹�'*�f��N>��dŹ-V=���ҍ��xãm4?"��-�[�
�B�n�������$(�!ʚ��="|��)ĉ}4ƈ�!�v�rl�9��{�k(�=��8��C%ə�dP1���?�t�z(���L�o���g/�ݕ���%�N���O$�0���qSz�Qf�G��|6W�%V�Tݢ ~���o��{o=�h~8��Y�P�\�XSI�?#�^jm~<� �K���0h�� ج��������l�m���Dt}3W-��Jƪ
x,�h��|So��K�7�T�=J�X��i�䙯�;�+UD�����Ă�W5�"���D��?��,�F����؊���t�����JH�`���.���l��mGt�Q��vN���U�z��!�mµ�����缴��yB`���b��x�:H�v\�.~���cJ���0�z$�W����A�g�,�f�5����~l!2T�+�00� �����������A����
��EFy*���Q�AZ�D����b��NOr�J�[�L$�i*	�M6~�J(��dl|+��@Y΂|�\g�u��T>eJcF�AX�S��6�=��so�.;�7~�T��8�SL���>Ѣv��!�p6VU�ٳ�WF=������Ҳ$���5�����8z�/)F�&� �~�ڠF���w�I?�>n����5ݶ��VX��H�<]��7�i!> �j�IUj�+H��t1g^Q���S���(����/t$�h7�^VL��>�'�~!�^�]ރ`�>߶ܰ쀄����&�7�q�?i&�mM�,������.IB���ѵc/�+�!j�	�ȑT�/j���M�u�YU>k�w�����jq�(�_?�����M;_�]�*{����3{�^u�A��#�X��h{6 ��r-�)�n�::g S2�&��}�=�L�ۖ� �.E�a?/��`c'k�F�<z ��:�YVοi�Z٤Mڦ���}au�N~�U������������˂r ���:qW�R\Z��G�0�o9S�w���I�5�{�$�;�J�]��Dvq\k�P��y��`�OkJx|��J�걼:oh�o�,���-ӛ��RR�乪5�tt�?+�=ҋ�q��$�Y�eb��-�A�k�Y*�����uW2��d2�a�����Ɇ;]��c��Ђ���R1�:�<��T&36A���
���� ��]�k~i��vd��l#Z}P_�^�V��X�9�j��tK_� ١}cN�g4�3�ϖ-�� ����jU ����lѧ��z7�������|�Ӭ�m�P]u��9j�&N���r�#�(C��Yh8N0r>��k�u��rE�|73wz:����u�Hfi\���$�j�I�����Ě}��tG�|�oр[r���b��r�q��m	�"�|���Ox��~0,^��.M�e��~�Ǣ�`2a#;Q8�:���Vi�q����V�g�]a�zW��򩳠���bȚDM2_'޳f�T^!<AY��ڶ�SW1��,�$1��,.�x#W�������N�;}ͱob�Ӡ�Y��u��)�m�2�1�g����I[���wE��l�����"ݸ��u��>U����<�J;���+��.\���F	�x�8�����S��+���ssC������L-�_��	��=�O4�8�l)�(m�YkFt�c8����5=�4_4��7σ"����{R)�*�S&�����~ ��RK*�PYΐ70qJ"��`�\��~�PN�A�!p�d��|G�ǈ���f��K����%�φS��
�4g��
@6�������0���(V�JW��i��ǽfReHf�/�J6���b���Ǫ�ࠄ����ǎ�#p���ϔa]�ikj
�<�Q�-�!�K�
�:��'�O[9`.}R��@����1��%oT�B'�쿘��>�����w���)f]�|K܎��Y�Nȸ�?����TB�mA���6���)f��c>�jp\uk��H4�hޫ����s��AT��(Z
�&�3�!f�h)}���[���MY�� R��D��mZv	Hɞ���)����V�ݷ��jWW��z��	m!.0��1���5O��(�Qw_��Je�`s�k�����5a����Q,�_܉�kΞ����UQ��B��P�Q1m���@B�w5ծsd'���Z�4HS���{�K�t�8<T�5=��n�x�<0Z6wN�0�Ձt����(��o���p���(2RX����@�#׍*o��R*�&��iO1Ly0��ƹn���c.W�`f�y��2�-�?��O��#ԁ�'����Ъ�uCx]�Zw�`:��9��u�̃������(�c���� 
l�������=Erʁ���W�����1�?�յS���OK��!��W㮍f
��#Z>�UK������m��v�$�f�*�K���W+�1QN�[�]oX�ww�����t�e��&�t���B1&
�3Ŏ���%��j�k?�Q�ȱ�.U%#�'Q��[�ٓvb�w7=���K���~_f2̙'�	ฑ��;����ݹ0�ír�� z�Й�����ݧi�d&����A��+M%�����wc�"��rxHR�JVx���ةH�w%"��<.J1o��9��Mqw���*{����=O�k@e�������`����nRꯊ�� / ��ֈ<)�Bv�`��(�@(�2O�Rd]�f�`)Z2�~�%�b16���^�j����`��gS�d6~��}Z�̈�!_#uH���t]Jo�۟Xb�BB��E̶�Ci�}��q�.�@��M���6�?���b$�_l�D�sae��H��Ξ�!1f�s]�g&�V+��ܑi�N-���p�1[M1�M�Fa�NVV	��e)������m;�f�r��Gu)'���W�W�O.n�8��UO�(��0�@��5b��y}��;�f����<�q!�c��`��?���A��m���j��&�6d���L���@��ʲ@- �+y[�`��V]eL-�nǜ�PG��2(v:C;�\�s[s��fU9qn��!��f{h�ӯI��5W&	5ao���a��"᠋e���F�	і;c�$���"N��,��G��P�Z��X��w�x%��J�d���7�C������CO[���T�Q̿MK'��PZ
$�U�u����y蒃T�B��naS���<��{��D�c<����^+��T�%�Cr�j�8��i K�Y#��D�Ο����_*�SQ~�b/lY�78����@h�|1Ad	%���ѧ�%�/G���
R� `�ΐ���\�-�#�#�#&<~�%K�cϺ���p��U��b�ǽ�����࿇�4q����ԴJ��E���hG"@5Z�r.�残��t92��2�wOyE-0��Srn1�� �,<�8M(*2��ٛ���f��&��u&Á ���:g�\a��h��̺� �qUx���32="�Ƅ�+���{|�2RLζ�S���喗�gZ�Q�$�k�~ދ͜�0��>�c�JM�ޛW����z���d�o�t��LC��	eHh$�5%U~g곃U�N'E��� @����j5p �Y��U?:!��07W��?�T�O�%��Re8��0	����%�I��\/R���g�u�)��9�(~�c˦���g>߯�����E��dd���aDc��L�&>����
(1��Y`��"0�u�Xp�J�h��7J�7ݗI��-�^%�]�)�co�����`�t��)�ЮXѰ���1f�T��!��)�m*S�*�7�����@�2ݟ)�b��D��٠���6����'X�O�Q$Ҁ�Y�W~*�kC`��s��P>L*���+�MK�И�P���Ǧ(\���CU�S��@z�!f6�����b�6�w&P���)R���4�����+��0Ұj�ېk9,S� Un�duwSp4�,4�y)B���!��1�y��~%�$]-��m&VB�Pp�/�g6���-�$R�p����vZ{�8K����p4ᑽ!���mJ@��~4�'X	��^L��A��pqVOw/�Űm�����֐x�*�];W�ۡW�8����*���K�mobhj�	��[Ӕ�-|���@�����{i?�WO���	nu���
�Ծ�,Mҏ2g��a���e�4����f�����iz+���舁]�G��N��L�F�(�z��РЃ>UY�c�G5�U��Z�ڛg[�m�x�w��.6T#�Y�b؀����Ȅ��	5�EX+��P�҃���p���k�3�\\X���_o�8�8x�Pމ�����2jh�}qZ���m ���B�Ar��u�q�L&�e�ԛm"g�3�&�f�n�����[��{hu���"��%i�H�b��C�lH��п}�gGI:��(������F�G�0Q����w7wkj�$X�nK���F����uk��k��Dd�>���w���/���nܻ��"��j �e��*�q-�Rr�[�6#�V(�0�����t?�
7��Gz�eBZ���j=?B=sv��p�2�x����F&�|ղ�,�>%�{$�o�0��L��-��֪H�+�~����BVr��F&[#����w^���+*�Ŵ�Q7#�B�a�Ή�C�ON˼�����KCj���v��?���n�{��0�^l�5ԩ ������t˒qu��� E(�}lk��>ⲫ#1N����]sA����H��B��O����s��;G_�dEg^F�p;��:ݥ�8�D���AP	�j&���|o�ޘ��'�~ʋU{�Z�J��Sl#"t�G]��@a�ƀ#�>�)WKXXcT�8>���	�n6��m �3�H�k�	p�hd���/msܑ���:a��.���Y�x7�n�ݮ��q&ZhR����D�C��to-6ȓ}�1�U+�{U�FS���5��g?ef{b��F�� >�^�ץ��`1g���dqJ�x�-\61K��eЬ-X��L���,���~���藱�fK�Y �J �8K"����T^q�Y 2��g�l]��P�� �L�\nIcH=�\s9�Y�����	Tƻ�	sy֟���MItTs�x$���L�'el�i��-��P.�E�*���kV>Eb��'�؈�w�Z��|s�T��U
&'�WB~��hz�C���GJՈ��p�-zY�!�p�|5�<k�<14�����6ɋ^�u��f����vT��y�k�+���-9��s�����p-,,G��+l���ja�9�������d�1��@�k��"&�ɹ���@�8P
w㘭�p�/��+�{�܂g��pO�W���o��C����{���@�0S1l:cR�m�Y3�ˑR�"<7�M;����΅�4T�1o%_'~�p��vBT�B�QR4$����:QN��z�)Tc�KѰ��M�r��b�M`�";^��[�Bng���������,�;q��\�r���X���O)Kx?��8��Da+^
M�U�6Q�����`�f����/��3�f�8JG:�i o�	�>C���^Y.���d �te[�J�����둖O<8 �+H�F�{/��3ȞycHm��p% ��l��?�Y�څ��Sv�/����ʕ�(,_x:�����{ha/�|�}=��:(�����h倅��ʷ��·4����c�Y%븢�zY�mo:T
��fF�C�U��Z��OkM�[��A��?���}�>g[ ,_�ݽW,�k�o�ū��#��:oL�m�oW �if��J�j���?�'_���1��f$e��8[�\c�
���X��1���GǍs�lQ��jr*ř#w�K�],�F�[/�.kW
z�	�n|����	�@Y���"��Y��ȝ��|qkC��o��Z����_��,�d����Y�JW������[�c.��Y����I��"v;�X�C#jcü���C��W��kq�_#+�;Ӥ�� ğ���$�yotC���I�ם�����3A�-.�u����tk����އp��*�r-{'����M��>@��_�iB��%K0;8�US_Ul���"���,˾O�nƬ4<|]�*�q���}�:k�5=��3s�4�oU�VT?{��R�������Rr����%�մI��F0�ߠ	;� d>$QX�Jb��z�ǏOx��?4%�ۦ�Qx[n�M#74!2��ҽ�[t�M��d�0��[U�Qb��3�n�m�o]���vmF��5b��.K�u3��u�pB��Yt��%���+��?�H�|�R�ࡋ�?���	�.�����,���C�5��� _[�l�Z����%M�[���(��<^��u��� >K����_���Ր�;�m�o\�+�Y�����Ÿ}�S?ń��A~���{��.u>��jּo.@��"��Q&��Ӓ��A�G;F�|f)�oʒA��[�Į�d\J	�;n�Mڿ����h�]YWc�=ѥ�t�sT���~�jI7��k��N2OC>�T��w�����bBu�W��{�~�?(������]�"Lڞ"���>Ap+4h�Rݥ bT�N#O.h\D���س�'������0�i&��\��以:���!�b����#�I'��|��R#��y."^��8�%�����.l��E�|[j��WZ^��@�o���M�˚T�A�J�TS��9�Y؃�U#��-7#M�qY��D�����N�6�RdF4X���f��AS�L�A���f�T��C�N �����J�N�qof��3���C��9��%�/'�pdVh���J�Z��/N���6#v�v���|���,�4,:�$q�Kb������@Q��U�9���t�\p����c_��D���Z,ӈ�9�WUR�x�#ȊF�xb1ٌшQԈ��b��[����Jw�d*����C��*�Aa��%��(^N��V�а��W�Nq���P�z�&e����,�rc�&j�G){�P)�PBo��-�my+x�D����QuV~b �#�}�SE�;U��FW֙Wv0����)6W�~�&���!%A�ᔡ�ݑ˰0����MuE�$
���5��8�m��Z��?j�LCz�*��|bf��g��[9OH{�2��+m�:���:Ub%s��d�P�@Rʹ��q��_�a�9K����<"Ϲ�U�j΂�����>4R�������E�ɯ��%j��s�AO�e��}����61ܩ�!+�@�5�̂f���P�Qh��Mq�I��R��#+��^��H�P:��7��3L ʙ����F�H�c
c�!Ԃ=�R���#P��q?�@����H��Q0��d/��M ˧W���kX2;aR����,�w�d8����0�7 ��c���"�_�F%�K�`���*U���<[Y{ �n;��yH�B��O~�Ox���셲�co(*[1Nb�=?���r�pb�d+a�n+J���pw3W��Z��;��)��L�G�G���^�����;-��Xӫ� pT
��rLZ��� �*�.���������)�!]�z����U"9�Gvz�=�[��KӢs�	���]v�����^m�,���"���>���rU|�t�M$�KS��=Lurz.�a -/DZW�1�E��Q%�ZF?�u$���u��e�x�{�����7*� Afs��^ ����d�2�H�ў!��>}=h'%�������ߠy�$L���f]Q,�Ǫ���1(ά��l��me�� �J�_@VG���#��p��0A�?|[Lh��g�L<�R��-@�w�6��iA�����^�������h�+�8��P痂�Ƿx����~�MoҘ7��-gm��4#�o�T�p�J2c��C��I��!dE4�����ս$���\����������f��A����`�)��B5G�?��b�Jk�޼���-ȼ�����8L��a��Y��ձn�rL��i��f��;�YF��G�p�L��^)��>*��ũ�W9�;u���s
h��n��a� �>v��q/�qW\�L��p�����c�g)�C��`�)��R����ʶiMz;�3��P��3�W���U��hط�s�\A�fO۫kέ�E�FX>GK��[���0b�Fe���Z6_
~�\�
�<nm@� �x�L���CVN���7^��WVA��c{j����4tm�G��͍��ų�����>�c-�/�=�\�E�j�H�f���XbF��±��䮍㔦;�&>���8�ċ~�:Ԯպs�/�&��=���7I��%)�@Ǥ��X�}1��0ҙ��o��OF�c�f��[鿶ӣJ�Ƿ�7�s��:t'��FZ��܉�"v��Q�� oÇ<"�w2��� E-���a�Lp��Vr���;y��v~ɱ����ҙ�y��Y�N]�-��ش�h�pAG��3�}��%�m�z��F͗�y�z4�???�4438�>����s�#pY&?�c�:�7Ul����o���	��Yxg��O�wB�����2^�>�F(��m��δ�j'��T���w�=1�\,^���yyv���L� �3���>�T]\���ң��U(������8���ȁB�X�2�Z�>��01���"�Yܩ�L>�9�U,�n#�?���(��d�$��!�˲/׍�3��3%�_ҙ��8�>�F * 9�h�S�*X8��1
��HR��+�.eg��i��h�Nll#�A�<p�|�6�ܜ*�_����D�zD��aUVϐ(����B�<��c![�g�ֺ�Q$;9)��o�5��Hǜ���s���h�HMǮc��I&G�+�5}�%�B.�5���K��ad`Ä�l�N#;_o���Fd�yz��m�[d1��+/�\HGJ��C?}}_���1wJ!�Z��H�䷋����U�!�%���4B�ڡ��(�,���!�o�b���Hn𓛹�q�(C���#K� ���ӿ�Fw�]�C��xC�3O4�]���p��2��MA[�}@���1�E�n�WbJ9*�ER��r���ya���Г�_��<��R��-�q���.΋�泍�m��r�ǹ9�e����a�҉��%_NmW�o��ةy2��:Q��R�*1�0�Z�n1_V��L`6	�k��O�h����&~1��a�2��T�����7ʰy���h
��`yleIa��';*A��Y��J��Yuc����L�e�9��<��I�BrN�(���g�u�DGh8�uk2�pL�~Vz����6�8���e�-tJ��n/~�Z���F�И��-���I��t6I��^�f,���}�j%n0ꔏ���~���c�~���,��<��>D������m��k	�4��_}< ����ָ����r��]/��������e��N�{��Q�9�Y�kȘtH��P��sU7+�vڳ��u���y5��!]�)H��ʥ���-��ma;���pw�Ҍ�~�����n�q���ٻ�4 �I�{C�|�u���tz� #(m����j�UsD��\l�;
��Nר&[I��W�N�'�5/V�Oρ���Mf��0�r��\�{�`� ~-�=�N����[�W����#'d��i�F��p�w,C���uA&E50�3�,#h�"�����YZ�_{�:��\�}r֛�6c������x��7���ya�Ex�M�Y7�[L��r�I�F�,�V����*���L�ޯP�0���� �0ү��w��V��2����:�U�Y�5MҹX��5^F�L�ާ�ګq�bl�/b#�փ�e�lX%.�8t��c�4���frV-��u_�X�o2qAȹU~L�?��ˍp�g���-�}�P0W���^��j�|��\	ު�-�:��
�\[��>������[�;�5��UX��:}z�5�V�1\
U��;b���`�_���]9�/��D���2��[�׋��y��p'ް���HU�]b�bh6N��c�c��-�'LD<r[�W(��\��i�'��f.ϋ��� �I²?*�I��Dm��)ٛ+�-N->I���a�즵|��j���:<G�%P�@����OR�g�Oly?��@�z��|����8S�]� <�\b�y�w�ȶ��f�Ѐ�F�4'zg�� �~�:.o��3��4��չ��~�w9�@@�|k��^�a�5~��CɄ~4�bd�z;Vy�횳O��S��<� Þ�1��� 	�Ĥ{.*���{�6�s�}z��t�������'����<��~#�u�򑢉��~�B=��Ϡ�J�O}m�q����u�����۾��=<�Q8��<j	��J���WχN�����'}%��x�]'o�E^hw�8y�D ೐��ll��-�P�"�#�P�8n8T�L���Y�tw�J�qƬ�C�h5?za��ʻ"� MN/U��.d($Y�Y���BV�m��S�s�n�^�(�!]�2�X�9:�f^i���iW�*�CY/�[�;5g���6`�>���m�%w�h�7�o'���d��%s�!t�!n�}��Xj���mX���0�������R[�8@:i����S+�������wPD8A���ptf̦3��r���%HFwx���2�����X`�R�X��`g��c�os�)�4��}��	+�z遻4 F���ZXԱ�$�S�;�>�b�V�0�o�a!�G$�ֶj5ѷ��{ȶ�ٔę@��R��/V-f����`�Gd����vV5!�\:�]�a7���̀�uw���5p�K�z )���|֥�^]�#��#�z�h�G�H�w��X�͢8J"�����:����{����&����ܭj�"�]6H�m�U� �;�k�1��g)7�l�j�X����1D�,e��Y�G6<�TT%�&��Z-����b�h�;t�fE�Q��H����V�+ƪd}��>�gq���^����C��EEY����=���<��Lf�@:��$+.[U	��f"r�t�9'Uf/����\;	E[���?a{`I��U�ۻ����^�ڼMk���"M�s�+G������b���N X{����!��a�\�G0@C/54t$�.<����������3Ø�.Q���bI�X0�A���c�`)}o�2�r?-�����]�&��k���_��S�DV�Lj�5�;/���y��
 <\L���)"N=*�Y��z
�,������{׃�?��|��&��P`)qd�᠇\�rgw���D�Y[���y�E�+��B�HJ('>����f��bKRU�mϣ��}��{�b�g{��u�&�/��c���%8�P���4J��Ŵ�.r�_��N�hjfH:G�/7�Y��T�~s1�I!h)5�R�%~ac�����3j�N�(*��ʙ�ڑ�_!k$�"�<l���A��7�C�.lq��(�A�����{x>a$VD��GR���̩�� �C���/���O��e��#1�v�vp�mXKu�e�b�]�ΑF)�_�"8�`$�c��c�f+[�gG�Ǔ�mC�zw���V}�[����1E��q��?�6}����5�G����Hޏ�_=��Y�����A^�{�M&4p�A��B��x[������ }��i�i�q���?I�i�c���>:S��F�=0�v	D�V�������n-uc,����E��>��wW��Ns=^�!w]T���{�H�)[-m���KQ����Qi�%�Ǝ��I����C��>\T���^6� ��_BS�������ؔ�[dTR��^�x��8������<o��F��+�u_t�g����Y���F���yfݰXOf�����j��4&Wɮc� ��������vr��q� ܭ`�e��_�$0zX<�e|ە�(Fާ"�@���\c��ЧBə� ���)�c;*>�	R>p:�����8��=��Ƀ�X�R?�xDj_K^T��dÇ
u���-]��O�e��b��3A��A��e%;�3By�\�hL�&g����3�~ˣ�ʺx�!r����Z��q�^�$��:���^(��l1·ل#ܰ3��	iT�N�z������p�pE)1h���`eC�s����&~�����!NZ�-|AS��������I8����u�$|.6f�Z����|��;o���g<�^�`��`7���:��_^��X����VZ�A�w�&�o���!;k�9f׀'��C�d��ف��$�����h���YK8"��)���R����W��H��6�D�AF����"xq��ͭA!�k��T�;M�r6�?�V��ct���$`�2/={UH����u�˖��[pN�ӜL�m靏_��B0{�~M�eǩ��
��i�A+�?�������N�%��Z*��^?�	�!P��c�c����`�r��q/jw������$ܚu>z=�̙�/��3�{)-�~���kB�I(���ߗ��e4܎�XB��Z��xN�!��z~WFiU��L
ԗV��
�aZ�fԙ��S�Ԃav;~��E�a��
J4��FY`g�b}�b'��#��w�7��%��Z��s��*�1�li�	�5���t�Մ�|JB
@�����uP/��2{��e�O��_��]�^"8j�G��>(�����������(�\���렎3�ͮ�X?���1j����c��x��=�$Z�o���l�ԴudX��&�X���>���d��=���lF��;� Y�},���!����9.
�bz�=;��{X��Q ã$R�v��ˀ���;�t�s�[HbE�U�޴�!���׏x�dYLt���K#��S\E	�2��+���w ��@�^�'����(1�7ڟĭQuV09D���4r� ��cw��p�C��D�(�m� �@�@�6�����zwG�UB�~�i�������'����&����3�a��:#	�Qn!�L��!��`z��DN;+;��c���AЫ��-R�o�B��!���,�X�����A�P�˂��I��J�|�('%���"
t3?�����F.J�" =��J3t�X67s�}�;�~��
��e���F]=�����g���O�$U��3��y�g�r�Q�O�@^��S`N$���9OUz��͗���1/&�9���4ُh�_�Blp������
!�D������΀6�~�9��f�k���q@���܀u[���Ǿ_�LQ�S��2�����f=��E�L�P��lsh�M��,�ǜ"�j����Pj��fV�]w8wkH�y��Y;@��6��"[���vb,uྷZ�?�=�[!`D����Aa�|�%(�t��0~.��w-6π��C�ja�
��݉i���k ��_
~��a$���õ; Nt�Q�3߲��QeA)E�^�Վ,n"IB����J�M�>��!aTK%$�WRR�]ȥ햦��Ҷ�4����,Y��I�D`Xǿu&�q�]���#}z
Y���葸�O�4ݦ�9�"�&��0��g�Ar�ѿ'�|@JB�	�Ӟ{?��r+�d���f�D�Z�PǱƾ���^㝨�~�'��~_D����PĨ�!-h�l��I1������o~���mfI<�%��C�Mh�:S�\�Uj�s2��8�Tp���">�i �Gŗ��|�9U�0@U���x�q�(Wom�v��*�Zf��UDp�LO��~���5���)��3�jn�a�y�f��_"ѩe��pxm;�E�PQ�T�"଺4��ҩ�e(�B����t\�)�aW�|=`� ����{�����B�w�5]FuфCx�gH;�:&�}Z�,gR�ccn�ᄉ��J1�#���Ƥ(��r�	��)�V2�mEo̒ d�u�Ȳ�eﾨ��	ڢ�	�Ťt�&5��b�NX�o�@��ʯ=%�C�tsL�f3�9�y���dr�����/�_L��;�% :6h�ʯ,�>0$�'߳2A���ssOC�Q�4~�dҽvJy�s��j���K�������jlL�ȁ��_�f<��#u��6�>�Ρ�T�8;�1Nj�I׍�����k��=�MC��VQ�=��x�b����E�"Zm(��寞Z�U�Y^<Z�C��K�'�sN�/<9vj�w�!G3L��24!�z=0*�
��r	|�jIWq�����	�2����i�#�-��>����֤d2~V��V�TRY�
�*2������(Ȝ���m�5R��]�7%�$��w�4�U�0ƖpƤ�8$���h��Ք)�d���/�]��뱗����gX	�z��S�E�r"P����k9St/��>@�6�A�Y��ڹ��1�%G���qZT��X���N�ݸb�(�RR	���X �%�+�J\cZN�v�"�Z�^%.Ѯ�+�!��O�WM���Ar�R:*�P��`j��Ȕ,��hEF�@#
�G���p~�9+Fy�azEG��/Ю�w�g;�Al�&��yy|A��Z/ͺ�8��c�!@5Y��z-F����\�c��dv�Ou���=�ƃ�xE�g��r���ᒉ��0 ��Dɽ�:���İĐ����{��*G0Gq�?�4�;ev\�4�}��%G��y´�oz'��P{i~��pp���`�5�$>�Be���<k���
��&��XTj��f��g0�o%��&5��0,�[_1�o�g4.�h�z��uz~�dkD� 6P���S��ĮQ��d��kb�n�ZP/ݏ�$��vGU�:�|�g�u�E�4o����8=3����_���� *�0����=�"n�Nr7Å�ؒ�8����m�{R���wא����]K	���B����A�~y��/���4�qkΞx2nN�fH�]k�0��vn�c����q��2A��6	?J^^D�*{B,��K��T���g:;6�L�qam�x5�H�
�G��tN��;�nmǕ��Rmd��b[z�-
09�������$��0�oݍR�C���GY[`�Av��D &cw�P�5�l0!j%����q�� ��J�^���|��Rd%`�X
����ń��TV�K���������O��rA�m#uk&d��x_���[�J�[@��/Ux��OY뗪C(���[�F�7�>ԡ��`4�1���,���m;��n&'�5�,�U�j��i�x��y��xT���ʛبu���E�+�ΌrLayp�����'U`j�a
��b�v�ƭ�:���ĂWQ���)Ա^�Fm�L�݆O$�=�~Rܴ�|��*�l7�2q�GDgJ��`zcNf?��%�MU4p����`�K��o��R����.�9�Aix�t[NW�ϟ�&��vF.J�g��
a��xm;�+��x��pϼ�a'qsI'�E*Z��F�zs�Gn�*��=t~�,�|���y�D���T����u��Mxgs�s��5�-����ᘬ`5�,�1�P 1������1�?���LW�LB�P�JWM�Rշ��`X��\�Y��!!�������G��&ن��,�؎Yրy�e�I��	:�G���a��E-��0�<&eF�����2F#~$9?�ʤ����8�c�Z��Ρ��8�E�d��-��������6���^Yܷ�]�~ �,�a�a��b�\��y�x��?"��u�a�|\��A2T##"E�u�z�$��?x�]B�+��LB�ʒM�j]��y�t�)���j�03;���q�l�6d勤��{�ٷ0Z�[���)^��R�FeG��������,�^"�e=�q�9����OfJf�Y�.rn���9"ǝQ7^B�zC#S�sE֬*�"�	%����J��U�aZ՗d��&ؔ7���}~(����F�J��uq� �*��R�u�Y�	:.����;E�0�r�xz$�B������(Uy��2��F�((��u��� 6��꽔���C���`9����[�N3�g+�s���-�&X�q���T;��l��u^!2tz%��pl�(�[fb�e�s��_�a�|�E�&�+�a��jۘ�0n�Jܭ�;����)pt��(]U�@�H�T�x������Z.�LDU�NVc�+ıTa!�\����a�X$�]C4�ls��׷U�~]�Ƃ�[e� 3W<�7�`���hk���'Ze1�ⳣܱ&�t�Dq~?�F3�;"Ii�|�R$�խ��y��%������W�� �H���Y�GPI����X��l���Xe���v�ş���m˳�a�Y$��)�@p�h������(�(ٓ��l�A���Et'��L�{�!%�R4�ͱ�[�tc|�%/�Ș��B��q����[H0��{gE��umr�ЭF���"6��P��d.���wCM���
U��7�@����f�����\a9��o�w5��T�p	�dHg �)i��7�n��pY��O"�:�[�[G�u��L��+�Ö�S�4!ѥ�L%���H_�D2S��6���J<�-�D���POBZwwѢ����� �M����F�4=)��|7*�C;��=������3m *`�t�?"�Jj^�,�Ӄ�{#��N(g�᧣�tʞWX')O$݆�U�D�H�]�m!>��,��?���ݲj�-��j[�h���n%�J:�@{*�T:s�K�	��m�s����@
j�c���� :�2B��#J�(���X4S]���)�M1�Z�S���oo����h{�b�s�zx�:K���UP���9�[@�^8��9�6Dd8h�|@��F�MkXE��6b;�����i�OI�ge�B�%�!����3B���� pc����×n�տC�?�$�${_p'�Y���0���=�k��n����[�L+�-V+�����GRɬe<<�5�'�ިx�����I����I?�1��(�k����)�pU򡰤ؘ*#s9�SU2�v��ڎ��c}$�ѽrQ���M_hX����m�HZ9i�$;�!���eU�1�в��#g`����z� \F:���3��:�(<�+���Q�)�+�ni�%G �3OR��N��	�8$|ck�VU��`�uH�{uv�橅�
�3�#r"�Y	�a�Q�I>��pOe�\<�~�#�`D��a�mN~�0�S�˗��F��{�*5pU�P����Ms�������}����	UJ#_�}��;BK���T���Q��	#:�V	ax��#\�"%�C?[cv��N7��h���f<9k%�r ��up�+�B�n 26���4�w�&�>l|�	�E��&dɡ)C����cf)p���@-���Q�첇��^�<�B��m�R`ړ����e��d,Ku���{��᪣#Y}:�LN�����[������,�q{�"6<	�����v3R�4{N!���Jً#7uOd)�n���X}w�+ϽU_���m���w:Qg'h��b���^\@�Y�QS����y6p�_ľ�)�O)�^l����#O�w�GD�i����ܘ|��g�h��������� b֛���A��Ġ��돟º.�D��A�U+/��+?��kN�H$y�D�5�y�s:?+��PY�j��	�M,w����*�$b���[@�%��-�n��:��KZ���Q`#,���T���\�v���Z+=���Bj�7e��$UhA$��6��.�&�Υ[%X+����{���y���4�/s�=��uP-��W ߱'$w��܃����(k3c�UW?����6���������2��]���ò֍��&�dٍHd '�^�_��!n�����B[��K�亄��8��^+���L�~R!��,Jc�p⃯&��?�Q��x�?�\@jN,�]Y���O_Ci#ϕ/���e��m��{BD�Q�E���XB� �dYw<~��6x�C�c❹��T��˹��Y�#H���A�ғ�?U�dV�#k���������މ��	g���sȒ黤��/x�ۙ�T��-*�U2��)�ٓ�@�?�0{�l����~� �aZ}�UhT�"a[����>ާ�%���i�8�_^�Ν��-��Z||;�N��d�O�4��r~�T��㩼-l�%̗�����%�]�F[����ҩ��k�.&&PĿO���{O^va��:�ڂ)z��"GH6>�NX���%��Qq�X|��r��3��t���!�3���<)��-%��%^ v,OOV�xU��>#�&Co�/�ߵ�O3�=g%�	���x����KH5�����I`�'%J���1S/�pa��u ���0�8	�埄��~��'�^�tm_w��I����P�;_��F'��4&��.	)#�%�:ar8�����rg����Cab���+|����b��Ba��@Ik�b�����L��>EyS��IӒ��A�E�Y���)�qю\~�ݹ(����(v�����E�Ӹ�W��b��8�/�?`��H��X��m��z)�e�-P��I��s[�`��K]M���\��.����EI�r��,�E�+^�l����1��(_(����+4��볬[�0�Ί��kyʚ[Т������M�Vs��*���(�.8�L���L�]r}���~�w�)�͓�4�%����O�9�$��hYt0`��a,L�v�eGȷ� 6�J����$荠l�_PֺnYkh�]u�� HÉ�%J�j1(^���pdh�'`u���8�S�CO��HA�Y8�-8��_w����\ ��6᎐'(�C��1�& zA��� ��R$V���X��7@�<�W`���[
`�β6sW̙�o��D��`v?"eJ��p:����0�ʠ����z�Ǘ �n;p�&����y2Y7�A[��>*$Lx��4m3'm�=n_���ex�Y�+N�Z��s������r��#rQ���c[�4�!&ڳ��u��ւ�)��M_N�E���(��"����ܚ��"��S4����}�\�'���{��{ �򣒍�������"b�Qkp�Ǭ�c��p/v���[�̏�0���
�� WD���^-�SR��Zj���i����v���,s0����t�)��ý߳-��;ߴ�ĸ��O���x�7a���|�u�d�,�H��l���E,�0�F!�@&(2H��w	��X�=5 #��`舕�V�������b�?B�ĕԒ�Ǚn�D�>e�5VU=�h�����<l���J5UƏ�F?Â( r��������-��9��X����p}����H�ja���O�
�?z�z��!;��tP����tL7;��5�:����J����|�M�v�p0aW[I+��۲��f���I2�� ��B9 ��{R'���@`�]KJs"댨Q��utrg�2셜q7��uz����0ҊJ?�x��1�����K"ś ��Z��+<�%�qa�5i?-�N���r���d2-E��T��K���ޭt'�����;_����i��F��d6�%y���L�	�Y�)o���]S�k���b�Y�%T��W���[z�
W���N;���W������$4��+��C����A;/�~m�ڌ�����牵F�l���m� s�O�B��j���T���7����`����Ts
�u��AȘ�R�B�5y�>Z�(4�,��`N�amd��l�jb�P1�.��>��T���r�A/�����X܎�Y	�=�-�r@R.a��v[A�ӡP�����,Q��S���K�R[�6c���&Z�Q���(�����SǑ[ۮY|���`P%n��8#O�bj�C�u�$��5l��fk����`�&�������&cTi�͹��˭�ʠ}�yYs��(�{���e��}8]�To��P���a���>x%��s�e�֮��BR#�����bn�S��1�%hЮ�@�69���y�S(��Aʹ��Mm���̾���d���W3��/$2A�ly���)�q
�P���e���P���ϩ*�HD[�-��E�4"0�	Y-��Q��;w�z�nJ����d�K=d1�z0���b�ٳ;O�2uY5y��uW�M��b�{!������\���L�M���^��$��]�|�&.z�H܇Ԣ3AtA]GJ�s�!'J����2K��/�QI�JCf��]���+N/ˍ��2�i�t���"����`f������ն�����x,���f ~-=�ʮ;Vh���6"�����x�o��q��Nګ�����R��㉼�A���ώ�挕Q:����e���HM��1�L�I0� �
`���fR���7��^W�?�YJ�:�S*F&�M��t�j=�v�L>���;s�R$ ���\҈�FW��$Qg��&���&�c��+�bN�- �v�n_c��Y�R#���0�3��]rXi\�MV�;%c�n�X��
�a��i�N�cus/�G5/$�(��aMn��X��^��ReU�ķ<vN�({
� D�ϖ��U�/�P8�u��7�]���=PT��3?k'��l�րGk�CmqƬY{�d��n��W�F��qq��&!M09C1�9����(����|K�st1z�o9���t~N8�'���&�j1�������TM�in|vdO���\��H*�q���B0^����z1�=��u���k<��X��\!/�W��e�;�Ga~�}Aĕ�O^�7y�072�3/��t���Ǯh�c=���{�
)�t:,��GG��FI��	,������ CL�F���m`�c�j�ǚ9���IK��p]��
k��uD�vhA���@ߟ����擪55��[l5;bA��y�|A�˃�@��WJ��V*E��8�=�F``�N]�g��]��D�_�4�$�mƻaՏ�q���)~���f�"�`5])S��H�1ת�5��Gt[q�fܩ����]�T����Q?m�FT�I��&e�At��؛�^��޶�$�*KM��%�t_���$��pj�Ǻ�Lai��'��m����˯�io�A�4�~�w�>MoV�&�6c �"4U��mީ@GR��P@�g�����@�%'��[�Wa��cX7���� }2|�){�=s�/���1��+Naќ�� p��
f���X����Q��=�����K��=�!�Q��5� ��Y�C�tDahqwj܍B��Sav�1L�^�|J͇�����f�N�����05���t)l���/���%?վ��k0e����E��{!����׾���-¼����.*��9Qu�h=���׭�9�����e��-����B��+���ȍ�)?���м�%��덓$�[�:��u�=x�-�d��8�j�&�fY�L�� �I���uۣ���S���M]�"-�����:��`�{~V������@Z�b�|��o����E�ͅ���;��1!.x9Jj��R>� �mxp�B'�^��̮�#r��1忤��LP�\�%��?{٭����"�
 {��� ��B�Ϲ`���}�ǔ'�0Ԙܶi�-C���6�M���:˵6
ga ��[��	%9%NEY[�Z��S�|7L	�����I�.��5����҇}F��b@W�
1�ۖ
!����6?�E�(�	�O�8D�5&�ƕ	�\"&TH�"5B���h7Q1KN���q��hn��c�\��(��?��/�St��=����Lp h�����+��M��]�ezjv��k�zD��'�UeK�ް��Ո��4S���r~�p�{>�٘j���vF!����<Mf�D�r�'r' ��pU��n1���)Z�q������Z�nru���[�{@pi�L�2���K.�;���P%ur*˛�ޛO�iz,��Y�q�ҩ�k�S��扑���S�&������=9��qf��d�WW>Q�h����~/���§WBp�������ϰ��D�M����/|��P�����ƹ&R���4b�`g7B��+8�A9�����܅4:G�8@�=A�CX�c�v���r[�mc�����~g�%+4"M�aك0k��:�\�	�*�+I�fO��/$�!+B�_,�V��aNnm2�%qؙE+H�s<]�U
�Jq^Ѡg^�786�6���-��m�+�>,ف��|�O��	��*��%���C�Y��x:Th�r��� �e���o�02JV��,�j���Q���]Y4Y��p��-|p���s��l_�k���/dV匑�3DT6��-I����r�C��9��ݗΈi�X��x_�CX�a�6&�D"khO�<���de!��|ccX�uO�d��Z눚 �Q�֫�P�|��27C��!l��sa��!0:�eb=[<=ڡ���(�%s
�ªѽ �� ��۹KA��3����D�@�hr�a�Y�lf�'K#fH��w��j�*J�ySP;z��S��"�_� �pM�����5o���}����y�'M ���'�N_�3+y���i��!W�X��Q��(�Ψ#2ՒY���3��1�쮛�2��=�55�\|С��/��oҟ�
��,_x�w46][i�%�Rդ�;A܆�k�*x�l~�6�����j{p0��2RѮY2�,����	��Ӂ L�e�3��ne��T*�T��o��%�Am��:��j����=�
j����*ng�8}��ߩG
#��<�5�5!��Ά�W��z�d{��kdt"7��"���F�ME�ٲL}�h�I2�rLz��.������k�e7�"�r�_1�-F�8�z�32SĶ�6�DKT��u��X��&�q�� ����V�������/���M|:'3
B+�O�݄s�pm	��C���8���s#*d*cF�x���[��G�<F�š.˶c!�PQ�yy�L(�Tn%��3�D�\���KR�b��;w����~�eGzX��
Ӫ	�������L��\_�%�ִ���*ĕ�GY
��xd�V]��G�3�Z�E��0ݺ|+Y����8����&�[�����v��j H*���~ /f� ��}Y��@��ۋ�b�tnH�&ج��e���QQ��x�3u\�bZ'����t��,zy�퐔��
�A��^���C���5�zC�5O�\u��Q���Pm��`�fK��&T𷫁�3�^�B������h��63^ּ�k�Z�����P���A1�NE;��S�c�����ʣeM����l��!��U41@�t3���ɇ�*7>i.�	<��/�}��\{�
�G���r�۫E`5l%�&zHg�H��=̟��7�r�¹n��Z�â~�7g[�=��^��Θ�q�;��p��� 5)�a*��(�sSpn�͗�ל�'�v~�����0&=#ƿ޺<�X�_���gB8:\�~��J�~�8�7R�A���R����C/*�v��n�n����G�죷�U�2+�##���U��jz�������N�Q�����0䭡-�׹�p��C�)e �'�k�+ş�(R$v0��]��=Jn0�H!�hB�T��<�}6���y�9�@C�ԑ�s3aV��~��+)��U�+T�BX��L���i5��^A��%l��o�U�	��Fgx�!E�M���IN�N���M�vŕO��jA1��PAZ�;��j��C����K+;椠z�WB9�2v��_�Bk����_\s�	�+:N�i��P�q��"Cn�wq�]L����dm�y�Uƌ���U��+^}��Gl��;�PDA����z�FhL�Rx��fK
>�x_c��rGg�Q���:#t��S_��@�vݤtO(�t��&-���DN�kS��.�Mč�̟0v�#�S��;��iϥ��.���&AOb�FM�Z��v��-�XεP�]��"U���Wk�-�`�(�h�i��[<�[e�"y�Q���/�	����d�t�zt�E��� ��X'�i��]��#���G�[�ۚo�^��L<q��md���5\���������2�Ԏ�r0ɮ�B:�^�3@��)(��2�C�e@}6-����P�B�/���þ��˖�aq2�*��Ry�cfk�e�=����Նf]A\����:����ep�Qp��6[�F���`���<�-X��F�O��m¼//z�L�&�6���d�U��s^���Pn�oV�p�Y��G����W/
�]��a:�����Hs_���|�a������f�yV�������.=��8�Ԁ�9�l���e����U�G���MFy"�!ĩw�D]g��l	�_ֽ��n �+^�{�2��T�C��"���@�`����n�,�%�2 �������3Ƥ��j��!bA���:ji:0�47���4� 9�����/��A�G��eD͂'qHa�;A�r� Pzy�o��r}&�!��{x��c�s��]Xİ-��#њ-�ư"M;���-��������s�И�ȳ1}<d�W�ʒ��W�W��L#��"o$�t��Zu��c����Fh��!O���:8Gg5]+]�E�w%��}j���N�:�%ZH���s��W�V���P1 Ct�� f����f���:�F��H��V�V�F��]$�[&>_'t�4����.3q&�(�(��c���c}����?zN����W����`G�>�HU����
��[3zޮ��H��-���nmx3�MH�9�s���dQҩ���?���9��)^�������d��Lu$�����д��l�5��@���������p��ci��i��0�T=^^�7x�)˰�T�>{>aSZ]��֙&[�ȱv��7��8��\���f�2_X@0�@�2v�Ճ�T� �9o?��Hh��s��#=�wƪ�q�^m��A�)��m����@`? ��+�?�Y�+�צ8b06/:;Z��!|�t�_�8���
�k��ˢ�� �T�ս�mtT��T��P�e�.�Ƣv���
�@��3g�Jo�{��$P�B|9C��(�(�|�u!W�,Ozy(f^���e��0'����߬�|C�� ���z���U,:���b��;ՠ���=����\����a���SoA��7q�u9m{����b�9j�»��ڲ_MQ�z~�L�oX �A�r3Țԋ���"��`[���Q�F�E��
�V߿����k6��4(�2]�P/�����g�,��L~�W�~��ђ>?���ʆ�P��K���# 8 ����d#��SS5F��!2#Zצ�%A��`<�%�h��@�g:��ӁlTW��AP�l�b�h��2v�����0��䆾M����?���dޞ�Q��N/�V3v%B�~�Dp8i�&�r�S�ul.����wڀ�O�0(�	�A>h�@w�W7��JkW��{(p�̦��=�/��z�C�a�H��6f�i����V�"*	f�i��(������+�	&>�t������~��&�~0�d�I&��[B����z���l�J[�+d@��@2{S[<x͍CO���ʇ�<_v���Ϛ�-�x8�b�G�� H�gt�- �m}5*��0A�9T���w�n(�K��2?/�q��ڟSEk4�"x8Ǧ�Y|��*�o�͸虥��nl�tS^}�:�,a'D������M�5RKސ����k\�C�U$*c�|A����dU�W?ᎍ�L)FUhRKc��~˧ ��� &tԯ��.���l����K�`��@�@B���$ �u%�ཷ憿�����v�(9�δߨ����耶;Z���_�j��$���gu�
��L 6t�_>��&�$,�an3b]���b��Y/�j?�2�:���>垯���4�oj�$�:	�������t��j����-�|��;_OQ��k����={��fVOW4#�a��m�$e��n�
���!�`�k�x��z$�U1�b��a�3d�����+�M�`]8��g+�ˋPO�,v�,�!#w�j��^����%��!�x8$�x�D�������t.��:�O5j��[�F�=0��Z�瘦Q��uco����0�߸�1�/����IRȋO�^�9dv@{�"��c�\�g��a��Ϗ���(6��.tp�ܰ'nKI�����5��~코�y>�/W�eA�Y��6*��i4AUi�p�u���yl4�x����u����@��a�&M���R{7���4�T�u���.��j�2��ŕ?ߙ�.c��x���(�#k��튪(�P����t�F��R0�zRa�1���E�61��5���ÚX$
��[���'���@�f�?dt��Eu�y�F�`�'���Ё��tei!1�Ǔê=>��V�wT�I�����yra^M�F�[4��3��Q�kEᇅ�8�(�m��@�,�@,ِ�������@���� �)����)*qj�@���ع5孫�R�{���Q�p.�\I�:⾽+�����/_�Ճ[�9�)HX�483��B������SF�Ƒ���O����nä�-�\tM��)����"	��ֆf�U�rY�&姁��0�Zo�zJ!G`�W6����jNs(��8f�2P�d-��ݙ	j�l\G�iT��a^�=3�����ӮbR���Q�f �����O��$���p�j{ }��~��j���1g"J@-��{z]%��ǔ�AM�LB]�v��o'�.1����o�N6�a(E?�V�@˜�%�� e�
u�fr�"t$]���##�G{�����!ϧ�Y�n
��1��>����K_<Ɓ�z5^6���c����˯*���'A]Y�Q�e�ʟا��C>L�D4�O\��[��[O��kD翣��& 9)��������w�P?��_r��x���2�����y��Z���Y��q���|)��85)�DpmV����;}���c����"X����@S)^�LS�o��:Q�rЋi�����݇OX�,��(5�Q2�pD����̡��Gb����2�d"��}�b߬_�+'����t6�q�d}�)�RI��IW��br6}3E�:@���_�K7H�3 �i:��$��4Y�SWL�l�jX(�]A��p���|������[��}�Uf�"u*��fݚ��0���>KU
���]yx�L������ 8��H��隖"F�pf៘�U�:P_�	��">�3�O@Ǩ �N�@���#��.�f�Lw~�X�^�.��-,�	�ѻ%������C� ���[����_8�ά�+D;����e��+�4��t�y3�ց;N������Q�q�)��1fkk��?��@���|�b�;�ˢ�����~B�,�a��͆�s���LO
�݄�1���k�`>�R�A+�H3N��ڙ�Z n��&�;���="�Ҷ�X��;�N��ݮ��-U)k�}� r��.=�8����m�zu(�>|�6B` '���|�c�j�u��do�V*NJ/��<�:�aW�k�6�(�cp�Ì��m,�YF�� KGw�`��Vg1qH$n�;E� ᮎ�R���� I�R�w�,�����=���6�O`�y�<#*є�/������`���6�Z�̰�x9t���=?�ru���tbvE��Aq�4��A��ё��1�u33���8�1�CF�'�Z+�����&*(!$5���`����R7pN/H�"c��}v�� 0Z�|B(P0�NMh��\�^>��[R�Xx�بGU��@��	�,�ߤ���}�����>��?�b_�uK�p�)�.!LU�,�������z���W��Y<>u���M�u�Uߞ�v���n'��L%���r�W-���[�7�\uw#�3���^����"�ٚ���q풴x�c4����x���S\�� �Sr[�܈ 8�/Jf���?h{��X����x�=AŌp�۲�/��r�;'��b�j�p>����#�zJ�K{����]�!:kq�������(�K�2�$��K��A� �(��I�ks4���I=��O�q�Dv^�)�sf˼4 G�Q������< �HwQa�G���6������J��k߿ �.��
`�X��%����- ����y^�Lpe�f�$�3b������<�Vkؾ��o68�&'�KU�j���{�����w��|�p�����M���1���}d8WNٌ�Yx����"m	�5dT	EÞG�;��ʸc��n���e���] *�������`Q��n&���!���prq�B����"���+���;�Y+�*�!����j	��.�T�W�3ہ� Zs	!�`�k3;f|3��D��L1+z�5gR�=�6�!�M M7>5�q��Q�Z��Z"�x�[�3x̄Ժ�N}�UK ԿT�8olf�+�m�R��%�����<K�nO�,�1t��q>�������8v��J�������m�Lt�g~lZ{'kuª�k!�>;.����u�O�C���2,b.�s����P�������W��V��:����¬6�;h`��$�qg�-ŤB'����!���?W�$�R�׫ %
��W���w%��O�����(@ �@�����D��S&\�bš��l8��a0� 16;h�Ne�l��<�my-���)�ʝ��e���YJ����Oܸ��V*���h�It�hC�CO�s���-�/�Q�Rv��5}����H���e��O��3�Y:	�	Bh��^s��FD��0R:d
����,��p��,����`x1��5}#fJ,���2\u,��Iۊ�͊d�T-�����v7�t&���ټ��&F������If���	ʝ���Y�}����>s~�.�޺q�{���s���1=Y	��;��|�33�ުY]#f��Y)����N׮���������Es]��:�ć��� npQ�s��Em���^@A۴�R$W��5e͌�|�=f糌$y�*_���^���hFa��q��'Jf�C�C	��sFX+��)������t4�m~�MGs�l#]�~�,��G���$���pI�X�_�J�j�k[�7��ؐ}�� �{�fI�y6i#��"�b@�F���=��I\�g+�HP)��1!��"�<Υt�q��a0Ũ�ߦ.�E�Z�#�痣���,2���)b� �\��ĭ�˅$R��E�D+�s���L�ڦ�JWp��+�:�;�Ĥ+|!c�@F����G��,AQ�,���Ñ�H�W��7!w��h�G�}!�n��p��nL�L%������5�(dZ2罠��4|����TI�!�{��KGѬ�ki��C��p�.>,�zK\�L�`�J�Y�5���jv�Sט�L��@�FH%��,C�Gc?���k�/����Y1C/��u9�?����Ձ{�t՞�ӄh�4(z4���쬶�ѵ× ���*dտ�;��7.���R�|b �/8c��W4/e�Rؖ#��˳e����`�� �!] Jb�M�w�J� �kҦ�}w�1�+��O�vȇa�e���74�仄��Iڃ���.�)!�r���ꈑa�P(�y)y����tI�.K��m�*%���w��0~�p_��l\�3_*��3�憠��||��d���9qǭy�����|TDR�C�˪���iE �~=����W��U7{�$�q}��@���=2���{�,LR.GK��<O��W��k\��ϔϞu_t_�6e�����ϟ�/|v�S��o]���+�z-���U����ȧ�SM�H$n�كEݝ��Bq>UOe�%�H��C����4�}����z6�:03	=>�D��A��!.��,�\2q|6�����������}�[�X@U%���*�z�<�5ow�3#�t�<`�K��Gߤ�;�{*����x +���`L�H�PfN8؊(M3��5�X��qFAsW�D/��`���}<��pDW��:RdO��v�1S��FSs��F�n3�w/��v54
��jɐW�I�8{9�r��3GQ�(s�e�� C����<���&M!�o�����v�#q��Z&�zroMk�Q|�M�luDe����ڼO(n�;�D^4G���G�fŚ������akr��z&6�ƅh�蹔�5�uz0�)x�.��^Gbw�S`�kʊ���%TI�Q/7�{X�|�+�^�^���Q@Z�|�ᏙY�
��w�^�����[�o��ۆA�=˴��fF��"/����:�IVJ)S�®zhe��0��D>���߬ɹ��9�2��@,Ȋ-��x�yi����K5�K���%RO���%�Jdt�;�jh�RJ��X�k騞��j
X"Ee�[d@�ԥ�i�эZRH/�`�]�!��"3K�
�-�f���/�׭q~k�U�$@�q�֨c$��N�$o�`��Bһ���'b�)𳯡@z�{��"{��e%∞"�0�c�,�Q