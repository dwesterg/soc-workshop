��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N�]뭀a=@��ޚ��#��铉lyAk�М�j�ܑ���gToj������W�P*[�I`rۻbҨ�
���VN�#�R�h�II��4ҽ��B��-���E�,!G���9b[r��j���̐��~��#���"��I�X�H���o�Uwh�l��H$���p�U�_\g�x(����T��u�p�y��n��
$�2��J��A,nھ3��Ok�PO���CXGS吝3s�8Y{i��N�������B�m.�M,�\I����i�ͭ��X"Q�[�e�`pj�tq�Y�๠�5?+̼ZN�S%Y��j�%rũ^ľ�:G�hJbm�^�	��V�`��/q��3g.��#�Jn���O=�u50��GP�&��i���,�>�Wa���e�>�d����3�Q��1�QR���CWLS
�D����l��Y���I*7kma\����.`��%t$t��w$��H��ڽf���c��v`
C{|��}�B����n� �7����v�SN��V
��u�8�~O�@-��KBB
Y6:���l��~~��0�ۢ͠�1�,/9�k�q}ﻦ�%e+T~[��em/� /��\/K�G� 5~�H��&i��Y>م�ϗ�h�@YVώ�=���p���`|�6Qp�2��l_W��(���{�%;w�;eoJ9^� �U����ܗ��Q$��~�M�4��n���`+��8T}�Ѣ��ք��4�����@?��x��{�<d8!�mDg�$	�g�����d�aPj<{��B������X��οkZ�!���9FSWG�R}R���ǿF���ܤ��v�^�`W�4x�i���u�b�t�fcV���z܇2�q��0M�g�ے/��7�3�&[,�V^�����뮋��6 �*puP�@�ۂu���s�Ғ�]4�Z�)(z�J��rMU͢���Y��X���wΟ��rx��{>�{��+݂�?kt/�}�e���Q�g�57��v��#�Kk��-�pX��fH�����a4t8�ےCJ��e�^E�q캑�7{�2	M��*�r�Vc��Z|r�^a�e�����";��{|�I�(��Q�~���yƮ�?�֊y���?�Z������>e_Uh����q�Y����9�Q�N��~�Jyq�������HU�hmW�V���p�	-�����uBY@ż��K�@v]���%��	ު����v����mM��ַż�u�k�`���x�Ւ�u�N���pT�;�,O �ܪ�彭��V
)�ð���~U ��G��)tZ�H֞D����\��U��~$/V@����,�D�Ě8k���R1���0n�V� �N^�n+)L"T����ٍ�:��V�x�}	=P�U�����\�*��T��S7���?O*`���i����y��)���)+����m��w��g���f%������v�ͭ
V���R6::"*ٖ��c�5��酺��V��fZ��zH@�9�@H��<�kJI�tX�,���e�W�?�wUhܒ����	�$q~* c�ҧd��o
U0�8�;y$�6�