��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌ�'H�TԀ�YI~��\�4��U2�� �	Q��SPҭB�ڈ��@�6���DN�Qo�#.�j��u��(1U�݉ҟ�h�S�K�8Wp店 ��!Τg#�R�-)D��9p��8+<�oG$��tMB9��i.��g7�i������R���kTQ�.�]7����qbK9�Sv�Q��]�(�Amv�R�0ҏ�Kg[}������Qv��p�%���xf������!*{I7��b�-���C]U�Ԓ'0ޮ�6�]"�G��⦚�����V����Jc��i��ؑ�R2
jcU#�����LK�f" n����GU^�l��� �a����f�4z H�1�U /���!i�`3q��\�#��*�=*|��jf�J�x�*|��%�W�Dp��<M@��@Ȧ��� ���{I��i�5���?���,�pc�.��y���N����c���3��r��!2!��[�FQ�J����4{nD.�#)��0�j�_/�F��t5�4ֶ"�t`�&��\����9,��3FoK��{��~���֩�����5]yi�v�k��s�K5��49�lo��I�o�EFyyp�m�i)9J?٦��k,Ăm��$�<��R��v~T��*��XL���3T�5�Tj���5�4���R;k�S�A�4�y�C<k*ض2L�G��xfޠ�[��"�e�l���!�|?�ᢶ����m���H�8q>9E�H���Vv+�M4ЭT�)�Rn@'�������8o~`����eO�n��f�<�u/1o������"/��,�,���]����\Z���=QJcw�H}
nh|ňA���[����̄Ǎ����dk�ky��������0�*���ב�ua��w���j;"���O�6l8��4N@���O�.��/Y���������7�u0s2�X��?��&R�}X���F��D�|&�7�u��J���Ƒ��O<�z�|w��͎$H5�P�S��s>H�s,���J���,Ʌ2�	@,�䱄$����.��n���x�R7H�a��A_3uj�WHՋT8]��R#zT_!�%d�Nq��l�Z��	�1���P���NS��~��fN�����˱��G:TB��'\%�OI���k��ED�b.��,�Xؓ%⩽���Np��jdC0��4YH��+L�`��\�����q���`���D~V�`��	(q�iJ��Y�_U���^J�k3בb��a��嵷�8�����"L���A����L|��J%o����3ǝ�	��F�S�b�,��R�R