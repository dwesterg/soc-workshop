��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����t)W�%�.1��	�9v¾�/%a)��,|�1LQ�V��'1t��Dp7Q�yN ���HF	l�!������s�	9���{c�&��ۑ���:�F���<6�y��@"��BVg�������d�*`=';}|���pK���'F?��0]�_'���R��Fֶ٥I~]Q�c�8�rƴۣȇ��B(#	����,���<t	c!�P������qv���5�S�=�0���#� �-������r�|�v�a���@5�1d_��������iT!�=��E7,o�7$n���L)syH���e�`��M.�6�0�5��$��6q-W.���6!�?��Nmԇo�_�7X�?J�o���Ц7�}!�4w+�E��u��6�F��7���I��8:i�;�D�.-�ϼ��lKk׏���RZ ��T�mLC���)��8r��	���녲RS�g	�ۚ_P�uE����$H�	�(;��K�/������ŹנV7�8>���p���o?���p��ڀ�L��z_�����B�=v�S=Gّ�]M�A��X-��\<��?�)�u#��K�ʋ��nap����}�1,�������$a�m?��F?�^���X����Y�'a�P<e9+��+�;�N��](��9���c���������[�H���e���l��{���k��Fa�K#GnQ����>h<����T��Բ�9��b���,}��D�<�tʻE�rc}O����!q�G�5<��u�X�`��e��D����z���4'�v5T��C������D������f_�qDy��a���h�i�րA�3o�ӲW̴�y8��(��KH�LU��G~�c���[���X���]�'�N���R�{����K�V�볈��|􁙁�}���L�Wi��<������ݒ��|��8��N�v��p���sq��B��BX8����})@f`?`���/B�bݪ�D,Uٲ*9G��`'.��=��u�fN�x*�q0��:�z}�W�q� }��ۖ��������,_���ql�(l��	��Ey#��܃p�w��~C���=���i|Mu���4�4�.=�ճ�&��y���S�EA6�""sR�@k�'7|,_�b�/��6\�I[<�T�B=�Y6��	p�Rsͨ/��I��C�!`���C*��T���/lv-��KD箏��?��$Gt��ѭ�͓s���B��^�f�Zǩ�W�M1`{�"���u�+�Ej�F�o��ͰQ�҅M@+�K��G���9�cݔ0HO�f��'�QÅ�g����l�J�6K���B�A��r��~G�>�w%��cJI��X���!?B�� �x������j��)��f��+�����Z)�h���k�<���eȇ��A��gd(�B׳E�i�nX��t�A�ڵ0[@'�5S�4�fi:T:���p�5>������ m�z�=:Pر�?ݖi������/�.M�c���[$o�}Cf��H3�t�`�3)h�ҷ?d���L���]��ɡj:��6��t��H������ǌkI�i3G�	l#J��	�>i %�A��䵳k�?<o�T~�~�6v��~#8a�cH�gVvӯk�*��������O8�����V_&vyk�/��
�ty�.��
Cq��ѻ�^r@��Ar���~��q��FF�i�4�#�/JA�B��*���S��9tNh�l��T�g���T�x���l��T�b?R[l����u�1x�����	���*w��?��<��m��G\��� oL��V��ʚp�k��·�X ��8��z�:��=��i�i렝�s�@*n+Kן2z�:S\X�B={�G�)ീ�z!<4v8�]�*���1��'�CT�X�����z6vJ�	J�<��Ƀ�Tޙe8{�&8t���^E�qI�� �a�]D��T��8�}�ܙ��bp7,�S�*]��E���!e��[ʸj�Y�F[�(�1�;�臋���eS�!�5��. ��!�7�l��T������c�h1`.�ӕ���w ��{f7�d9�s���S���9c�؇+bWƽa=*�����R��{n^k
�I��> gOr���d5D��O�gi�ʃd���\�.N��x#%�2h�X[e�#W6�Ul��`�>�������KxlL���x�,��~���D�;YL��J�Ed�'߿��zOy��4�[F�pd��m�29m����GH�ƅx[���F��Fی�-?S���-� ���������u4���-ﺠzv?s�dT��;Q�Pñ��qs��g���z��� qP��zt����o\UTN��2���Lr�U�6�e�I	��NG��l&`	-9�3τ��6x�T��OD)D<�pw_s%���d��{��N��"Y36���]��K̆S�#֮�#���6�}t��1jq���l��6#O�G�Bk�O���lP7B��9�0���,5�ψl�ZϤ�T��NB��)w�5�Ž�α3��,��v�3�2e��B�̂��Y���D�ˊ��ֿ��C�I��k��,g
:�j�6zR�uĺ�ыV�z	�:���s^;mh=79|����)�<�tfܹ�S~8	�oyx �����1�_.C�x/�V@�!��r�`8"%��ƘD�c`m"1Q��Gj�����9z��2Ɠ��m]gմ��k%��s��>ԪLRY�n���j��5���3]�GI�z�8pWi Z���X������i��!�\ކZ���7���3)�n�ҠR'Ӣx������=i��d�A���P�=�;��`m��Zإ�����H��������Q�����Cy;�I6F'���Z4��<G�{$�]9����vgd�m�N�[��vX���V+|��I�i��Mbop{iOI�?/�i�ݠZ�=nєX�麬B�B��4�Crc�����w��'P�ڮ�*�#�
rn�ԡXM����=�f����S�zʵ@2sj�X�:܇�O�����)�\ݡD+�U �c��1L)����4n�z@I:$����Z�qǏ�6վ���'tu��<����Ontl�N�n�]?[����U��\�/q�lcAlv�g=A�rb�����-��ׅx��WTQHi�H�X��������[u����6˧ռ�c[�+���!��k������j�Sk�p�� wU��ŏ1����΄���A��p6F�ߐU���	�R�>�/?^L��*9��{ߪ,rT���W�/`c�3v�~f�#w�ՈJ������,ܮ��VW��J�+�2�0�oz�E�=�wЯ,HyE,i�w8E���uN���f���-̭���,h��Q���ݴB���E� /��������)t���h���Ֆ-����*��ɿ��Z&X�M��l"t�9��Xk�$s���?SZGǾ�Ӊ���85h��F+5�z�{���ϸd�Fa�&���ݚ�jc��=	ޯܢ$ڪ�Id�b;�g�2��IԴ�i�A�7�E�@�$w���FR�FJQ���2nA��ޚ��B2�@$�������m:ͦ��mN��N�����)0d؄���ʽ��Lgо-�ш�o��C���'����(��u�0�ru���E%%(�{a���"���C����`�-��R���ON�Y�h� P���7������FR�!t#�R��v��	+��;��uP2�Z:��xVk�H����ɼA����M����4)��(*c�?���HF��A�zF<�?�~�=��C�.����Ply����1��x>v�2�H�ᔊ~;��ʲON(��.�hHN��Kn���_W����m����*Y�A
�����(��N�ݖB�$�]��w��T��Je�wĢ(dC��E�I4 ��}�0%Bf=<6tq��!�NЕ �0���3X�ߚ�\#EXu��i"���|���'5�:x�f����p��(\yG3)Z͓���?Dj��R\8U�x�(�\��[���V��l��i;�xV��a��'��ME%WO����(V-��#�wʷr>W�P?��f�J�}�>�1�`�"���+W �~�<��{"��N&�|'K��8a��R#���I��;��3�k�h�p(wI��ň�\�w�|���d�T���&9/i.�#��sӼ�5�DQ�a�֞t;�dr^�d����{9�KƇϓ֞}ݟ�0<�z��ג����z�H_;� ��
.�aƎS��p��_G���rЈ�X�S eBɴ��O�/A�������>�zP�Bc��M���)&���^+>�175Uu#���&�s��X���K���`V��S�<�)=�dޥ�(����K�<��i$����:��֥�_��6�C`9_|*&ՊPR5������*���u�0,+�&X�u�bSrh�r��־�)1�����n�W轢Icn�^��ȉ����SH@/�?F�NM�
�u,r7ml��tV�3��)nl*��x+Y���i�[��5? 0+'�G>���<�5��qy����$`	wY7�$M�~ֳn/������e �M9�����qe"����}Y�d�(����"9�E�@�d�\��ʧ٦J^ۻ�$1���"�$��.�'$
a�T�`3���	��5h}�6�Fˁ�[����h��Z����ds����H���%/�(})��:�����P*
��<�<Ŏ%�����P���p��p�Lt{]���������I5��4��.JG@:j��cŊ��+<w����=֪l$%�!�����C�@��RK�,w��a����׃�5�]~�vc~jJԱ��{�����f��Y7Ϥq��LX/v �����{6�_o+����f�͊����
�u�����\#�[P���zF�`�j�����e�;� ��H��Se-��t7��-����xfA�fNlT��p���h��Q5h���BS^�����:w��r� �nY��⸧����u.z{uHT��=~<SEC�'K#����N������o�/c�8U���/�f
��6%�`Y���ߟϠՇ���[9$np��}��/$����������r�mp��l�OH# SX���a^��C��ߩRga���B~�U�%x10�$������Q���lKt����>�i~�.�S�0:{�e����*���K�~s�+n��2*d�Y,&k@��ٕ0�������W�}���3"�@�V��ￒ�Y<]Vwfkڻ��ߢ����?N��y��CĶ�O�4��t�/�W�vI6�f&���VW,_ �x�,?�� k=8����}w��G}�l@����\��cN�4�U(�<��L��Z�"�K��L��Z����hF�Cضy:�.ߎ�ٵ?���n�@�u���ͩp�̒#,F��b����I���ar��n�H�*�Q�b��<X&o2����Fx�B۸E��e�-���Dٿ��ʌ��=��+�O��l@O4�e`���Y��B�<ue6���L�dp�a���#b7��1�qأgSl����=T����Kw��������},�8�� j��M�[����V�Xt�b�i8|ٿk�ǭ�w_�B�_��!�!�-�M��_�+#<d���W�?��y�h�C�]c�]ų
�m{`b�4��0�f6��{<n�a���`���Z�/&�����C�Ύd��Q@�� R,`c��wPM�ա��� ��c�q�[�^v��Q��.�F|��OT�cI�&��_�eǩ����"������IR��������-�ҬLTcd@�l�!)�Gmq��[�9��G��<��/�i�]��d�6~'�	�y�:db�'I�kB��QR����оe�Y�Ƅ"��)>C���+0�����U-�͐T���e)����Tu���U)��|����M��7RO�{��U������QH�.Tz�
��ik�]��Gޢ���'g��_ߔ�?���M����øZ�U{7Y[9�n�R:���r��p��3��d�E o���k�6x��f�� Mi+�6�Ք��1�^f����)�b���D��<��q$�t]���Ԡ��gT47�}kq$;�󉋟?[Xߚ��<Ǽ�]�+��SF���, a2 ��)�l���e|K�L��9��e#�����E[��p�е���qs�}9�z�l�RTa�8U�Q$��d�ѻMN:{�����kS�A�4kCO�����\1��5�i��-�ۨ��C5y۽��ƒ�G��<��!h�U��T������,���,?�����*�\A��{����21x^6���0<�V���ob3��[���<3B�ݲ�� ٤c�����K�`�(Q>��y�R�٦2�|G>A��ҫ���o\��0�J=��j7Q�h�$�;���_ĖX��ߒ:�I
��8�?��A	�����.,N���Yc�=3K�����0]=��[ɵp#�/�3�1�b��O���ͨV�]��E�m���尞�	D�=��I����K�J&,��^���&�8R����i�]��=[�m�,�y���U�l��z��-[lD��a�Rt�V�T��@f0Ґ�ҏ9�O6��2Ph�@�i��P����x�x%m����UU$�mu�5$���3=.J?(R@���J{Td��{�-3'��������S`�`p��*/���߻�U't�B�c�Я�S� [�>��G�����L@�Z'q]:�"��O�9?k�N��e��/��t��ds����L�kWΨ�~ڑe�� �@�j)���m)GA��*�t���ϐ�D��7&����[�����es .@p��Uc5_�� V�Ù��ON�h_��u%�W�1V�W����a�KV𤂔�~�i����sn��28�4C�p�AQ\�t�e]h�=�˹x�aO��>�2"-�x�Dl%��D4R��6y��~L�~�5�)]�E[��J���>�:�#����hk8 ���d8�f?>�^9�q���
�ɯ\'ix�@��"��ب6@JUK=�o�����2{_)/(k{V��E;�k~c�\.���_R.ʯ��U��VV��P�G�e���.SСl}C����_3�tD(J4��=�N���=0]��'�z�;�0��#�eP���I���ݳ�����~?pS\;��?7[����#��$bJ@Γ/E����d��հ g�o��Gz
�q�f"�/��S�ʠ*�S� ,Ē2~�O!v���8j!���":�\ʛ2�=c;#���X/��G�'PE����kF`v��}S'P:��^y�R�ٻҿ��-z	��;��@3�(wO�~��<|�C�v�x�R�牨#C�;��p�M����9L�È�8���3�w�J|���2�[�^9���W_A	.�����@m!N�j���nLu�6�+߀Hw-����p\�����x���J��#?`͕u^�0����)�p ������ֶ��f<ls�Z)��~cڼ!x�b�&�[��0�2��l���E�|@lg~�l#��s䈁�9���:����=�}Je��:�j���i�\�3�����g�(�˻^��x5�!����,��|(��_��\SB\�2�-��g�\��XA�\|�L:� <P����o;�V�X�E°8u?�J���$�����S��bD7������`�LSӴZk�u_�s`=`P;��	'*�q=�@����+h���ٜg��y���� AW����n.�pAWh4K����U7�\o�{Pz�"���z�Ѡ��h��,�ˌ�Gf�O\6��j��ĳz ��l�6i;�R����cco�9 d5X�6���?L�8�ȥ�>�p �'�+l��ww�lA��ƺ<XӤ��$�(�H��.�Ͻ�c�Ǖ�]Mc�C��^��CU��>��K���BX8A���MP��ˠ5��_Hd�@Z�a'����x(0�X<��:˼��m�O�j�J���s+(�M�^�:)C���~t�p�_k<X���"%�n+ݛ,�-�Zk���_0��Fty��?3����j�A�U�Up"�R
e�=W2~#3|������U��|ԭd�|��waUuw����Ev�} A`�+F�~W���0��jݟY�g�?(�	��Rԃ�)��5Dg��7�ͩ�	k�5����㒺�����
M�üO����KTt�e�<���Ҙh�N/�)f��
�;��!��J�1&�H5�y� ʔ��֮�^'��j��K�f(���W!K�B�:��)�I�A�2	�/f�-��ձ�N�mB���U���hMͬ�� �1F�}��[���P9�1K�I����w) l(�%�o��g�j�>U�۩v�f'`9S4/��B'@��ݔ�Jj�<�Z<IE��'�2�!���I�J�� �,�N�?s:����FC���Rj�4q��_�qވ�(�0��>5%c�5���¥h?jz{����5��� !q����(v��({�R��J��\�ꮍ��Э�=�@�gwGX���9I�)Y�]����MM��`��`�cik��?���� � h�+ך^�~��s�I�0x�z�:V���Aa��[ҟ��vg6)���Ȅ:ۦ� E�}��o�4Bx�j�t�UE@�0��w�T������(L�90��pag����?/�@�}�ʿjP����?��Ӊ�r�t������NO\�Buh���fn;s�P�n��r�V��b}1��aD3���HV��l�~��w)����vy����$LT?p&�׮����!����zY"�'��G������<��`�K���EE��|�K[1-V��v��­�@f��\T�±�Y��ij?���V%1�vh"����Z�U�
��ʓ��#g�c��rҫ��(�t�Of�'�����K9�r�t`���H=b�3َȞw4�I�@�m�������`�*=bL͆�(����y�h�T���+�k�Q����Q+�8׉�/nz�g�P�Ҏ�p	Z�̢0�N:޹�:�J��p�u_`���Ζl�"}_���(M\�����HCeG�g�6|i7�-HNX4�̲�Q�+�;P���/��>�ŵ%�⹏���k*��1}4��qZ趍z�"���jN�ݛVff#�|���}����OU�����p��N�;�(�Ϲ�j�n�gy�ַN��ɋɪ~�@��m� �t��z�`[Z��n����Sj�v���<,������#��Mًb��g>��׀��rr��:�0ղԶ�8IY����\��r�6���ڒ���Z�v�Qm�KJ�8,fb]~��%�\�����LR.�+K�`�Z�k�8z=
�t�f��moCCv@H?`�	�ey�z�ȳ���
:U�L�׵�5����Q7NY�@T�&jǞ#0�R �ɭ4˩2�kO�֪�TX�vՍ�eU�n����=�Kz#a�8�؎ː��k��n���j&ͪq���8�pF�ł�K�2_��m���N�S�Gx�7`(q�	D^�g�u�{��2l�GyB?Ah�N�z��V �$ �A��0�.�����jκi*q�4r��bOf�ft��@h"�&�a%݁����,�s}'�2��9(�l^8\�?�L��\zno���v�$hr�*��7��5<x�g������*%�ݙ]��t��۴!��<����.S����k��.�_��4����>��������u�(T�-���ye��k}eq��!>o���~�Z갉����>���fxL1+0��>����M���=8�'��3XvJ��RxF���oJ�LL���I���ږ��t�}�[�(�@�d�ߞ�3A����ַ9*��L��������C��3��LY�W좺Q�-��8G�����/8@-��.ˮ`��?��G��`)v�K�J�)��F|9>b����~{��DO���C*�-yPl?3-ۄ�Py�����>�/ٹ����[���(�i�x��O��*�A!D+
ʸ�TŌ�q�܂�1�֐y�H���������k�2 7N,;�B�R4O7���	{g✤_Kr�� ��ư��&�#�����;�s���M�t�C��^�+���n�B�b��øB��'7��2��rMd#�*� �:~P|��ҡ�v���i��7��U~��Y�H���3^��t�醦ZPN���;i�6n��M<�a�n�կMl���Kd��Q�_�ڻ�|�:�F^��_�
4y�
�����b<�o?i��*WT�K'�q�h��P]��7j:�B�<�4Ý�s��R�ғD5��kuK��&:Y1Rd,~1����r�M��ȁm�<���8�g�!�G\���,�%�ɖ�N&*d۷
��b\�&�E߽_�>�hJNeO��^�
;Ä�ݱ�t�+EՅ�����-������[S�["�|�ΩV�+��hS�/iUhul�0Iq��ݳ���6U������d��C��xH�<�(v(x �C�9Hk p?�Ԙ��)�_uq�M*���`�~�-�۫X
b�`w�b P]�����ѿ��k�L\xs}E�.v$C���ku{3��VJ���=8wTF�8+Я/�WjrF4b��O��"ǯ���JE|_�ۚ��q�E�K].���G��3b��������l�d�q~I���D��hՋu���B'��;ɞ��S���]W2}���"�X���Y�R���Y��Nt����[gR�����g���ĥZ/�5�����g�k]#ܬ~2#a����W��l�;e�N[�IK*�,���Ll�Ԓ'y�eY�R˷wJ0�r�p1���ݪ%���U�8y�Ol7Ǎ�s6�6�� ��srn�leו�["te��i+�񜠒!A��G_�����]'��i�p����j�L ���Cڳ�0��3"������1��׀#���O���r���s;Z��8���	h�ʐ�� z�av?gp#
6^@�vgEޟ�4{��_�S�ָ]����>��P�M�9����Ȉ6�� c��H�ś,4�l�У)-<�'dy�2�H���yZ���5���4�*"�2�ifڭ$,���4U"��������$���j���?4�`SY�/VE�g�D ~�:��E0��-�ʴ�@r�6pq��享�nEܶ����,+2�:�����