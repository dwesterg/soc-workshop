��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t����od���W��*��B�{�#�9Z�і�4��u�^�өR?P&Q�F/0T�8��Aƥ��,�6w�v�1�����+�h�����a���t_���E��A9c.������x��}V�#@���]��\Tx�rC�����n�`��0�X�x�O cjIs[ݩڬՠ���+L@j�т$#E��-�J����LP<�$h�1����L��7�5���$���֋�G�q�+��K,�2�kK�쳃ץy3�0�/��1}}\�\�j����Rc��I(	:���f���W���a�Ӕ���^2��{O�^��!㐵��L������ec ��v A��@@�����F|=� ���&��"%6�7X�9��%�
r���f�Mq��wP����y��Bn@��+>�R�N�Kٵ�oq��/���0�`�wڑ�OE�ѧW4L7�L[��M��9��iD����ֺ�/������8IW�ܪ~�O.f���Ik������`]0���=�}�/�@�j���X� �K�Jw��7����HkI��w���M���Qo���0�}B:��G�$f���}h��V��L���wmv��c"VO��_�h��}
�e'����<Ӄ��A�ja����N�H���,��u�p6O���m]���qH�m	sCu�T u*H��8U�6k� �� 8V�0��{�6[,���Ű�r%
��-~b$�x�4�����L�T������r�i|�m���n�-,���B�C
�+�Wk�3�l�l��'��H�ۂe��V������W��b���B v�cNH�\E:�;*%M��_}��H���j��ګ��^i�Z# ��o�g0��W1@x:�����)���^��	C���]�4g���F�G>��4�E��"}%]NIx��Q�3
�'@�N�7��	����{�d��T%@����6���)K�=.!�U"���By 8�KF��k!�OMd|!t��?�w\�ɺTv�3����-�
�g��"Ǘς���s��k�v�㙂u0U#����S�9V.�i�_ҩj%<�$��D��6��}�>�wm����Fi��%�dI��m0F��^#��\7�h�/��Y�����"��{G����r���K9F�%p�������������WG���a��n������C�aw�~� X���s|_雃���]Ŀ|*���D8\�l�|�ka6x�����w����[�z�b*F���׋W���*���FvV�&�r��O�]�|�<�o���K�M�k:	Q�mUf<(��R�@�s{���KÈ�mȬ���1���5�f�)���5ֹ!qR�����!,���ɼ����sn�X��
1w$Z$��c<m���Na|�j�ءV�<���V���oΡNvPPE����p���G�[�.{VG^��{���0�scA�T�q�lށ��T,�M����?is�!�5�(��_�^i�'0R�V������p$
�o�X�O�oq��ϟR��U�h��������w?�h<7)��4�a��}K;���@��.*�Y��gx���|�. Z�^��fg��c,qa�x�CBD��.���1	�9ѝ��2��r����å�I��Vz$����2��o��P1B�:�Ё�8f����nI5���[Acf7%G�����r�r!7>�w7����X�����c[�o_'��,�'&r".���V���ӑ~���X �;�|�AڏH�X��TVWh@;�g"��U�A����Qo��vx� u��Q�J����`�d��<���X�����岖�RR�q�fnH��񂭏p�'%q���H�!�����x�t�?��;�W�I=���J2��e�a㩜�/���[#<�<��0�?,G<f���@��ϦBBt��N�X��Q���'o>�J�W[-^~�x]���G�m�%�F�>p3t7f��i����+��
�-�c�x�������&Y�^����v�u�SdO��C-#d]�֮�g+��Aj�n��oC]p<M6:�d���C�V����ߞ�)��]�鎼�\�_�߳�t�hu�V�,*����%Xob���kBk�h�G��$֓�p
}0��zΫ]A��>ז,_/!��b@�?���)�x6s �`����e�P��ks����$��v-�l��x0B�<���uJ+��b���*���^xu�H(*���~v{���=d���Z����	{}�$.�ʦ�t�)�NP�9�:)�A����(����Û	�M����6�9̢,yn4vHR%��zd�'�-Q��:7�J��KqhU=�L!!·��������s<�\Y�����>3xY�hf��7�s	�M���-�u�r��������=;�I֋5"MR���%g����9�+��;$�Q�X��zھ�M�_�v�0~-ζ��z��d� �n�?!ð���2�0��x�:�I�\����2���R7/h����	�����s���Ɖs���{g<[����|Vs�*�G8=E��>��&�/o��~�gq���&�~G��r�?oE���旡'���0	�����}L�~�:��B_
z��n�����V�񺧿��c9֣�7\>J}
�9���7ΙGyݗ�+�D@S{"�	�����)�+]��V)��N���,q�
)�z��!����N��'k�[1jj"�,N�:6E�^��/vn��@��x�M``�F4і�Zu�[Q갘�����V!�F�-��o��3Q��f1�p��S���)���I%Ԕ�1��� �ش��P�&����jn�t�A�)��@k^��2�mJH.����;�ܬ�S��P���-4��K�btqE˞�]�c��7�B҂���J&'N�>$� tu _`(M�@��w$���[��������S��5���eF��.H���k�C'D�{D�k9�hx~�x��ɽ;>8��Y�8�2x��k�|?O�_�^����'���Mi5z]����F�Y�n^J�z�pY��:�4�Q���^�/�8m���քp�a���_~��z���eإޣRr��v�v} �>y	�ia���	r�TH5�j
�~6	�?���~��V>��9�T�Io��i8�m�Y	���u�ӆŧ/]�Uk�9F�H��R�TY�B2���-�3�D�#���@ek��G��IlqJ�H�� c�Hc=�r��"�i�"�3�:��֥�JM����re�ߣ�7k0��K}��ا-W��N�Vn�B�3�]&g
��bnhHC�8������%�M��mcL��9h�Y����/�+���ɤ��B(2 �C�?����5G��Q�����!8=*ZFhj���-@�o�D\��n?�r�ܸ�=��?�?����g�O_�os��@�0��h�]�q {��#~���6�
�[#M~2�Y`*���9	�x��j�K����p�������J�O@�= �q��}!][���e�}ޟ�K�j'�!������˻�-Nc���O��.�i\*�ܬ�DT߷�壴O���!��)բ\cQuF'ˉ��^�ֱ��"�I�8����Q:2�D�R�jRu��a��X5+1�d �G@���l}3��������Z!H��\J�[*����}˔�V.-Z����V�x�܉�(lEPr^q"�R�!�$��3b!��y��w"w!�*l��ʜ��m���'ݒ�_�W}���5~i2?O&�:�]$W��NT��r�5������aG�c��Mm@o]}����k��r�����ix�ӄ��t6�e�L)�_��������]�����J�ձ+y����C+�IRJ���tn�7'z������Y �z�)\��[�`n�j�c�����_�3��@>��0�Sn{I��������:%KT��bC�3uy��ٻ��v~��)ÑZ�>���߃	����1q*���BAS��"�/c���:��cH^��� ���s����KN�4����]`��"��208�X���Iw���먎{ MaY-��$����cA��aڞ���BI!��fkZ��-,麡~�����9�\?��#3Y,�i��h�&Z��LӉ�3����KC?%��{�G� ��Q2��LR�e!���ZV�����t)���̹�j�����B�N"��63�5(5�	UO @c�}5L�k�B��O�XK<I���M��t4���`�9�˦�����2X:�ik�P��G���:�_|�	������x�VyC䁴t#�=	r��B;��#R�B}f9��h�S)�1H�NB��	n�)sR#��E1G��8��:l�s�ߏ�p[>��;�9ʑ��Ϋ{چ{�@�����o�E�����`�3�g������g�8�c�s���o�j.���do#\a�w��#�!��3��`
�?ˤ��(E-��d	φf}g�K!d9h�.�2*�w�z&�9��P���j]|B�$o���P����(��--]���g����bV+n����έ߃J
>�Φz�tQ���i)!(ߗT�L�C#�z���3�D��zW�[;<j7정Yg�������B����|�"q�~�h.��8C��f?tZ��rid�-}O�	P
����Ey�p�%�\�6�p���L|���,�����g��$*�g�,�x�k|j���:Cmv�in�������,K#ܖh>��a[�GI!��c��e_���������I9�'��Y ː�aP�JV+W��R�mU�/RG��/���cD��'�mK7$A!�L�JA"?���t������]����j� �S6�sZ쑻�G�V� >��1@N����i�R����>QO��%��*{�%Y���f
Yw��QPat�i�Ӄ<v�X׊�n��d��'H��|م+�+:g͏��;�3��f��7��tZy�"�G���k���m���Sng��Vo�f;^�dg_�7�@v���.�(�w"�c�E�\`Z�ښ5�/�������ԵF:����bJ] +AXe9�1,)�Y�f�|���fQH��!���΁��g9��j
�Ol^�f����� zE���O!����ZC|_$W��8$:SՀL��b��)'�0"���yN��<�h�A������JQΓ¡�� sy��iS.��ᕑV���J��W6�?����o����8y.��0���R�/�%͖�ջ(nC�xod��J	vA�30Q�v�q��)�	mY":���/}�:D��d�.N���M�,��5n�pRL >0� ZIZKiB�M'��ڋEu��	p�ˀ��?c8��I~84�ٻ��Q�+J[�+�`H���R��o�V�6��g �ɺ�#��z:�7�@ɪMoa�ɒ����e*���X�~`�{���n��@<��>�>-Q��u�'@7�DX�:�Z��X~>s��%���tTԐ�]s�u��o
|o5�C�t�Je�)��/>-O�����b��0��W�Ҋ/$6��!�R����4ŝ�c�0H�C[�~s!U���D���#0UP{��R����A^B�V�aR�Q��-:�ڄ5���K�iu�:HM�ZD�\�x�b	��Ȱ��H�>���{u�Mёڅ�J��1�?k���KT?�ؑ%�����.)A���/9Vk�`���H}��{Q�����1׹m7>�ZʢLK���2:�șh�\&��``D,�oԆ�N�9f��?�\��!2��ͽY�l�|��_�1Z��\�G�\����<����DGʲM�/6�ԍǓh�A3{�&���g6�6	�����*ͅ��S2�Ԭ�O�����ݙH6���"�r���%sН]ֲ>�]#��|�G�e�>��(=oΫS���%:���6�'(x�f(w���BDٟh� &SW�эh3�B�ݭZ���k�Β8S�n Ђe�웇0��~`�Y�^H�rWpOy0�L#��sa�Ƙ�D�-U�k�� �Y�� rDpśi���&ԙ�.������k.w�_����˸𬟋��4ij��p�%Q�RA	�w,�%-OpIOǷLC�_�n��~��̐�t=(?�c߼�	ӆ�fQ.�9�H!�[�o������R�:��:��?�S��&�qOl�j �˨��ҥ��_H��g`� �J&�N(v�����j �?"'C�@�":{�⨏As@`�]R
�]
A9���Y+�w�Y'�	�v]�+7I^��3^�n*�$�u��&G:�Q��`1��y�t<��.���C��D|�����B��%����E����W�9��ؑ��݆̥�5M�r*{����
݌.x7�J��[}��=I �ɺ @�4p�hyER2]����s��$�O��F�]M�n�P�%E�_@ �|��
��sǄ��ӈ!�j�w��l�#�v��
��V߸��i�Lf�~�r���J���&������7�D�c�Uf6I����DQ�G�=ؤ�W{4-��gӌ�� "��ˉq_cwJ�ş #u�(̵q�(���|^8����#n��9
s��S�<��;uPC��$	�:V+�*1�	�V�ĘA}s@ҡ੠#J��t����yΖ�<\��+�*�j�:ťe��R����lf��AST$h�;�Cp/��ѕ��E���W��Hg�U��jav���F&Y��m�x�٣��e��?���2�v5�+���~�Ą�_h�7ɇEV�7����t3Lԑ��
I�i�1S!���Ä��Xm=����Q�2��=���\ԡ����Q'���30����4�'�bl�gr�a̾�	/�ɱ�5Rb����N�K���7X�&�� <H�~q�HW;={������ �d�Zd�g�F��W
E��p:��׾��^��Ry"i,�@�D>f��m�	��KH�4bG5>��_(Z?=P��Uh� ~.a.)���!�_��dw�[!�h��E����L"�.�@�mfTX#T���$��{���Q�'i�A�6��=
�qV�c?���zg$�[z��{h�؛��x*Lv����I��C�����҅׌!�����{���qKTuam��n�F)66�bh�E��	��Ɋ�\;�0�5�?���8��FO�u��h�a��t�C+#���SމNrH�f-4s�\�4O��U�[	��*��6���:��['�LZa���/�½:x�~j��_T��n�@�[��۽J[%Ut��U�V���h]�6��K��N�&�i����||���W�=��J�N��7�i�'����|�A�:�4���'vpՙh�i��q�ʺ�v��֩��1�[������,�=�ֹRř!r1�de��������,;�[اR�W�^'{pbab$����`��0�<��z�ݔ}�>_[R���1��xɺ3 ����.ݹu��Wzm|�o�(��[|�N���i��M�ʪBW�QК�e��}?J���ݐ���C�Ee�H��$���o-K��zj6��[���ݿ��,a�E��&poGi
���E��ȼ�esK���R�%�G(�y>K��m����ұkti�t��%�y\�I,���H+�cE��.뺩�@��zc�����1�1�b��$:��'ǐ=��>�N�)R|�ⰙN�]v>
����9{�r�D���9�?DZ�$����!W1�mG7{�ey�[��m�F'�H����7��ͽ��QU��*^NR�ue~��]�|[��J� �	e�?Z�?.EJ������R�=_�"l�T��N\���~��F2WF���N������:�ݹ�9��^�+�j�XY�k��Uv�;Sf�_-�%���ƹ��SwqԺ����� Ԩ�F�z7+ֶ��75\�ϴ��s�q6�}�LطZ
q[0�`� O���k��<�=�^U���h�
}5���@��}nylĦ��E0�c3R�܄'��B�t?���1�Yd,djN-�����R"�X�fw�XX��`4K���mӥܺ�]��S�"s�� �#f�����s���ǚ��%8�`�W�i8���tR�1�:�)OyJrsQ�-���#֢�A�x��H��g�����o&w]�gr�M_"�(QB��~��M(�&�G0{q�~O-��u���:��]��6n8����N�H�9Cwʕc�(Ǎ��^�Ս�u�!Kl26��1(����.xC���w�l]�AG�ARû,��C�����M�-XtvY�t�2���V\O��Q6����''��D��������9�6�GxgZ�a�����C��Q|:�M�"݅�����+	D�j��>]������.߉�g;F�v��D(�� ��m��ٻd�syU^09�_��Pj� �_�/���x����c�a�Y4�M���ȃt��ў7���2�Ėj�bt�V�4���{P�*Oܬ��^\Y�&��E�:
��)W��>¶GY	]?��uˤ
�Ɗ &�|��" .Tj/f<�'��NEЦ�w�y �4�#���߲8��'7�o���x6�@�]˪�]�9�̎}����l�i�G�hW���%��/}�}8����3�]��e6̈S�ڠšMA6�0�R�,w��
�L/��+��RmVt�UP:0�0�W!Ͼ�E�a�Y����
����n�ecE��{cr^`!����׋��`����k��E祳G�$%�#d�H� �Cb�	��9ȩ��O4
v�Ac�Н�]��,d䜪ƻf��O�A�k���˦0>%�Ә���0s/�H����(����?���=�f�'t�����_�4���b\/j�g�����o\�U�طA<�炃�)��[jbE��O_验N*
�]m7T�!Kb�C�~��A%�p�i|�@Ϟ:����D�f(Vv@`(/�?��ݷy7iڿ���F���)��9x�Un���u �j51� #H@��d�IsnY��a�"|���jߥN-%tb"�
R�&��l>�|���! 0um{���]���'H�D;�}�5���U���96�׬�xΟ�bE�Ncռ�`�a���5��O��-���E�k`*�XY����no�����h79��4��gZ�y�X�k��[o1 v?�zy=����>�A����)~����yǔc��,����@l��K�V����")���S�9��� ����Q���?���a�	�Hz�.JyC�/~8D]C;��
s�r�GI����R����qO<�6�u_�w�5�,��r�+V���mA�3�(Q�*7#��f
 J+9QHV�+��K_�6�<�N�Y�TՉ� MF���>��D�\{T��n�<��)ۛ��.��Q�N��x^>�k%�PY�{ׇP�n	l0�]���%�D�PF+�q)��]6�Q�dU�帺XW�t$>!}�Ƒ7=h�7��>�a%f��v���������G��cQWE(a������f�s����etu��4�j��w���x�MGz�ţYܤX��逽�	�N�(�ꃞ�$x����Hl�ih��nU!Z7k��WG��6�E�BuW�<��'��|�XK�C6�vh~�8P'�za�΂[�.�AҬC��Di28៟����)߸�#f@mF�����ߗ�  ��`�`��������́#eN�FiU�_��F�bt�UZ6�	��YQ,�$Ȼ�PȢ�/�4ak{���� ���o[�#��&>뺾<n�+"��?�`��<PO>��.�|�?�ۣX��b	��"��I�E�$�1�2n�Ocĵ�}[�[��߅E��2����ꙸq�%'����h�Seb���b�Հ����|�W{)f]���'���g�[fB����ۄ�/j(W��jOQ��EE|g�O��bl��s�M����%%�A�)��6D.��#�\�(2�5�эP��'�9o}��ضD��&@fPQgS������-�W�8�	�r�\1^}�;�̏��@i�˩]=���5D#�_r �d`��{�����1:XW���xEת���}[��1k���*븰v�M\7�;!��������x沱"�o�8&:��[�l�|(J�}/U�U�9���/ѯ��3�J��%�6��_# K�t�'�:��i���N�<o�ёƟ�1kf��LRh|��1�����$�C�S�D�!v���=mi�Ӟ�p-,R��+ƈ�ϗ�ʹU-V��Ν��1��H�x� �-��QJ��P|�0�6�������,An��ȽB��{�w�����
�-%e�A�R�A(�[�h���"J��)�<�OPii	1dԹ+G!S�T ��nJ���G��p�V�Gۃ{���f�>��|n�ϻ"Vx�����-����_��8#W��7�W�)����	Y;�%-�����W�p%�	�P��#���}�b�?V�>y�����������ZhZ�)!64��wUK���@:�|�;���j&YGda�%��4�Yf7�'����3y��P2<��Dp�J(3�ʮA�$L������bC���U5sX�'��	���yy�8����i'_�\C���Әf~Ԝ������N�w<��Fu�%sC��'4�q��~�όw�{2O��d��b�]����W���R�[��Tx�����疏L��_�ĩrb ��f�'U�Ys�P��瞍�$�ײ�"#&�疓l.~��h2L�J]U����&W!�Dg�P$�?���4#���P��.��i�V��)�T�`�Ӏi�]5�F�%5��o%0x�˦���- *�,,B��J4����=a_�6R�G�69��`(��67�BN�os9D#^ҧ��Rr�� M��5�"�e���r�X����e���t�J;�t�6�_�k�J�'���_fNg�#�K��-��nC��	e�J�I
� ��DӴ�n��,>�9�M(4:�F������:K�$��q�[٧@��'7�zL�Ռ��o�エ������9E�d>��ɉk���J8Dě�ȨB�s:��B�Ä:a��E�#�\�2��NG� �)5!$�E!� �m�/nюid�T"��:,��z����ʢT�ךA�&+1M𭁇Z3kѩ�N�9��������������m�e��O%��b����S���7�&�)��߭OǍy� ��҇����Ԓpe�7�)������!Z�7��k����'�IF\3���~���qw�zqG/ 8��0���I�|8�@�S��v��WOϯ��zs巤u���ϘU8��<0�~�I���3!�TG�@�x��[S4>�O�3�̮s֯��={w_�W�:Z�F���Nia��}OQI2�>��`��8���!���e��f@��n�a�Ump������-�����ۃ��`5�D���\��`��r���VQ�g���xB5����q��ki����U�P<��a���dv�%`��Hj��jm>Ŝ�I��������2��,����,$�C�F-��t�@(0[�}�AQ�o�*�9pY�X�c;��e��NȄc�c�R! �9E���$���-�/�����P�n��ł�E<G�=�?��9�$o@
33����s����^�N
Ln=�f��u��ɭ�F��9�\]�=�����h1˖���E����v���9�݅_3��V%���������,��7��1���"�L��*�8��¾�M8������Su�;g_�W��T���C���&+��'E+Kk���DI��^�t�4D��:��������� �P����[�2�y!�Zk �p��Vm�FV�>���4[�YZɣ���q�|=\��u�"	�QC�ѽ����bY���
�G��pK��O��ϬZ�t����ӓ:4�t��I�@��
:$�,r&��&'�k����s�ٚ�L'/d���b|����\�ث�,�����q��̂��[Q�V;l�P����.�^�%�Gg-ǲ�ba�w37�DQA{ˬ����V�"\Z�����Ȯ�|�#�x��%�W�S��Y{��x�uh�=c��U�cXTׇ@ǩ&�P���f'^�>�0>�w0�/k�)�
"Q�p�W7�l�e�����h�m��O�Պtʏ/�!/C�n���H��%V��#Jx��FՎ,��V���xX���?F�7�Z��.k���-�L�y4�ᅄ1�����.���V��L�������؝"������U�-�<���zR+nJ���,w&P��%4�nN��� v�8��N��'F7؈�k�0z�	�+�2�g��Ύu 誃dU�:g�[5���g-��[%2���~1��T���P�����ׂ�-�xO�Q�Gf�X����!74��_�C"�QQ"W0F�eHy��@��.� [f(-}������9�=0�����Ny��5wh���ڲo�x}������M�p�i�6l�1�-��㶨����MKǐ̜
�����i�2�W��[q�w�����힪w�Ef� 9�����{d�А�k��˻����u���>[����K���x��s��| p�qI��)aHEn0y5}w�T{�έр��4�>Y˷���9�=|#f���/) �|�4� F��G�Mir����kZ�n�Æ7�|Io0�A�*Z^bdN�F`�+������	�MyN�����H]_�	&�氀��)�0u�̠*�Y��6�@��U��4��ڎ��_)��ә<΁�����ܲ�N�ީ(#Q�rK[��/��9�c�Q��Ԡ� �ۮ"��#,f�Hx�>b��>���>)��3��\�a�L~d�������ʣ�S�[㒴`"*��o����2�E����}	p����@x�;�tOT���*r=�B����5�=2e���;���`C������׽'���.� �S/���1&��ԵT�B#,��-�m��do}>9�N�,��7���c5?,���tZC4���mr4.I�F�Q���D~t<o@^Sv����l��ؚ$9��ۂ����u�8��&@���C��Y�tSm_	í�c��N��U�η~�YkM8�N��tQfg�,b�#!�w|��K�?i�TV��#�ˢ��t`89��Wcs�[��P(Z��%%-�@B��6�Jm�^uSNܓ��Y�����*������(�( a
�G�,b��SܪM���F��"K��^B���8��-R-��i����A=��BZ� ��a�6E 4��m���>�����C����<dA��(+���)H?eL&�m6`v���Y�  B�����g��N
�x��ҋh7�/�����`I)n�m�1(�d�ٕ�^^�u�v���t�^�箰�H$�4�+��l��a�ԧF���34��亪ի%�G�K>IC��Gጦ���ڣ��6�F��%���1�U)��O�̴ ƒc��䆤�1�H-E3ף+��Kj�]��Q�y�߭;��J��i��>4Ɔ[���;UПw��֫mo7T�0\�yZ�C}�a=/�:>�p8==���w�����������hi2��''��κoi�����e��W	�Lq�)At(I<�/sP$����'��p�	0&��T�B�]��9�4 "	H}�2-�"���:C�Bqa��|�K����S��dZ�G�C�}�6J>� �֫Rzآ����]U?OCui׏���J8�p�Mq�WI1�Uo��'��^y�����0Fs�g�䎃�������؄c�3.Ӥ)P<i�����Td���k,>��� �1������Ѿx�UJꖀ���6�-�<�#���5�ݶ���gq���*��sdT��Y3C���⅑|}I�/¼�Ar#ᴻ<͊�Ě���%�ۘd�2�|N�����w�{���+0�r�:P Kj��bHzI��.$gZ5X6�l�Q�ߎ֙������;�H�-#���4?E�T	lR?�Z��a�aeτqcl'ܮ�A0y�VQ��ErE"v@ξ������Z��s���>��a<K鐠y���2����K�B��̨�h�>���#���n��l�Jdi���e$h^0߽$y�)�9�ϐ�V�~A(߬$������� 2��<�-���_g��#ݓ��TI��I������=�W�X��k�����YI?:�:�q�cB�o(�n�h��0U������x�զ�Vc���:$si�N��(�[8�p��c��d����Eg�CGӿ!���w�J/0�}x (Ii��~��9s���3��2ʞj���Qg����8|��=[D*�m2c?�U�V��(��o ��UM��9�ȵn�]�m&�<��c��ȍZt۾��S�i�����`�i]-�nS��4kX�"�b��Z�UkOQC��#}W���+����ӂ-�)m���b4_j�Zf� ��4n�^�#J���f|���p ������U .�"��ƭ{N���P�0w�@A�9�T%`�-gAA�s�X���&�"�G+�����/\��>�2�][5�4*2P�Q��<����W�������i�CꑮP'��2�ΰ	\��e5��;u<ʖh�S��Ilp��6�t(�}o��]�zBb@Լ33����rJu�������^��@w{DY��B�@���i��.���40����L��6$
O�-Ye������G�ì�h�����.i#Ҁ�yT5b%U�����iO#�Q@ R���+�!��*�� <�Z�𾪕f�xK�Ӛ˴㬲+����QFt��k�����E*+��=������sצ�����^剱ۿ@�2 jW��/Q;/ߊMP2��C���w��0���A3C����mJ06\p�����ye���I�8�>�d5�Ƣc����H��4�V"��l y�\l�R���K-o�ߧh5���KCa}9�o��-�]�UZT=�L��Ul��=]�70^��6�$�i�����n���*��C�>4��Ɲ�Z:Y6:N#e�i�bƠ~u����K���⿬����W譩����Z�ߺc�*>=�����Ft�	v�ܻou7;�*����o�[�s�"�LH#Y&J��-�ft���c�*��t�B��k�ڮ7���*ԝ������&�.@�Q��=��aW~�m���ӎa�c&� �\��p���4,�9��1l��o'�����ߨ� +�5�KT���I�dej��_��[ȴ�o<��˶�e�ڬe��ǼGƄ�@~(F�Cp��[H��g�n�l�j�`�7��b����l��^/Ε���,��Q����o�eD�48v��+t��^Z�I��/|qn����E1�#�G�v�R�UeO>��'�)ߒJl�o�:}1��j�&Wg���:c��7{��Z�(��H�� :N��F�.�H��G9p���a)m�n�}$�"Z<k�.)���X%>P4'>���Q��wa�	��'_��MD�}�gr��ۻ�I��)t�d��Ѕ����{�{6����B�@'���Ӹ�l�-�[L�)��"����w��|���0�'a��;�o�?��@E��l�f�⤑�E{ͪ�J���M�^���>� ��r�E�MW�=�ǖ�F͘�_�G�Y n؁Dhc��U�BD����k��'�oL��y|#O+&��F�ZO=&��eU^&7�.S�]RQ�+����7�_]��*f@�t�\�7����"I�-�oS�&�<��5i͇T�i.s� �l��yQ��	���f�j�(�nͶ��-KR�隳����*�pw|s0=R#sA�6ݴ�hZ��E�u/��4�o֜�[m/0�{�Fw��X����A$0���	~�v}{�Li�R�F�ݫ�_D-XK8�?G,q����s?Fq�]��[�v�nƁ;�2e`w���H���S�,(�U	���I+����c{>��y��_��l�Wx嶷��y�3�U���Zx�T�Ĉ(�����@�ڒ����Tb�����U��b>*YU7\	�^���H��wˍ���վ�-���wެe6�K�v[���%4������@�&�kc$��FŒ���'7	J/�իy�A=P�Nu,��O�aGU�җ�yJ�ؿ���
���.�����]��%�e���/=�����<��>1�NV�
�0O�Gv?�Q�c���	����d�oȖU:� ٪X����V������G��rE���;���0�<!Q�0j ��T��b��@s�K��G�9�44 �$[�qkҲ��e�?k?o�gq�D$άR��������Bӵ�H5��[(�WԊ��d1�(�+�_3����%n�=��Ə�����l$ԥ9ɷ�-�o4�2��F���I5��kZ
�J�{���!V���^�?&��mPe����05��)(Q�Q�ՎU�S�,bn��݄�0�8�����=G�AK�;3��NjTM��.=��AI��á�C��;�1��B׺|_2Yߧ"1{���Iy^>�MR;��tL΂���ͳ�N� �Hn�CB����7hBƏ�I@���
^��F�aK�ZWj#����L�ڢ��3��ݮ�)c��G�8'�-M/�|�	�kZ���~j�v�㊻s �L*T`���W�UX�C��ё�q+����~�f�]2>���m�\���1�Q��J�ٲ�V���ڣv�Jkg�5r�;��!����$0��L%b��G�'���:��E5���#H���Tߔ����C���s���m�A2�z��62̠�EzvS[<>��Bp�\��u�^���߂���Ն�Ϻ�&�:�E+yD�:�~��Lv�7@KIB�"����.ec=�3ܻ������ s:�	�Ø���a:1^�Z	���aB�U��1x��:6'���$�쐫�&�)��/[bp�%8٠��jpvԽ�i;j����a�G�O����Ǟ�� �}y\<&�"Q��O�J<�"�#b'#Ն-'N�*�Vt9d6�����������A!�Lo�����~x����]`V�}f�y�xr���q��n�?��ػZ�JŻ�u��M�f�V|��UUR6v6��4����͆�fr�6-.�;P�7�~}��X���~����t�oZhz����a�,|3r��� t���&f֊[!�.AuB.:bX	��^W����N�p`�_$��$��� �ؑYW>F?u��D��������'��}�
ХX�:J�!������n�W��f�f�b��P� nf��q�6)�N#i��[CC@��J$��o�s[-��P���*.��r#�^��h�o�&nu*UY���>�W(�M��kh�B�_��*�/=���˳~+��nH�����7_>�<��v� �^P�:_�ߔ�Jf��oP�g�%�����̖FHL|~�YTʣ��0�?����=��;2=AdN��U�)kzC���h�g����6��9\*��i��LXB���z���*G2'�Hr�(�+pe�s���w%}�����y^U�Gb=W#�g��T��z��Lj�/,0!x^Z�W��Hgs��]��TJ�צ7�DI��c��þ���ՙdp_4��9h�� م߯��R;W�nBcb2d��+���w�]3S��q5�����,28��3$� z
�8�����c���x���w����q?gP��S����+R	�Gfݪ�i�ڼC���̦W7_�[���1�sH� m$�Y=��K�{�8b�6Jf%ʥ`�\K�|[f�l��ݼ�m�kF���G�Qh���5%�� �j��k���Om���˿��+��k�8�nխ�n	���䥗 |mǎgU���/W}���"�B/�˞&YkщN���٨c���[�;�K�C��9��8�12b�ߢl�^��e<���R��s�K�_KE�c�lK�����C�8W!~��L{��Q�^(�Y!1����������M3x;����v��«_`Xu�Kmm��"ŕ��
�Ɗz��7^�̌��r�_��F�]�
�Բ�(��c����eO�(ʢ	m�t3�T�%�_��"8e�3�F�F9��}U+{)��0c,6d/
�?�zp���591ױ	����<�t��ṻ��>h���т��@.f`��8A.�[��j�^��&����*�����b�IK���i�e��H�hlY�?��-���%\6�����@vHU`>MD5����Ĵ1��>`Q;s�y�����?�hP�i�����{�$.n�z�$h�S���)$�ä��7�q��p��Q] 3�gȢ;�ݥ�ŋ��C�.�\���XL|O��N�oT�7�@:�춝n������o$���Хq�<�o���Qz��,7Ws��*�7�[�y���f�:��f�Ī1ǈ���<7{P=n�];��?�P�F]��0q���,�x?�y5��=�w)�B'��#g�s�� ��nh���!�x[�4KbI_����Jn���0��d���|���P��%`ڃ���?AytT����_��U�ZȬ�*��r�ʑ���Xa\2�ƀ>����

�UT!+��j���>l�#�ˋ���B?�#a���L����h�X���$+��xE�\Sh(X�	v�)D`{R�� ����c�#�u��\�}FQ�V�-��H��R�M��{ �[W7�@�N�?�'vtZ=�B����7.���õ$M��)���/Ǳ\H�Q�Q����z�pvU�Jw�4���}��ؙz�
�X��t9�@��#@��������5�pTt.�@�^���{�S|i�:�{է�@��UX�ՠ�T��b�N@}y �N�����Vۭ��Q���ZkS���"j����'�*ż�b@+?�7p