��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0q6 ��ܥ�̬/�-��!djΌb0vѭ�%�b͝&�^�u@�]���&�ɼL�B5%�y�~k�㲲{�NH��m�=pg��F�-� �!�+����l�щSfz{���V�,�M��H��>��&���	#S'd�v74jO �b$B��,�Qj��icś��[D..��?o&q����9�B���N�o?-Pn���	�w���A�N)��g����Ik�={�ʺ��7Tc��@"��@s��r����L�"�m8�̏s�P�2= R󐢀�4��S����u9�����|j�dg}{�������ò9��e������÷�<w0*�$�-��7�7�=m��̓=��D�F�)H�w��c������G3|�B8��,J94���fv��S��ZD��av�]���� �N%�jQ-N�����.����P>�d]�3W$�r0�+,A�K�:��58}EO�#���%��k�^�w��\t"�����i�@u�u�@}����>�?�F��|����1F�y�t��2ό����0Ӡ��l��8>"�'��߂)���8�^����E��d FL�_�*ش�kqk���,$��k�}�l��n��-T���#�ht�^��C&���GZŠaL2?�D�R-ږot`�I�T��SB���<nQ4�����k i����]�0�o���bp�������(��ws(;���ʶL݂��6�K���_5����P_c}�s�a���ve��,=O���*~X�BX�aU�g�a�:�����WD�%�j['b��̇�B��{ �jd�Qx�Ɉ��)�h�ܷ�D ��8��VI�n��Q�����\(2 #{S��������|��D���M��F����^D�ǎ��k��d�HX�G񡗡"�ۇㇳ��� 	kQPBP�&=��{��T��o炕&�11�;���+���Xl4�%�$�FR�?۵�F�yݚD�C�!���ց��tԡ*.Rp�����o2�8�J�
��@5�N�bW} �F`~7M/��3��!�iҠ���wv��m�:*@谗��8�B����їj^�ݷ����#a��V(F��� �`2��LCD��
�B![��A���j"�6I�9��]hh1e>�8}�rR��A���g�&xz�H���ώl���E�7H�{�o�U�+S�h�[b�֏�����_�rA���9��W��45���
k��lsJ+����P=�~��j�� ���b_e
�1��<L�8�R���y�oID����`�?k ��f%3���V�S�o�����W�w��:�6]?�i�Ol&�s�X�ν���򤜁��v	�ʹ�JQ�q����*�F�g��{�p�����=N��B�y�"�
���-��s'�I��٩��^qȍ�@:��k���+0|�a��}��8�s��`7�QwGݧo73�>c�=�%@'n*sRwb���t�Fɫ6���g#*VhA�ʷ�"w4��%�l�}�	��a�NQP��JNX���Y��P\n��9�Km��@#}c2Y�L��?qT�b�ݽ%NS�ll�g����ܧ<�¯Ⱥvݔ��*�(i�d�K��v��͊�ۈ���LС��̂���ʆ�Of�9��T5��☇R���q�Q����è�-��IAD��l�M4'-'�jΡoV�U��]�p��m8�d�Wx)APH�/\�	��������L	g
J��r�i���-��ɾ�����AƎ,,z��tS����9���Ǫ�c�Y9�]د4�j��ѡz5p�˚N.��1Ow�v���wOk�|�nm�9�3y6�t|�A��ɹ! ����P��FFí���4�3��� #�[��K�jQ��ݣ4#�T}N���b0vB�þb�ɪ���Ů�3��PFs����/��xF����)J:R�Ww^�q���^;��*~;k�!S̯�����E�@`��hv���>�P��>JM�J�\9�fw��v��Udˮ�^����Ŵ���.��4L3��n$d���&���?A� ^џ}���$�ݔ�䏸M#I��nt�C,��m�=�I����Pyv<���"���*c�:�%��L"}��"I�L�J��s�Z��p��O��lN�N����~'�H�_5��g���#�7��?2��ʃ9o{�kH���w��J0��#�$�ɇ=�"��C-��<��{�u�/���OQm�h�w,��7��1Hwe�9ޘJ ��g�s��p%>�0b� Jճ��"�[]ڗ�"���Hw��)���m�ZG6�>y$�ڊs�_�L������Gq�44������V�̐pB�v������;0��v`M*Js�rʟ��J�L�L�U���/ j�tt�8��ԍd�ݡy��A2�f	~H��I�i�V঴������a�L��+�[��]5����0�j{� �{���OI�r�5���,�G��-k���Ϙ�-ն�n=���s��Q��T6�8�*Hb^�L]�����!��h�a�V;�R0]��㜃H -�bH��Z����2՚3u<���A�Bzs��	������_����'/m��{�Гe↸����>��2K��ꖡ��x��W�ˏ�'N�;���,�`��ƪ��Cq� �YA'-3��Qd��Qy;o��B왕��D��q�t�踍���`י�<0
E�b��\GAAܷ%�a#�ECC���L�]�C����L�F�N���Q�� �ԍȈp��#��R%s�,��fz�`W�L@{F�2�YY
UL�7Lr��-;�`9��
Mۡ�:ǐ���E�c���5����F�b�Ci"(^36R�5C ���8�Wqx���/���[�ɐ����b���^�
n$�c*��D�ly�}XA�=RF~l���SK'ڂ�Q����eAMЮT��]܅`xD�e�4u���=jJ�é�0E�9���ph��>H������\CM�Y"������$��*�� ���0�^G�R�̵b�`p����.>W�G�P�;�7$����8[�4BNsQ�)q�t�ܯ�̘$�>0�9����H5c��>iB�ïe�0u�-ī�`^(��J���FhԹ��D���x�Pф��ݮr`���/�
�5��<7�TTR9\h�s�L��bё�`���"�,@@yGHͅ P�{a�������H�R�
���!V.�w�_���'B;è�mꍛ﷫��
bMiܲ&�#�?s �1�@ih���M�����m���Mo�D�Q�f�%U�!�4�VPR��~�ڌ�D�D��e�%S�'%�$.��Q�����V��!�9�	��z�KR�����B�`�/yjl����۸��DB��4S�y�D�A8{�M/#J�Z앭�7��2�����H!Y��H��B�|��楸"5:�m
���:+XҌ\2�h1���\��א�<p^��ё�,��ECf���Y�4�����`rl�+�[I]��ò\@�XT����L��"�[ʰ����rD�a�=�\9����T.b�@���J�M�z�A�eZL�IЙႁ$�@�i�BAɔrd��3�6x�x�(���߀��+�Vˆ<z_���{�x�֖=���ug#$ծ"�f�Rܓ<����"��>��E��1$F��3�Ȱ�B�4����c�M�}�XyE�M�1�: +^U��2d�2�3S�xY[�%���p�ީN#e�ln�������N�����^"c��W�-��mLf7p�:G�D�ncM�6��0~I_u�R
s����5���x�y�7�ul��G�{�nR���#Ҿ�3)(`.�['�r��4(���ÌQ��L����*�p��+��Zw�cW�s��O�
}W�*2EsԸcky��tL���☳pD��$���u���P�xWݰ^��i'g:�@��:��j�-645�ی�5�4)�+���PPK��%����*�0�g�O6)�(-����^>�"�,��eM�2\�U1�
�:�e�f�>=�>�'as���P�k!������_e`���S@��"a�����57���$dz���^?j�Ƨk�8e��Ɇ�t��d��;�,m��סbk��9
���LJT�+��%lkC�\�y��
�Fي���BKP�آ�7�~P�H7��!��
�D�X�A�ٞ�������3ܳ;� 1lM.57Z�	ar��_����OȶJ�Q^ �j��E���e�JՔ�207e7f���d�,Lt����P���<�@O�����<.���6��NR�dM3/���Cy�`��D���0]8~�𨦡sɦ����NFx�v\��D�}��j�W�����:��H�ڋMwRk�S�#�A�)�����T�!�U(�����KIx��V�>CȊ�x��'kG���?�Q�N�~ I�Sga��Pm��Ʊ�`n�xx��_.�Af�½�@���YE|L^0Z1�c[h<1OI��s�5�A��NE9=�ڲK	�u8�ŏ�ͣ����Y���7(?�I�!N�o)��Oϩ�W��6I���+9'\j#�b�!�V�o����1�%���i\�ƛl�F�k�u�SE�Ā_��xp�#����@�
���䑾��)�o3���<���r�m10��҅���"}|h�������=���Y�m�y�)"�OF����L.��A˸$�sr!i�?��U9���9��a(5�/#��%#	(�̜ᄡ��փ������űb�'�#�܂D�[��B) H�<T�
蚞E��6"tՁ�S��ˬS� ��>��7y���/5]PF�e��I�(�a7��0�<�A���}xO#�F�{�w��Rf1?��'W�6W�,��F�i���lw+�\d��R'�4�]�Q�lx�L����T̞�U�Q1=�i3X�1�Lam[^�N�Ѫ{�0,�ON"gX��M��$D;�zN�"�iٸ���隱�;�G�Y܌$����P�~�`�7"%���
���.^R}�@��e��H#}�S�黔��f�3@�2-kԊ���v�e
:���3� ;'=�L5��;2��<��.�ޥe�@-��9B�>���4bj����wuǦ�O�j!�@�^�$=��h�@�E�oQ��������*��z���M��,w�$4��w�l#�/�,7�;C��~g����1��JG H�
�^�6��$��w��amv�-��*p+���x��ԅ)]����|�b��,[���?����ⵓ/�K �M�P�HX�A���X=���#h�Rk[�3اj���h�;E��$0/�������;�A��6FL禿�$>�C�i�����y�g�ٲHye*m�����'�	�H�0�i�+ԋ����j.V��ae����C`�1>}$b/����Ӱҗ��>h�xu�
�@t��oU�O��I��<�Nʳ��B��Ƨ�3�zIg-7(++!]�z��B!~>�类D=��1�d���44(�	�ߘA�0y�)�C��(Ye���<�Uִ�Cl�ϖG����7�Jf�ڱJ�7��=��Mԡ��_L���u��Cj�u���1��xWu�?x-��D �c6�gq�J�����d�+��w��=�f��Z��̑^MD�?���I�6�������-�=�z�}La��O�����������_�t�9��_
��
w|�N��J�e��!��UV�q��+k�ؔ%�r���1
O�d�o�˅T���%pKB�-5M�G g������v�H�>&:�#;��ڔ	)�}b�E߿�g�6]�na�a��τ�P:n_���� 殑���������\����/妠�Ά\�-԰�=!
��hT����2�(p��T��	����)
7"��D]L�p��nG0oc`�Y�r^V ��l�Ś�"Zd��Ui�PMT����)���:���7��	M�3Z4�oP��ߠѮ��R8W�cx����韦p����\򢪃�q��FCx�pg�&�>��#�ʘ�<���(n�gP����Ie�<}�*��d ���)ON����L��²��pN?&�W� Y�t�*r]*8}�!�����Zg���
y~� Ye��%XD��6O���%ڡ�9�#���_�o˖!:7��ɔ�Qۈ����:1ڭ~7NN\�/�7,�,ť!���Jd;�q.�9�@M8Z"c �4X�'S����=��#C���q0z6y��'�TݡH_�8}��,À����ȇU<!��R�5	b�L���*��V��<�	}�Hn�z�E���R|�������Ĝ�g�A��ٹ��9Ӟ�gEM�d��> #��5oY�	^�l����]'ʁ��h���,^���6����	E/�lH�-!� ��:�yAJ�6���ِaos��I��$�#�Ҟf~f��2���K�a��s�?��#]��	9B�o�S�x6����0�D^wެk�9R����_�4�lx1v�eGȞ��Od�x���Q�$Բ�D�y�8�!.t��gI�����Mg`��p��	���H�/$Ml�]8F[��Hv׺D�UT=m��eKkzt�٭6���Wf!�Zd ���q����[w@�43�G���W�v{V^p��7O(����>���D�B@zL��2a�u�D�R��y��!u���)���d���&Z�ӥ
-�-U�Ʃ�4���3y��O�ڹ�xc:e��Nz��{Z��v�J���s�Zp���hW���7_��؎�5��\�Xy.��q��v�caǦ�Q��'����i$�s�R��.y����i\2�;�
�xyO�F�!e�������~�-��u=�J�=���Ȩ�!�6�1��f;N"�B����������t-�+�M-�7iCdxw1�J�@�^�>�6�]d�����M����o^�I{��W9U4�Uq�-9��C�kgGќ����,�ޟ���Kc��������4����R���g<` @<N���,�2%�Q�󦸼�Ui�F��8��_�~j,��8��r�G�a�YLmQ�`��X�Y�k��� �c*�,[��?a9/Iaj�@�7��L��"����i�1߮���{Y��@��(
�^J8(BK�z(P�����IK���w��e�V0B<��Ibh�ܥ��+����O�GIL�\�8���q~4H����D/�o����@boݫV{ص�`Y�����z)V��Io��qٽ"����X�Gϯϥ�	����'K@s�Np�M�qyն�Sxx�}/�_Y��������3"�w
�k�ߵɞ��ٻ�2B�/##V��rq�-K/D����rt� W%jE�~YA��� 3l����F&�&�0���|`V]+��c<HNX�G�11YG���*f��i4V7#�ƍ>��;������q�PԀ��t�2�- �u�V���&ҁI�W����2gBm|x|�G���\�}�Q�����c⩠��Sx	㻱�$����m=�8���\|�v,r����{���z�8;X���N̋Q+i��V�OU[O��Ю'L��M�	�Y=)�%��<[$�`��Uk�PgU}�£�Vmi�J�ڒ�8��di�d��~8��Ƶ2�Ɓ�bM��}�<9�Ǣ�"�`��~�"�����{3�?{�s�?����E{�CVyN�a��r3%ױ�s��Y�k��]��q;l�U�Ɛ!��C��"4I��@Y�Ho��C�|����LP&�^{�!�,p�ڬI�����P�vnϴm�I�b�iN4�?�i�����J��*����ZI���*	����uDΟ2*lpH8�Q=�^;{y�ѵ���d�\���U7�2T�4��