��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`pc���e6��'��) \�t�"27g�#7�bZ=W�JN�W�J"��̳��O+�vi��ᓎ��z��6�yU�g�����r�����ē#� h1}�W���n7��x)�r�ez�Q��B*nn�s�a&7���b��v!����|�qp��Q=�� $F1/�}������x���u���Xtp'&�Մ�ԫ�^^�E�er�D^�E,��:��	����yf�0��=��-�&I�x����K�?�t���sh[��1)1�>Pl)f�5�9�F,�t���dM�=<*��O��G�7^C�7�{&#F?��gGQk�m@�.�s+�)/�A����ި�z�P0j
��I?Gi�k���n�mߚý'
��]����ʢ��b�L\���8��MaBl��a�Z�Br�禣Z��OR�HO���V�z6�U>��]��:*'�#T��O^�hz5�1l�X�>G�035c
��h�s��|�QE^ӓ�G5��GoiJ�!�'ztZ��0��*0�������ta������7%��e�i/MsZ�a#�p��wV�e8vB�۷[�d#�"�Q���
�>ά��W� oK���e�v>p|p���6 !����=� �C����3����;.�݌.��
ShϽ�������X���wآ�8�]d���|߫���=z�}n��=H�u��i��8�K6?񹫎�y�ݘ�T�N�'`y�\G}�(�!���{\*4��ep�?������-I)?LI6���s��\h��g�դ��c��Es͡ڪ�=�ÙEJ#�ҁb��5�^�zY�a�h=o8��g� Un�+��?���3��O"�/񏲖ђ� $e���9��Ӟy�����M�Ä�p��2��﹁�%�t���)���NBҥ��:�eUX}n]�q頥�j��!�-�}�ݟ/;X�c�agk�D�c��)�À��'�)���Qr�%��+��V�XS�KUf}9�:ݘj��{x߇��@�,$���?��I�G��fn2yУ}�0�2�Uz�]`t��/ �ADF�}�ukVw�'F����7�����J�f6fe`�\����.u*~ӎx��ByW�d�5�4�m�M�9uU�8왧z�ༀEA�iU,�P��b�$U*s9ѱl��/*�H#<���3����-�I1]eJ@��
{���f3%j�z�J*3pa�Q\��oY�$�����?�C��;��7k���v�pF�s~%P��>��X�8��4�����*��F��p�	}I��bA@Hk�~
i��/�?�WO��i\�����k+�k.�@x�ʾ)��9�ı 9~h\����&@j�
 ,�Ƶ���QK�'Ud-$��b5J�	�(&�'���nT;D��d��s��+v|��rCˣd~�w�KK�����pf�	P���w��Z���0N�:HG,7������h�-s�d�l:(��ˎ�8?XA���\!I�8�V�Dr.iv9ȤF�T�x�J0��;���*�p���� �3\�H�@{��� ̛Fv��ͯ�χ�׭V�4[��N'{���gr��w(�ˍ��|-�A!za�>F���u�R� ��+�4�Y3I�R�=oI���0��_���I�;�,�A6[h��Ԏ�<�T��f>%*�sbaN^z��?�`����d�2X֭���(k�p�J\�����<5����r�=�xCW''B.J0��_[�ʉ �j�Ȅ�+�-Y�e[7om�Gr�����!�,�3�
�o<C�m�,�0_����b�#mS��Z���#���*����KvxQ #}��D�*f&��cDB'yMt�k�ȋ#��އ�D����Yh�imG�y�<�
^]A6�j�����"1-ĂؑVޔo �6V���ks�e@��';!ؚ������J���	�R�5_�^�o��o?�?�!U�p�ܑ�߸4��yƋ���䯪�é�[���Q��#񻧬�h��F����\�J�yd���pЂT���|���oQ*�Y�KӪ�K�5뾺�ҫ�4\���Pe�^��Gv���֮�}�i�B;Y4�m��q�y�=~�.��9�C𥟀�.6Hb7vL�ª_��^�6c|c��9��H]�D��U%R)]Nm����rƎz���>*��Wa��9!O���m�
�y�� ��S�o��v��d��G)���'���M��B�.�� �cX��A��ir�_�\Js1� ��iP_b��d8�V�`�3��a�}&8|�l��c$�a��Fo[�� lCyN��=��Gh�lm�{l��jV�{MW�H��b�� B�u~; *��3���f%��E�p�q����*m�
�oC��{�����Oʰg Lyl�+��-���TO�R7U���
c�,cW�a�v=FT������%j`��,ht��aؖ���¢�p�{Ȋ�8�T����Ht>%�x���,���Au����'5A�Ǻo�R�RMH�͜�$oQ�1�m���Ɋ��W��?9.,�R��?�H�`�Z��ڙ`Ԏ��:=k�K��OH膼��lL��k��?,�Z���MM�b�B60$�E�-�
�֯���`��1g�h�ѯjw\'��,M!:5LUX����j��I���2>�د%�&��+�����o?譌Fޜdܹ��C����h�]
�	Mk���i��p_���Q򍥃�c���h�����s���o�kQ�O�G��<�Оn�ޱ@�
d��|yH�=F���~v�c���x�kֻPZ��2=� �A�1xa�9HcL1�.ރ�c�j!����ry��qNv�5ϸ��d6�<ؔ�Zu��
ݼ��G�+��N���@7�p�~���j�$j^x}|�2���p�m��<��G�{���4�@RW��+����U&��=�!z;�X���&ߍv�GW֒3������h�6�K:2�����������o���"@�~Y��h�/Bo�����v�wQ���u)u��oi�$NDz9o���/�9�m���v*h='�#�7�����m��T�3n!�Ҥ�j�k
G�����t�cř��n�ש�>)�Q`���7!�uV
���+6甄�O�6rQ�s�K�����Y9p�Q��Q]t����	�E���9��R��S1��`�j�[�f�3��#h�3���=%�����0�geP"j�׾�=���Kr����O��;?����%�>K��J���`�/DL��E�&��}/[S���n|��f��C7��N����V�OєMJ&��A)ੁ�R��~,1���lC	Ic�r�\���ӗms�����g]���C,��W�(F�+�m؎9�k���Ms�m)��M"�hA�,�C^m�������5����?�F��<�a�N?6�ai�)v�u�dT�~]g!7�q��?�ll0j[P>��E��F�~�S���	.�*��Eऱ���4Jmd͋�Y#���;�0�v 8w�x��q�s@V-�bL���]�"��,����Q���Ar4���*�"ɞP�Ȟ�b�/lX�(�Y?�3֎�yuu3���jO�	��8�����Z�d3ߥj3	�|����wD���#�>�yY�*���7�J�H�'��kH3E��w�ĥ�#0,�R��g��hD�Al�X�3V��Q��QN�;+����,�>!L�?ψE�4�>ט�	D�N��Zꂛ�ffY��b�V8_��Fb��qS2Zr���ō� �x�82��;�	b�K����JV�iC��͞j��QA��o���>?Q��R+z"�5�H��c��Z=z�S��)��m���oXew�dݝ�=�]g���O��r���S�ҊC��Kj�S�����ʆ5��Q�¾��@�Jh�u
P,(�_��Xq4<!���yM^����c����I?@�����Z12`�9��� ��CvaR|�W~nxvyJ� !�xM�V-W�~�Ӭ2�o߄Op[N�<|�5y�1���D�P��&J�(�L����Г��`�(����Y�F@J���w/�7�t��ƿA��4M�:A �g��=dWp<�'��������N�1|Z�q���ϟES��ާ�>�6��&�p[ &ň۔�x���6SX�P�!��.�e![֔��Ԭ��qĚY���C����~��Q�(����խ�LqKhp&�^��9�n�ic�Dlo��6����!��{^�m��˚���*P�g��]ks��Z�tϧ."� �z���'[�I�w�!EM~����Z���� ����j�7���Z�hM�P�w{��0'y9�m��Y}�E��]k�!X����-#���>rŔ}4c޽<"�=�J����[x]�|�����-������\ +��B+���:�q�[�*�L\<��8��Ves���f_��GA�x���|%�e*Y�цLy�Q��wL��(�B��P~WO0,N�#aa�:�e��غ���A�[eGb+CN��}�vwf�y�l��39�ф�iu�Vv,�#_ި�K1I7]>��/O0e�AU(��RB`-��{I��9jfe�o<_�Ԇp�N��He)f�{��q��� ~J2�uj�@Q���)Cϊ�؉W��#�ͧ�?'QQrr"4e[q��>�>m�ZG��&���}2���'�C��wfB��6�}�HϚ�۠��	���#n���>e��0���.2�vֈ*�\��m�x�@�Tܻ�h:�a�[������/�/f��� �S���]7w��:����� ��AT��?Dcp<P�nh��H7t�{kT�;���*��(�X��/�}g2*)�����A�(�wK}n��ζHw�4]�B^doԥ�a=�o���(i���>�}5͑&G7�D�r�]�*����ٸȡ\��ʶ˽H:�=h��q�zY����@�wޥ-���
�z�<Т�'ѯ�����Y.)�L|%]Z��r�ρd�J���Ue�m�G�EH�6g�?g�����8=�H-� ����/��(h�m*L�r��ݭ��Lw�&V�	MfHH�ª�l9�w�"ZkK��.c�h�F;�d�|s[�C�h���g�z����=���.%��yy�P����@Xg<D�����}?�:�IR��6.�թ�6�z�,�m�OB��J�s�V��f�����.�~@�A���yb0sl\w���f�a�j�]��&��[? �Bfy0��v���)<|��\!�{C�@)yV�1�DL���.QP����[�SMx��f��]_P�[��'�Q3�Ik����ԯG�����'z�k �j��N/w� [IxF�3�ꔴ���W"��eW S�K+�-��.�HZK��b�u&�Q�}��G��3�.3��l�A�U8	I��	��nrD��҇�:����|�V��������uWr5)P���
'��c�S��˩m�{�a���ühI&�ni�>b|?�H�$��~�s�}��̍�=Z��f�L"d�҉7?~�5��-�ӿ˲�����J0ʣ.�(0���&�
`Px�[,9���X.��r�3��Sa�B?�y{�%M&��F�u-wY�s m̟��p��J���>d�PL�:��=�^U�x���F����P�Mxt��(B��܋}��q﹥� �ם�ƭ�c,����D��XsR8}�߻P���"�nT�Нf)��4=4V?�	3�@�;�a��}y�w�͹`�f+�h�t��5��H
�G��.�D�.A���x��x�|��]�8շj�j�>Z�N(Si���	��Wl�,�/�����D�����b��ア�M�b�%c�����yrm�ĸ9I�g��K������G%�4�ٯ�WS	��X�c8�$�ԭ����.��.^w`�D)�����H���� O��
�L:�`@�x��K�_Sp�ȵ!��mmh�J�5�WQ��,@�q�ߞŏ���"�����[�iF����t=�?̩/Y�}������p;澤rȈ�; \Ӈ��*H'> ���֮�m}��[�I�sI��t+�w�꿫�p�� Z��8�\�ܪ*�V�\׽m �x��\y�On@%��-J���,��� �����=��� ���*<��}Ђ�o�~���F�ٗ�A$Ge����R��|��+�<��q�рE*��dÖx��8Ҹx�4r��!v�T��E�<7B���sDO�� �0٥���R�
'�&�k�'�v�ba�*���\
ɬ�
zyEذ=|75&V��l3���u'� Ԯ��\&9S	h� m����\$a1�z
S <V\�'�����9j]�5f�r���H��y$f���'���~}��?;�7v��� !SR��Д��Z6���ڶ\`[C�
�\�v�r,�e#Ia��X��5��}�-�QڍUqK�rq��
]�3 �_a��ecb�ҝ����Y���c�=|;^#M�.����$jBԜ	���:횊%�Ͽ�T��_�������I9�%�͢Ϫ xy�cka4n��a��K���&Qs,-R`�Ϙ���k
�+w�Y��H� s�DMT���a_3��af�jL�La��aI|�J�O����0i�뵅{y�����A�r�!�~�ݛ����=>��Z�_l�&�Y^����d�t`� _� Ahz/n�ܿ:Bp���7�n�*If���O$��>㊄[�G��pT�V@����n����ط��A���C��|Y� �ٓ���1_��T�k>�2���P����P#�Tp�r�������*��QO�]K�Bl�%[rfƈ�FǷh�꿹A)�x��Va����[��16��B�@��\��6/��,�?��AI$�!�b���h+T��b�~P|�U�<,�e��C�:�q
O ����(��1��`���wl�����g������ 0�Z�(pW���Ih`��KA��W�H���rS�z%��	�q�u���)|%FwN�6�~3 2/t0*n��F�����Q���<Jb?9eW�N$b�J�D�����������������+��&q5Ru�7*���Np �XYZF���?>��D�Oavgn�WU��9
U)���k�w:@���@,*B	��#c��Q	��ƽ�,�.�u��Pn
�L>��ޫ���Z����)����n�-�zi�$�X:�*���e�%�A��$���J�d�x���m�h���o_Dq+O���Z�������H���#h�?�Z� .0A�n�Υ��S��.�`��7�<�VV��:��|���5�++5��⡇3�E�~A�����dV�P���̈́'�����*��Z_ћ�^f噎G�����)}Ww�~^c�bd�����=V|\eLb5��z�f�OZ�b���eQU�=+��&Y"-����jJ�n���̔y��ca��x_"۽��� 6�p��OR��V���-:\��k�O�Ov^"��6:X��;�b6��+��MT���͐��fbw�7Zy@�׵�\Ԇ���gV�e��\?Y�2�ٳ���1%�X�4�^s�wj���ylRڤG��ʟ*������bmQN��{՝�O���8UTgC�c#u �$��?�,�o�����.��iښ��ڲ@�V;�|�Hܫ�Y8����)�2��ǆ���[�3A��?MVVZ9�m�!C�P����Y��:�|�'x��9)פD��@��]P�v��jؗ޼�K�N�iRShܐ|�z,κ1��t�!�b����r�y���4&�O�D;�ݓe���6;�>�5��]�����-e��-�k��~e���~`�C������ػ�H���Dk�;�ٮ�2�8p�O���S��/V��C��wZ�қS_\y-�q�`
LJ�����O������$�N?�NH/�|�[9~���6\E��v�PY�,)�
b<�[���U,�����վ���2IpD�`�:��׵�9�k��]ӺH��:͖ ���+i�;�5	�:�p�A�'=ڬV6XMœf㷽��	��̖��b����S_y�-3�d�{إ|+rs-�)�j�50������p�Mn�3��W�	���\�H�dX�QPt�;�v�f��z����y���$�%�`�>3�:8��ph�6Td��%�9�a|=�ԣ�t��^�3��jL�Vd���P)�>�Oj-�Һ�1��\�2)���L�{O���F���uJp~%�`1aq+��Gؐ��+�I1vP�
���3�䄵�����GW�z���s41�E��o���v�B�46� �9�D�˟�U�-G:P�|��'���a9Gɱ�R1�i�HOD�|�Ysz��f񸟙a,$�ש����k_�!�E������@B9,�e��Ŝ�o�Ơ ��!d��6P�!y;,P�e���³�t�m�����&��0Ȳ!����d)x���Ft�H���2ڀX��׸<���w�0�+ Ƕ�{����~��q����u�'FZc銘��s���d��}�� �Q��SN*�{UuHr�>�9K�c�'R�z�}���[|u�p�.0���4�Yw���������<�73�q�E� ��"I$@�AD[�"��Ӗ���/�xIzS�(E^�`�7~��Zh���E���F�8gL�8�.�W�Ý-��:����u���^/��x�4�p�ő��Q!�B�r���>G��`Tv����v��Z�n"Ne"^�\��ަ�Klx}���D@%�φ2���������#<8��<7��Z*���@��!n'���*j͛��g%���\�m?A��z�C:��j;4ܱ���^��.N7&#�">F~)�ؑHW,bC�{x��*5�d�y���.y{)U?�>m�{Ry���{��������gǀ���m����)'�TI�!�T�J%�"����"99��o�+�!K��I��0��;�{�t��y��y�]V�+��������
����S�+	�Q�6*��y��2��xZ�$�Zq�/h'�/��Յď��X����W�K<7�2`��z�y�CPi�^	��+�^'bAjŏ�GF��,���=Ra��~D�{LVU�oiQ:��å6����.��Xщo	tߌ��0�nQC�,�p�r�_�zN�S�Az΍L% k�Y�/�b88�N���N����P5�&���a\t"�#C,�ǦGf�� ]1����Z'��t���w�Oh�NQ��y�.�bn(�u�p;?u�?�ze��EU0�ܲע��݊����xN��ML�%T�n6��R�1�o�uȝ��(e`�CW=����x��W�/"xR��MH��J�7� �+�WQ9����Х]F�U�+a�`�-bwc��(/Ȣ [�X��Tȗ��ۧg��Z }:�44{@F�K:0F(�*P��yz^rfw�&�Ϥa%mR�o�5U��8�Ѷ��ק#�R
%�_�͙��A⮈�E�R8��Us:��¸@����97�)��Eت#�G�a���\I
���hv@�����"��q�o@�p��u�6��qE� 1�𢻄��F4��U7�l���OWI���4��㰵Ip`��v��r}u�&��)4��)%�"��@��< ���4��3�A�sM}���Kz�����4��I�ӹn�SH��;_R��K�����lR������X�K7ؑ��6�}�M���%/	S6����Z£�Pt���8x-��<��|�;�
O����q�w)й����$s;6+�������vzZE��	w��G"��l�������uI�ai�X��0�� �� ��k���'Bp�bAk����!�`ǯ�KO�����ӎ	�b05�$��l��z3.x�Gs~}���!���GϬ,:>OR Np��n@3���CX����+��Y9Eaq$�-9��N�~{�ǐ%�4��>�k��2�C'�:ᨁH.�6�_9�?����䯞�ʦq&olu�g�s�dEj�p�)m�Ƴi5������M���y")����h�G���
v��ޔ/�&�s�.9=����.51UP�;?�e��\QE4^䀜�6�AW�|����XK\劆L��8R�L/�ϰ�Ȏ��%!i��g�l�.��S�\~����4���:nr秤	B��&�͛j���i������G�q�=���0����L��&�d���/�8���]Z����~
��eC��u��,�W���.����Yݤď���SI�T����҆;���x����2f�#��Ki'���Hc)ݗ�QF�ct91a4P����>hez�=!ƾ�kY��u�����qb!�����XE�-�a͑��c��2�\��G��˲Nj3Z�M]���+�(9�N:�j��磃�Vm#R+a�wҲ^����l�;1�Ñ� EB�8�X)�P�76L����س�2Y�z�����5����"T���}T�lH�X� �������4_š!���������ǒ���'��!N'�X��ߴ-��*f)�&�6��<Xw��̜li�6�/�¯��G9���%�t�έ���8�|E��֌��I�:a��z��x��)��o��pe�Vf��5���ZS�V��5�e�Kϸ���*�_u�
�ȡ#���������G뗴��Y*��~��`�g�!�H���֕�t�͏���C��?�I��Nf�W
J��ý�9�i��J5��U��"�9�1�=�J�Q�e���-C�E>�� �	��9��&Ct�V� �먚ׅ�=���>�H�)��.ܴH<���_��f��g8��o\q(Ъ 5p�Y�҉�q;l#����EVx�7�-�/l(�y�ы>&QR��
�������Β�4�����1��
�]x����}�;�DyK+���D')o��`�c/,�x|Зu'�#qp)$]�6b� �Ƽ,^��쪮F�Hgjc&f~�le�T�d���i�e��п50������@��Dw��0���l��\"���8P>Q}�[�8�eSP�"v	4��f��1��7-���{��x$��-��g�	�夼� !V�������e��[J5{��Hh2��T?)]�j�����L����oH!�E>���D��qAh��>��[2��`���C���|��|�!Z�#�"KL��T���&� ���j+��������s㡌�`^"�#x
�j �;�x���s��L6�?h�.�	�7�Bo:(:ZN#��I�c`���>z�.�T��a��f�a�{�*_�� 	]j������Ha�_)#i �ۉo5Ha�~�F&h�X\��rH���go�0Z���K�����<S-$�������v�ox��"E�F��
ֳppy�s=iy�m�0�F�::�%�Bɫٶo��L���;���eS���r{0t��e'[�ˀr%"��~����iCx�4L�Nd!6�@10)t�r���F"\W7�}�_fb<��>��μ�H�oKE�9���;�nKy�~Bv�8���#��
N牻?֨����D�r�ך05+���8�VН��'�j�Un�[�l����XɃK�(�k)2��S�I���+M��H������ ����c�I����q4lh��ӣ�?��c���6"{�k\���JMR�_�<��2?�B46g�Y#�uJ�����:r]�����i��jꜪ�fmUF��O�.j��mΊo+r��4W��	��-�-��N��grA�"lh�(�E��=�r���o�n�~�����\;z �P%Ww8�U$�r&����y�5ᴭ_�F~}�B;�F�FE>a�Q5�*�Lm���(~^���j�^)��ެ��ף�E��'S�����[A��ޟO�H�f��	>�Sgͬ�?(�hTdܔ6{�l;�v;�nb��$��+��VdZ�+9�,.��ם�J����X�y��j�Õ�"��!Ƌ�Η�s��(B(� &5X�����$���N�Fb7ܚfz�}���^�$$�?~�B:^[U�/� HF��@g��)���Y�ɤ�w��(�"?�d��:|�6<K Rg�,�͸��>紩9{+i������MX��Τ:p�}��4�Q�P���Ln���	�^�t�)���1F��,5K�[wđA?z���̂sW �"u/%ۭ#Q����Il�Fx'6�(�@��~��BF�҂���0�嫷w������!�����H:��b#mD�3���M��m�u���S_?$��l��<$[�Xp���>2^����Ya.q�cN����?g�=��a���	�.����'�Bk�šA^Q2(��ݏ�P���{K�� ��o�s޴�/uGh��z�������}�H@�ɗ=�=�y��ŕ#��e��J���aH�pR��I��sc�&��$էQ���L�śVP����}1&g�����Lb��鱠�#��f�43��!��Y��/�@�y��ua֕V��X���g�*0��{�l���n,�=-��=�Ѿ+���r�@$MI��}�_m .�6�K�)1�`q��|�3N4l�(��v���\��Ş��(�ǽ���I��{��8�H���R�b�b ����Lnf���x�
olYi�GٴD/�ߨK�k��C[&��H?ex�xFgO˱����Wķ���)c�G�}3{u��4ߒ]�ש�6)%�f+ �	n�	�㉚��o��v��b �6%�m�����`�\)4�*��W�2�4R��:-0,@�0dMoI�9!X�Z����S-�@vJGjrݮ�̪G���鶃+���������֣	b�0�����s�'UoХ������A$�oQ��5��+��e3}����|�x����.��G<�Wu�T�)�t=�/��D��=�@W|X<ts:6�`wfQƭ<a�@1�{�i�,���9��#�I
��0���B9^,9ټ��`���@����jߎ����G]<�/1��l�TEx��A����n������G���.�du�(	Nń�hj�[���l��+IF�������&�4iQ�_vŘz!x{]C�#�8�m�����n6L:��_�A���1��� ���G���f��#�64$,��)'`��8-�q]����Q4��-e� G�T����#P_�a���U���i&ڞ� G�f)˝�q֥�i-J���sݑ�/m��$´?7�<A�@`-1fرN��,�o*vz�=[��ޔ.�"�P°�zjB$�ޮ���j5N��H�o嶡�)������k>�n�(0���M�~��.(��z�G���d���D���;Z��v���Ɠ�<�M uA-� I����(��wL����6E�k����8?�m�:��t��躤v�q+�P��"�NN����GqG`��MR���O'
����ɮהݶ��=E�3G�A���g(< '{��ܪ�K���dS�|��zcwP�����9��}�,��G{���:k"e7Irb�\�cOC�o���F��.Az��Hc�t*��Cc�L��q>��P�]�֭�ZW��8E��|ȩ�3�J|ȭw5���S�ř�
\��a��\��W��vί�t��JI��W����M�J����tN�dX-u��<��lW��16�[�h�{�XK���Z�%��Z�W�Қ=/�?������Ԫ{�0��z��v����=�v��	�bw!�_(���l��cw�Y��Tr�ެ�+�
��;�Q�+�z�i�g(v���Y�)'�r���h����5skW7gE[z�D���'��x��'�X��� ���]�x<8���!��b=�O���l 7_��,ٚ�|;����	�O���îj�U�q�3���l2����u/�8���7��L��j�:9T�	�g/y=Wg�n���
	�3N�l�k�;���e\m�~����q2]X��UQ
z;������x��W��h�|�Y�y�nS�\����Y�h7."�#�*���i�S���f��ߦs�/i8�4�����:����*�^i��ڛ�v˄�;��T�* Z �Hr�9���{�NS�(#��*�Ҏ�%f�n�i]�����twR�G;�+
�f��x�I9}�&�Y"���0�b=m�̻)��>����eެY�0���T���4J3pƏD��-3~-Xxp`�J������/�A��
.`�ɢ�ݽ���8�,~K��cT���Sٵ�@+f�W�M�Y�l������У�j�H��e���\�{�,�(�B��/�'�á�<(N�ܘ�M,��4B��`�P3+��c�.LA�.�P��rVl�y�O�8����pz`o�u%�}���<���h_��-G�]�.m$�Fz�r1�k����P-�
�i�����S1-��ռ�ǱnG�-7{�)��A���>j�^8<���U�?p&_5�r��A7�|B��jٹ��	�w�qWBaʓ�uGf�io�{Nr�X��<A3��Xs��ԃ������[ x�7^r[2\�P׆Z��,�B��4�n�~u�����_���Ɵ���b��ߧ�M���M�j,�|���pUpc&�`#j�J�&��D/FT={9��}/]��/��+=��Mp���z�����Z��]�|�W�?�ȼ c�<9���
*12��W��aL.�1�1��e�>�� ,��,�a*g"46���u�]hHJ�VC�F���փ��9_�lY0B��=�f�0���.pK� �n��]��-��O��J �׏�L^6���s�X>�e�y5|��X��/j��W�U�Ē�(�_�����pH��Ofu��qt��5�
���d	��ۗ�D��ZPvt���[$�Et��C��)n�	p4�TPL,�����ΛHv��B��;&�!3�P�z�
����Cb,��B�"�8��`�wރ�y��-"1Sց�j-cc2��di�;�Ϟ��x+F��f�\��zh��<�W"wF��ٙ����=�XC�x��Ev�?�E�u��0���G�n��LsO�ؾ�x���Y6X(���_��Xվ�Lv�>�O5�BCq��r���6M�Q5,���� .�d���b��u f��?}F��[�>�3�י�T�|�DvOU�s��r�u�����A:�ޜ�׍���3�ہ���k���P�q\�sf�J$�+BITq�U,�/�6���&s����W)Y��Y��q$�%w�;��y0�>���U��`�C�{��(A��E� 2o�'Wd���`�xv�Q�_�u�M;�ұ:Q�h9�ꅃ��dڹ��h�z9:��va���M*ޣ�l���gS-�53C���W���Gt��\�9��Q�M�-8�.��(����nq�jڿ}`o\�4�C��q��I�|;��ƋIQB��W�T�ړ/��Mw�SX�\j��䠙�X�v�+^'=i���Z>����>$��u=����#��.����`�^o�Ige?N��ʓ$uD�JQ�h�**5�}yE�Ŷ���S<,�g�H�؇A�Gt>�����>L-� 9����N��Hݹ%�Q�*���	��D�>��!�{]�?��׺fס��vٷ2��B:.p�Oxi�l�T�R�Ӊe�=�:OI�T�����#3���Z�S���2�s�b�ϸ`1}���z�K�@N坥r�Xn�{˻��-�2l`6�7��I��V�<c��(��%����#B/�6�ޖe��o�*�#�ܷ2$Cx#�y�af}T�d�jQ���z�S��HR(�|o�0�]��z/���!��V��fAB	]!a��d, �Ж�+�BA���T�/���<��-���f/�-u;̞�إT��'���Ը��U��9����E��Dh��$P���}�|��u���s��8�Py�u���(�H�I�+3L�HͰ��������?�Fm��x	Q���A͙�DU����]L��NKH��@)_�.�U����_�`I��������P�}"�T��[��&�p4)DJS���G���XV�=*�)b�	���3���!W=���64o���X��$繘�������U�2|x��t��_mP�3t)2w���t���	�����CH��:����D�jDh��zHi��*=OM���`����9x��T�
���w�S�O4�G�c����ˎ��(|�E c^ޜ���vM@�F��\=��Q_C���8�W�d��xz��ͮ*�D��dlqY�م+ ���H���܈e����C�O`�Lq����؝=e���c�Rq>	U����:ŏ{w�;�p�ý4S2�����k���0aw>>��nL���;�4�6�(T�P�L�>B��ݙ�\t'm���Z�1��B�W#l{	��m̎��N
-9���Z�����`�C��W `�u���(ON��j�*����մ#cs\��oM���6d�^�|y~�����d�I.Q@�kC�K�5�BZ�̏0B�ɡ�T�_0�EH��%p��=��[�OAQ1������U�V?�U*o�H� ���F�������W-�hp�٘箯��?��Q� ��UtO��r��.i����Qg[�YĠ�[�-��03.��g��#2o�,�3�~�ۨ�	�i�?�W|;
yvV�s�ܑ����P{��fA��9˭����5�W�
6Zk�=�y����@�G�>h�Z�����c@�ˍZ�6���~��5Q��
�x�u/V[@�͇��n[Q����9�݌�Ի�O�)����Eٌ�X ��[5��]f��F>�����B� &|��D��ð�P$�l�h��	��*]N�a��!ؖ� a�7 �y� �H�-��wV��K%�}��ӑ��)5����+�t �L�A�&����Wa0�Cǋ�F�ٴ+�K�q�����.��Ý��";���ml�WA��t���`��J�MY��7���//C�ÝH!���\s�`��^-zH�v�[#3w�Χ"%q6N�;�� 8)��@� �g�\hxsf�����Y���R�������.�>�Y_�|G�G6�t5���0֛υ
ཀྵ��I��9BB'g��Tƨ��q�~1���ă�7x��[R�5�*����Ur����Q��h��qM��I#�i`�$�)�5 ��~�L��&Q�J�2��nqJᯁ�D2mZb�����k��7�8�����x=����HSy$7ǭRWI}�X�� �
.܆�D��ޟ�$��Q���G���k�8&k�_�Q��-U��{Dg?n����E3"�Bz�
:%ti,(b|QG [��xoB���H�7)Es�z���pVj�������]R�L!J�|�����M�.�{�Z�k�:8��A
�,b�@H<��=�p�ti$4@ɨ4�]�ibɡ=�Cg�o��D�BK���4 �\��~NXN�#����4��U!��i\�W�E>�{�S76|��>��5"c�_t�ٲb����� :�&*��8*�.��~ ^���F�u%;ópƂ�|��ğ��n�3WJ�݋�(TB���Ui��Gw���%J���t5� e�e2%k���cꩈ�BOqhF)�3��OD�E��5la^9n���`�[��W+ك|�dcM�m��ojʩ۳�����j�l��P���P��pE #7[���W��ae'�����r,bl��}s�Q\�<勮$���� ��8���ib��h���fR2��Uqq��Ii����v���TZ.0�y4��Ϝ��㫟�5hӷ�["�Ձ���P2����Ru$����ݜ
B�F�8���R�gIb����k+]��hߓ&�����5�-l5��N�*��Ж� �y/��8:$���)=z��Q�{�q����D�2Ϩ!�����/��Y��$k5�h�8̙� ��}ʀ2��'�w�k�zF���7=N�7�ێQ��0�
�=���CJK�fv>��Y��b�/Y����P���օ�����1���� ��엟n�j��AA>\
?��zB����؃E�i"S�
h�e��0r\w���*6̺��X?ռi�2}�A���t�>�M��%�l���r�� 	����`�S��^��	k��[|v�U�����k��.O?Hthp`�>�W	N�5�����v�Ugs��.�����b��>� ~J��I����ա�l�	r!���R(�s�gwW*���t��F����i+�a�c���Ѫj��dz�j_D�x��-��T79�(<1�c���!��@�R�?�=�W�|�cCu�s>x����p��C�U`2nlhٶc�/ 1#[����.2�"P66��=��K/>5T%V���=�O,cڝ1�ձ�5�\o�_zIfo��V9!��
D{C��V�8�2�<EP1�^S�t!�N/6���<1�oy>-���8���	�!5�@m�5)il0/�(�$���z�3�S����$���I�
W���[y�ǻl�{]�N�>�_O�,ht��o*J�!���-�[��Դ-�}%�T/W#������2�LP�TNZ���6@�}1S脗��{1�R�:J/Q��=eK61����~ؗ4����k�1<�~�1�$�p�6��z7�X������;����x�q��h&c0���9��;�TX���c�E��I�E!��&xB���	G'W�d}�k}]M�B��.�������D�_���J�]����p�<
0ĕ_�v�H�;V��k�գ���V�;��W�Ŭ��`+���=���_fn���>�π��	�
܂��#�$�E �s��{�׾��l |S�'��D�c
 �<�KB�G<�,:��?ld���� \4Y�c&+��p�"���χu���L�t���#����mR!� ��fp{����h��&:�*�������r���tQ�_��џ�iiY�.�SʔZ��n%�~~G�W?��[Bזt��>�RX�����}�����UE�mOq@�I�86���@� [�o�$f�|Hwfl
�.1�n�H�,�ͣ�) ���1�͜i�Y��"� �].i)��������*w>|��#������"�6;��7�����b�.��s+fq�����.�~d��ē&���e�X�%�{��snS�QQZ�:���I��\�Q��8�����}��8wo
a�?8��Xl�k��N�p	���~���a�U��]%7l��#�ѩ�p�q��ؑN�[[�U(�_E«V�n�[*k�CF�]��[%�=���RV��d����a�"��nwJם�E�� t�H)"��#1�)�(��mr���������uD�$j���F}�|�\��w�i�"4LYB%~�J��ف�ņf:� Ck.����j�9<����[���d�` ��P�E�! ���fq�'�`-�4=w"�-�w�[r+&�糲3H�h���'��{�H�i�������� �!c��"mY�Ѻ�JgO=7��ͧ�� ��\m�� x�0UE��׆O?�:�:SA���W�[d�t�[)"vW��kU(�e�:�^x|١ �������{w�9W1SM�Aw�S9�|6rYgS��0
�?�@�q���ʴ��'� �����d�زG�����Ȧ������	�{'Rİ`��@��}�%Ga=W7LgD�	7�H�"ຕ�x�n��(�:k����5b���cG��Ҟ$����	]S&B1�d帥aOB��\����<��(����zf��䫄#�3zt�2Bb��^H������"���Q�S޲��\�:;�9<�,������+hh`�&�p�I�\����6CYZκs=Nu6zT�� )��*x��=~zR��c��K9R�Z:�\��~U�����X��];����${���8_���V��I��GS�捨�!J4{3s~���
�t� 2G�������[:���nc��s�y�r��A!����F��<)�*F�����p*�G����xU���U���v�^/<�1uźF��ۺ�u�['���n���?&/Y"���W�^�[��I����e#�Ҹ�����mt��5D��<}�vl��^_p���=s_�Rhl2~\���c`��}I>H	�v��;���1����
��M��[ҠkF�{՛�9����=�я�u�Ϣ(-*��X�:A딁���~ �����] �oRӇw��w[��a�|�\�Xm鬾��,]�F�9�0�-F얠��r271�{�����a�f�\|����^�<K@�!q6'�vT�ߛ>2�aQ4r�ϥM�a�4Bz���H���N��a�O��I@q�R�s�5׮����J�oE���DCIA����X�y���jǶ����*�}M_���s� �( A^����7/B�w��q5~ӈ�c�X�'�\͐�C��lu��~�6oc�~�&��=%di��TW�T6 �>�(����E��K���M���R,/�5:�� ����\�Vr2��%֕y�N�5���vuK;�A̈́�Շv�< Ψ)�!M����V�Qe������X͎'�#V&,3��������܎Mn5@+��f�3}F%G}`�K���%H\_{�I��V�������Hg�@UΆ`�!I�#\�u!i�۴1G �g����a+{�:W�QI�V��T.��������θ�=�%Z���	��؅8gSfǭ�K��!��������&O�Յ|w��I'P�rG����J�,��W�"#�ۈ���Ik �
������~:L>ù`l�yx:�>Fw\Ld�d��3��L��-v��u�;�mkO8�����s�ː����o��P�VS�6�����)X!�DI�ָD�5�ρq85M
�,�F߬��#0eJ���ā{�9nŌl6�:f1��)�)-M���
/�����d-LT��K>9ߖsh��FvO��pv+vP��+7E�_�	H��*
�4.�pr:�#����v�!o$Q���&zE^���u���H��[�'�Fnh��}����fE{>�e�������:K�Q��ߐ�&��50�sNi�����-.k��G��%ݽ��t�x�N1Yڅ�i^�����t8W�ᚻwÔ�;�d��S�Z��g�8�1RI|ld1M����&��gw<Ȗ'\*�=����)�1��#X�����u�iď��uC��\%p�C�vd�鹯��f�.��b��T��x�MO�z}9�س\J���R�X�o�b���q���L+3���>_��{69��҉t@�Vfʲ�=�΁Q�d�����������:���J?��چN~Lv��8��˒8� d:"Ol��#�����.
e	k����xXߴ��l���43QAHeSK87���Mzc�[+�z��'_�b����8C��O�\/T������<��s��0#ny�bct�5��}'��'��
�4�|�˫��8�?���7ࢴ�3�J�@<$���s�㭈���τSw��~z��r���]���9���mzh<�;]�ʤ'q�͘�y�:'>�8 �7��cD6�u������!2Zc��q��v� P�K��"F�\@x̚���Y��h[��I���-���W�-�c�/UOzA��(��g�+�Ij��������l�;��V�]u��y6� G����Y�B��{�/1��WZTsh�[)�{4�Dq��`+K���޽u�Zaoأ4���������b�y�	�T�]g�O=�xv|��������DE3 ��6V9������+���FNC5�>wH��s��v w!��J���0�ٱ5�a.�\��:'����<�v\��
�)��ţI��ڞتL0�V�D�b�VD���ıY��S"�Y�u���WGZ��$��\mR�ڗ\�4���
S��n�c�)�\���N^։�ç�Í��t^�=n0��>�J
_�������O��,9�j��v���'.2n��I`�'�7$�0$΍@%�h�q��`Ͼ��Mه�f��cx�ț�W=}��9�Z�����#'o�`�_�r�6�	�~�KpI�����&�����>�HuW��:� ,_
߸�A�,����,&�*���_�CBV����}1W������(5�h�X�U�5��{�H6<� �z�9�ϻ^�^gC��%,ɓΜD�O?X; QL����D����*�x?�lTh����܅���ʃ�d�sx�UQp:�Ci��r��v�Dɭ0�$�B圾eNX��9Dp�ė!���E�Ͷ-�	��.�G��3����Z�@c���=�Ɉ��� qP�
0�9�W���Nm�W���ڛt��F70����mU�&�9[{��� }�AőK�?���9��;��t�ֺ��|b�/����]lB�}H'�e � �A;�m����l#� 7����g�%����P���<��_�ټ�0��0t��\f�"�7� ��-F�� z:l�}?�n�?Ud�z+���>�ԭ�����S@6b`ll�g)�SF��,���X0J����R��c`�Ff�Q0W��$�;���ӍOZ+5��n*�M,�Y�M��A��Gȇ�����=�}�ն����Ѹ�@�G�����%vW�y�$�_e�O���X�喭��~������XH�'8}�2�	ŉ$`�[^�=n̺g+4�--�3�ͣ�e�@�'�v���/";��5$'5s*�q��h�)g�1���F�p�2R�ĎۢN�]�)ZD�{����|2,���Pa�Z��k`|M����]�|�m�a�E�e�n�I8f���5M(d���$ϴ�����;j��URaE��s�D�o#Y���(�t>y�9�N-��n%}�*}g��#7<FI/�uQ�����VQ�>5��&�QMTf��Dm���Z�M+BJ���+�K�$̵	w���D�`�� ٪�Yq�Im�u�n�b�̓_��ՠӼԛ�X4,�?�зɓ����ЅM.q��:�\�`�����cڥ��L����(�w�F?>���Y�����{��-��mjC��� <�%��F��w@V&���q�;�R#�%z.z�X��F|F�*�
�L���Z��[�:��]����?���Xi����������v�MU;�,�ԣ�#+kI��}����%����j������D���S�z�?���K+)֞�Bؖ�"=���S+_�5S-� Bv�*�o�=R*b���׻������	E[٫�i�(�=�8�sIREv{"W͸4�������y���r�\ĂȦ�} ʘ��:���bo�|�r*��6:5�P��ke|�n-���)���W�ԎKV�#�XC�E��)��J�~���'|�i�O�G�Ï�����>$Oї��J���G�-�J�e�p� MW_��Ҫ����ҟ�(�\�@?2���X��:��������,5�����!"$��L�K�I�x٥��Bc;Ʒ�;��-�`�׎�>��%�yU
��M�'xΓ��Fb���T��U��wXٛv��m�8zRv��"�G�#�-�EJ"���|g��"�bﶮ�ke;@ٰ�3���~���e?�]]���\�[쩧�D��T�{�	tF:pU��Ҏ�� �c��4�bF�N�vq@L�hh�=x�p��=mTc̯g>�r�-6h��]HN�Y<�M7�|�d�I�5ڒ�<��gEj�^Tߚy��´�m��q�T��i���;#}��_� ��ڞ�8��cTK,adؠ�B��\��V���E�<�Qx1��q��U~~V�v�o��Gb�,R�5
�
�8i�b�lJnbMw�1�G�������-h�A.�fX`�o���kTȃ�`�a�wX[g��3�vd��>�-kD��fTn�,�~���q�'e�K3�e����4���O��:N1�m��_�Q�y���x�P���rY�_�������鉮���{��9N�|u(Y���}l/(���p�1���֌o|1��!��WV����R{C�pK������E�_�݈A/���	!F�tG5l��>p���{���q��w�U"x�wC}0I9GǇ����Δ��x�����{}W�����V�ay(Z�BW�O��o�4eF�IzV5�L��*�1Hb�#��J�ౌ껈�hϔ��T��������i��*���aL]�y��E��wǘ�'�m W{H���ݹw'�Ҹ�̔Һ��mMz����F�(�	^H}�Q ��z[��:зTa��@=siq�т��{4���^7D��K�2�t4�♨���f%Ǜ ǝ4J�n�E�?ã���7ڒ�HWRT2e}s�1����;.�"��sV��^�کRr����W6HV���;&s�Q��q��j#	E�R�jP0�<�NH6�(���b�����Zl�  &��TL���sK���:ġ��$���T��M0��5ɗ��~������.�T�*f԰�Tn�t��|H"�>AX_�5��G����Y7a$즣��)1G�_i��������3�C6-�I&@u	�����c�K�&P��
d�q�Ȕ�6�T��vU��uڛ�:�r�ȭ���T\���bx���s*!b���I]̈��\V־����0x�6yx�S��ɓ=V�ٵ�0�T!�����#S`s��~�X��4:+�*�ؾ���@�4�EU�SF4.S�1a�ڙ�}	f�������bIH����v��m�wS2$)��\(`A|'��U.(I y0��7mHE��$�f���ծ�D4$�d�����aX/�?�@�y��o�:���}�3�=�v���J��n�	叟؆�uxC*�\-�&A���+7���f�c�Gx�=�h��}>u/�b����T/���س��="�j	�Y�@W ��]�'�q�����2������ʅT�Ly���T7��Eks.B,��.W��?s��=��K�{���(6�X	_ְfo���lۢ6�������w`嵣P�D�l����uL��lRV�/�m��I�}�;�)˾�vUv�Z����xމZ:�1�&R�B(s��={�o��[G����N�;���F�ӄ{˟��#�o�A�zj����@di!��}�U~?r���á��
j�6�����S����BVXTY��fA���ۈ=O�*B�Tc�Մ|N}<[T�����s"��\�ܐBH�gU��!�^����ʭf�_�]�����z����N�
'��O�Й.=���eQ�3��*L!x^�3m{P��p3V�ąg���)�"b�E#��b�#�Ot�Bw��4�vA�`���´���̒21����)D�.�t�?hf�f�����hS+��Go���<B��&��U&Bv@?}wB�؟�漃����X0R���Z��N��6���d/H<o������e1��-���5��T����柊���#��z�+\�=x�aR�_�ʢt���~���C�x`�V{�Y愊ۘ�cL�������?&G@�g�ڊ;�j�qmo�e5�*6$1�f�e7`����NZ&�X�1B�{5��]u�2K(�'_lu�ʑS����Ʊ__�	�᷒G8���I���ͤ����ex5�L�Y���y'�=��`�����2���!K�<HE9-hY١�P$�k�;G���`I�"��E�勫����)Y7�^a���}���&��eȣw��(���"��^�D�&v�i{gk�M�k��}���-�b��=b�5#{�͝e_��&w x�p��5���Oݿ����.a^��q�h$sp��O���|���ED1�L}�;�K��v?�Y�ړ�������J�)�p*��Iu�<���1+Ϥ�U�*�`�x�0��dx�M��{v#����̜��H��Sњ$�7O�'�/�**f��Χ}��>c�O>�W�"-���. �Mq�#�BŪuv����k���yp��*6Gސ��i��=Lr�����ra#��P ��L'z��Yvd�����Ʋ�[6�l$_�}��jjt�*��[�3{� ���/Ct��q�>،3����ѿ/(=��YE�:����D 7�?�E�ҩTp��Hg\����pJ��={��h����G+f@�F��ڕ�RJ)/����0�a�����`s�.���.����s��Q�:k�CB�����[��Sᑩ��w�w*X:�9��-��q�Г�켊��������2�U�}��s4��!+�g��RZ�q�F�����
�ˣI� ��%v���	6�J�'e�S鱹"��Q��휃c(�v1V�^�dr�{�P��A�\!����ݷ�ĵS�A\KH�?��)Jd.x���P*���9m�=�?d�?ʃ�i@U���`��q!d�T�u�y�Oă��6쟨�BM{�z��~�%�CI��K�;��`��qy�����&]�Yo�G�֤��gWW����v<��J�{��+�U1x�4o�%(kWfe>��<�� ��,����Wν��fǍtcp��]�|&���e2� �Lv]�Ov�֏V�.�E�tm8�o�G�A