��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8�B�#q�@�;<t��:�[-���&��5/(���{���i�S���?��5�c-~���*-�P�Ϫ���[C���Q���QpY�$;bؗ���s{������i=1��W֋�a�,dW��D��j�W-�e����1��ڭҔ����K�k���p[�Jͨ�bh�jݸ����	F�5��[�kKm��;���7�}žp�e��Q�_P���XU_~���r�@��W��v��]�Ƚ�}�f�I�\*|�;���1���m���P:��.d��Y9U�
�It�*_R�s8䘆�j�q�e�Xvź[{,3��x��$�����8PD-Odq��9�i��kp����Ӣ_��T���{��e��
�;����ȞrC��RD)/�@�t���;`Y:��gJ��;b�y�~���-W�x�?T�ʮ���k�ъ���� kj��X��7�g�Mwѩ�x�g���/���'��z��#�1y�mGyC���LT=�-p��O����kq:��+q�Am��e� B�%F�m�o�z�A�����J��vÁr���}�Ȼ,�g��^<
_e+�3A��P�ޟ�+�0E{XH���WW��X�A�n�k� �՚V��{�Wc�߇ç����P�5�p�jy3D�zq�Tyʁ[�<���q9��ҷ=)�]KG���+��}}�����
%?�J� W��yxyn~'�����V���
�c
_^��R�EP���ҧ��D�|$��).jh�aN<�5��	�9I�����t�w5U|����O�F6P��r"};T���4��
��a�vo�_��hz�����lj�ߜ06�I!��S��i�>i�����n�l��KP����c�cPl6���P��Đ�a���l<����%����,���>�)$�='�(�Q�4�5B�7��Q���y��M�k�?{"��B�����]�/�u��x��Bb�{�@^ߖ�W?��?/�u�{�=�8R:���%�mg�ݪ�%6���d���터��h��Ѯ������;�!�,UnK�a �����n!��C��I�;�����͞��)a��mbo,��K�6C�Ț��=�ԛ�\z����_1%���5��l��*�m��D7�тO3!�����#���aO5	4 ��&I�3�E�R(�	L�-C۴�rɞҟ~ؙH�7=��f2x��l��$F2t�Ҁ�����"�(˼$3ö�����$�9ց�Dk�oT�/\�{��^-�����<�G�����
�w��Օ�O@�>@>ٽ��E�N��1� ?i�%<��ϙ�͇��u��ؚ֬����udO-��z��t��lkPU�zvdS�K�X�x{�ʕ�� �t@8S%76���t�U�MLF[Q�dNt��E�ԞE�w?��i)T� ���!�mh2���}.x�#�~8�K �̌V�� i"N��P� ���|��z(�*����Fb�9FZ���E�D���V0_�'0:{"�Y'����\�����@�q&��[@}���3�%�`n���r���ΰ�\���^~C�μ.�[�-$��q�w����N��,0loC7��V'3m%x�������xA�1A��f��K�#З �@6��D	��1M�f�,09����p(U�m�J�k@�"����P���UD�JМ�&����0%���'���j5������@�D���
���3h�Q�e���	N?�k��h���kH�t~��Z���!(�{=��Y�v���[ �[��~��"sL�����t@.G
�"
j���*�d��A7Sß֏���*'9��Z+��U8'��o*`q�XT���|ȣ����kҼC(m�˅Í�!����h���1�7�4�KQI�J���z��҅�\���:~$�n�/��'�+8��Q��1�J\� ���>ݭ�~2��%�_0�:���^��=1a��d(la��&3E���i�k��3�gg�fH2�T��F�)�R�8u���w�D.t�1�PN�]�V �8� :Yy�gs.�A
knh:/��l�bʃ�i6i�~|�|�Z\H0�9�Sa����bd0��~lV:�Ek��~�����x>�~P��ڀ�����Y�<	R�@Fxm�9�H�4u7��D�<���ǳP޾C��?�CݵX!��Z]k�j�7������1��Y������y�"�Gg�FoJ��|�X��%����mSqZ|��;�0K6*����q���fE[1k1��
��e��OL�S0P��?,���,d���!�S˫�.ʳzh��Eeֵ��8�]a*+��_)K�@Mi����i���:h)̥���F�x�8��nWˎ�h��> B�� ��x���n(:fQ.�@g\����w���ѓ��d�pU@�Nڃ�e���_�x�vb/-wgQ�4!���{X�X�)����:�]'N��Ų˸��ʁaTW����k��B>b_���S,x=#<`ojOmT�����V�>x�pMP�
����qI��	�<�Wt�Z-8k ����;�9=i雟�[G߉zvC�u�� ��б�.ړ6�s^3�]���Je47u�S��a�־��7�����U@#YΑ6��˦q���i�������#A�����D�+q������t�^���6ٲn����u<�pA�mr��8���A�j�4dn�>/���	7rb�r[v�CR�h{}�*��lI�Y����9f}�&y�O�
�>�
��Qϒ	�@�����Oe���n����]�3�����EB��V¾�HC|�^�C��f$`�x7�t�>j���J����l9��|818���g[����u�����j9��5�Ҹ�>;J�]����ʎw�q:��ȩ~�i6�r����ۡ��t3�:?A62��!td�ۭ
rV܇��H_�nLvW�R�+L����1մb�~��O�R���[�����C%eq����]���EӴ���w<��f�s�β�~�idv
�[��x��1���T��6��?�����?�?������!�,r���C�g�ڰg����q8��u��@��Zү�(���o�^W"�y���P���	@b��;���B��0�S��vW��/�4l����v)/$t�g��Y�酜�h��$@�h����	�����7����̺�g�'�%G�Es�x����ȡ�������u��X�Y��x6R����PT��/��5�	b��`��~,�ܴ%��wc��xE	{�mlu��<j[�����mr���� S�~GC1���@*H�uޏ#\:�e���r�C/�]�D�f���2�zҹl(V��Z������ȥG�	�SbQ�t���f��"�y���j�k��NFf���*�3{���	&$V���)ɕ�_��[MJ�X���g��<l�����4&e�,��젔-5zd�(I����0{"=�'�3�5w@O�,}\,-+��-�O�V�哀o�J�eq��Պ^���>D)�K�[)�G�qk�Ao�\~&���Df�}��݋�%�;�7�����2Nt�ݯdM�AOk�0��g+8Y�}pGD%h�]�/�+D��Z����#Lhöt��ڌd#U�8#�r�*�r'�)�����/����Ax�����gXS���#2�5�-�y��ƙ��)(�)�\I�g�Yu�ND�
\���O���Ⱆֶ��@yz�M��&TJk�)̀���;!��{�}�F�Y�[�k����#� ,V�3���I�71*��N��gǪt�R0VYIW�>^HMS�&U��G\�lpU�ά�����mg+'D��8��?���ӏ�,mZ&��ψ���y���ZF�)��ש��C�X߽HW��vC
��	@���/V�)��6��3��<���b4��n��͙(b2&�謟��
����>z���8�n�*�U`+����v�-��2n$��a�# =5���K�V���
��e��{�\������O��o���+<����om�3F.5���g;�)$d��u�B��|�_D��hrSu�V�r3-��M��J��|���=~
dG�^Ĳ�HX�����z ���0�Ce/H��nkG��D�]ZzAN�2~
�dذ�\�ڑ$�L��p��x�C�d��
��ʦ���eY��8�6�7�wTW�l�>��J��P8&0c3�(�[�D���T��;r������C�!7���;�.k�"���RK�kr�-$�7Ȁ'UI�v��^��,ѵM� &�
t�����n�˖��;��bt'	�@aH��l�Yy�>ptU�o�|�lG�:�E����R�*��-�~�$��n����V&4yln�r��������)1��۠H`�V�U�qxPK��y���iUYhX��)���v���5޲��EULs���`�N��@�%��{�k��+���