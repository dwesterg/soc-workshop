��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+?�9��"qzC���0��tb�%m�o7�(Ɏ�u�l������`ڴgQ
w"%M|I�ۀ3c�m��r�����&f���v����f�%��i9>�*��6�-��k�IZ���Mڵ�a�a�xfH� =�A�o�A����͛VQ%=�	�@m��jA��wl���u�Xȯ#��.��=�#RR��z�����=����{-��r���8U�6��1HbE�4�����_�+hOs��!��ϔ����釐����O^�c�r�I�l3���u&O�OY.�wZ�8=�I�X[[S#4��C>HY`
5��{kZ=�y9��t�B`��$ R���y�O��HL�:X;e~��B���U��9���XX8fp�w����H^ ���d�W:�b�+b+ԑ2ح��%��xd~� �c�FT8}�W. �
�;�ՙ�3�7cБ�*���$>���.
*�'���Z4�4�^�֚ۥ�*�J� ���>�'&�'�s�0b����	�R�q�	�4��g����/�ºn��_�~��S�(�ŷ���tؖ��k��l���-�����+���r�8Y��T�\W;j���hG���&��1M����j'JBX����ۇA��Q՜D.����fL�%K&�j����C��e���jy�<�u����v�e�8%M��A{Q:H�|ئ���&LdQ'�)���*n��9��pz!/�i�R�.(��C�a��ڦ�; ��ֳ�w|���v�2�D͊$�F8�2#]���i�S���xJ�#���B^��Դ�j�7�Ry�'��"�0]�%�W�b����c���Ͽ��!�<�~�S���	�����n��Ӵ���ɪ���|��k�o��Xi�=��\�T=��9i�.�]2���l�U:��ް��y³0��Ғ�0H-A��+���׵/�N����U<m+M]�g�y5H�#��+��;��|~A���[Qm�Ɍ+�S���H_�ی%��3!�0Оڱ�(��,^.�I�#�Kצ��w�#h���Q��x��z	���W�_��O^Ex�`$'�ǵ�3�|tC�P�FC�GOhY�.�O�m�yv= V=��o��Mgi:�󫰼��}yn��c+�H[J	��S�=.:�vk�Q,�k䖗R!�^/Dv���W�_��Y���vM]5i��f
��-`��΁#���b�帓����wskc}6��V��Y���yOG�k�}y�]�a�]����(�1�q)�?�3`bz�Ta*��X����#q_>KG���O
�M��ª�Gd�vF��v�k=0~�=�!Л:;Z�@��t'&+PJ�`BzW���g|W�yh���r�3�x/9�i�,�F�+�I`�����Π�b�#=z�K�mF��V�J� O�XN��8�=�4=�q����Y�ѲDQ����IQ��y��zL��U��x>ݭ��3�VL�!�h�$��¤���5����Is��	d�]í��
�Pnۣ�WF�Z�k��9gA�o��Ǉ Yv<�PJ�U=սS�6|�aJ�9�/���Ɋ�+����ơs�q
j;߬JT盠E�[kX�m��*g�>W'l�]q@��olnD��&���Z\c�6��)�{�h`Ъ���(>��6�*��Ӊ�!p�u�xi1�U<-3e('�����#���׀�:W�O>�a4�c��!�zg�XOT�����-I����Ԯ;��g\>���hS��w�\}mn7��hL�/4����hR?HsQ	1%,4�k��{|��c��~�Ij�� ��ʊ�T^/ �}+{q�ReLSN�íj���E] ���0GHp�7�d�Ot��^P����`�È�W`5����-0���ڎ��-�� i[.~�.�~���l/U0j������	�p�]�1	�{��%�	��7c��-9|2�S��:�Z���������FL�p4J%��TiT��ݰx猠1uڕ3���	������#�I ��H�>���p��rnK�w
z��u�I�
l����]:�([|�V�՛�PIIi��Օ�����J�+ٙjh��7u�z����8B%{�ע�E!A(`N�+�ݖR��b.�#�Ş�������k\\e�f���(���<��SD	!>!�u�.Uw��N���Q����
7B��>�7���!7V���ȉ���;TZ�&}�
��L�`^��e��+Tܽ�iP�lI"�HB�g]b��<Ym��}���v����T�)&@��Œ�
\����!ܚ>�	�]bt~�g��W�]�;\+I?cFJ��o�.�1)
l�6?L{,g+��G�{>%mQ��L�	�]�������� ݗһg�-b��j�ן���=�r�n�>DJ��nOq�Y�˜����;��`���4H��=����9:����I��q��T�Z�����u�6����+�V���%\:6W�⟆t��<�Է��9��Wl�t{Ap1�R�<�!$ʅL�C�K�z�È~Ax�!rp��.�Τ@1ߦ\�]iR�z�-�ϫ)��1�/�8�?�ݦ�MR;�h�0S?,&���p�&1���K ���7�K0��;�S/�3S+�О������w���G�n:����Pr:��T���H[_��~de|_<�ES�W�3��/�mHu$7�ihp�S��aЋ$&~]����X6�m�[�8�X; *����PN<CI��Y�S�MʰIP�9*���d�H$������z�/�����`DX<�YzU}]	>�u�c��Gݰ�<�1 ����\n:��ǟ���.��7NS��'