��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���KN���פP�����DW˜������v�6�G.ˢ[Ma�R��o'%�E�FT��g����/�^�#�>�ٛ|��W�<�V_��q*Q_��g�W�Kv����:J��g����s�"�|�@����JD�z��)�V�6{/��m�8_�w�����V���)���M�"���?�
�Ic��|��0��w����]�����Q���b��]�Nn�%��@ێ����}tc� W���aӻ��i��:9��'Y�jz�����E��,��'�'�@�5
iw&R����m�������Øi�X$!p1|��=@�]<��z
�;P�F`�f2G��'�YU�M���r�:{�^��P:D���u�G��U����eg�J7ez���09��|�/h������{F��Fx�nΫ�`G'+����4�wcpSW�f��!� ��6�f6�W�BYB��б���+�p��S�e�)�Ս \���)$�Aܸ�X%?�m����]�%�p��s�x���n�a|2.+^�*ϩp�&,���)ߡ�TWa��$v?���0ßE��f�6,.PG�̱��Z�����"�v���$,k�F?	^X	`����41�/p'���II����R],�eP�ƹ���C^�1�R1�0V������PX���p.B
����µ,Kq��RG�4 bX�Y��(N�n��
���|=a�49�H��1�gn�Ifr1!�$�0�Ah��9g��ثQa����Abo �����\`e �5�q�@��Ҏ� �^n"��Q���WmL�d��?�������إV�g_�~�^�j�x$%\I�L��<1 �+�����?^	������H�Je~������C�)��4Չ8��{=��3�<>g�0-�%���b��d�;��Y&D���Y!)Q#4�5�!�"��s��z0�~ڊ���p����w���)^���"�i�1�nQ5FK$2{p��XY�z,�%�����&��a�#i.��8��I�ԯV�k�ZI��#W06j�*��<0aY��x�=V��%��y]�@y�
�u�N@I�o���@�C���Osq�eK�Ymz�bXY>ǒ�BhPV�Y�1��A��.���]�-�l����F�c�gik)�PWͽ�^�0	�0Q��.=H�� V���<��:��g~��jq150�����1tq*P�V$��U����Ɍ����y���H��ao�7K�oC�Ox�>V�3#��-cv����l0���<;�W��u,R��Ma;�Rs���`Kl][jN5��iˊ ����zm<u��"��zdY�h,Lc�Z+�Pi8��fEMp�}��lle�;0�Q� 蹳!��Aɢ@l������:L��'D��)����)�9�ʾ�)jy����z�
I��0;�O��=yNԐ�tmVC��:G�� Ƭ��,�9NX���[;������^�������븛!Tz�0���j�f*��-ei���n�a�ҚxI���'�ZS8�B�/8P�+ ��B��^������	�����jk������Ev�Y�b�7�)(��/Q-{O؛�p�(�I]�5����m[�\U�>���[Ó�A~x�y�C��˰��\�K���s�\o-b�"�����t$9�(���A�����2Լْ�/r|^�Lޣ���]l� ��;4 'ݟjPa��n��@�I�õ�EΪ^h�޲K�p(�;;���&7�����ӈ:6$.<�<��z�GfO�*7����{S��|�oc�������x_��d1�W)�A��yd!a��q�i̳\��MV�g	m�yގ���9O1�g��R8��q6���鍶������,�5�瀆�D�K��?�랆�����EN�
�5��#�/]��H��p �V������6ۗ95�ӄ�4�؈���}�?ϐ����K���UYRՏ�
����,U�Vĵ4��O<<e�j/��7��BĀ�H2�4�j8#��T]NC�xF��� A|�+t� �Q��,�
_��O&��5��Z㫎��C�,��B�ΐ9�׵��
򳂈��((t�C⧭(������r7f�B�č����8�k"���@L��䄊s413:��ұ-hC��`����|���s��,�|:c�.^��.m�;
�rm��{��tMտ"�G�����G�^��Z�#�>�g�U�Ro��2{�ɋ�XD��'
kI���dD��y�1頠����ȸ��S �q��pO{�;g�sݑ�d�=��΢Pn���3��
[�z���h�����e�fC�ց�Dз睄��)��L��o��h�N}"2ml�'�Csj�����<ݕ2�ǵ?����XJb�b(���9���w�"u�&h>�׸�GH��2s�x�f[P��ۓ*��j�x������a���%KK: 4���"��E�nJ���
�(po�'�<��p�?k4�:¶c"�cK��)s�ӟ1�몯�
%.�4Q�12*�u���q��qWx?&�&vD�0�Eb��h��f��U	��'V���o�{KY��Oz�w�\�JBܕ�x5e�3)0�vaȖ2#�a�fU�VX��8'��2��fIH���B��z��Ri ���B�_�4G�$Z�v��&;�,?	�H2O����|�;ծ.���P�|�FO`�W-��"~�![�qJ�/f��bQ�0�3Z��G��"�Xی2�*���Gzo�<%�L<���P���R��ν:�#|��YJ1��5�;�jx^�YP��B�b�]��h�sQ�`P��`��)��>)2	�.��X���i`[����B=���jU�j��0��up����I����|��A[V�j�&�����Q6@�Q+I�t{�BM}��;���%N�e����F_��18W6F�^���]pJ��R
�^�b�� E
�wP)gAѢ!z�؃y��������4�M%�S��7��.���f�l��2fɆ@tѹ����:��֟�v*�uƮ��J�#(&H�U�=7��&T�������QPu	=?	έ�xg�����LO?φ�g�������(�j�.g{�~��|z��F�	���M����1�g�6�S4ĆCd2c�?-��P����ޞ�+��~����jȊ�m�=���1ym�ƥ��R��>�%ڣ'�B�{3;�pB|��QC�����l�wY�~����f�I������4v����(�<�Ֆ�y�y��ҋ/���02��۰�%��ﾲxv��-a��!��9�#l�?:��*Df����T���m DKL��y]Ο�����TE{W���·݆c+�5J�y�KG6�������,���D���|�߷;����=��1����8���`���%K��1F������9����N��c�y���ʏu����nY��to�Z8��;^4�!!_LY��N�3��v����E �`h����7��|��ʨM���i�luK�0����:��a��:CV˖�Q+���;�M��|�?�0<�S����C+i�9Pd`����$��Ho�fel׶y����9����p/��2%ŜXkz�d�AG�/x4$'�v�}dϫ��3�K�7�giw�a�A`�NA�*%���F����2a�jz~���,�����-8~�t��r�\W��x�ҡ���UeU��d��X��u�s��"yR�N��h[r'��Hb�~������5�:�F���;"�y���!�}�.�0�7��{�txJ>�	f��ܼ�nG�<�ߠ.`��B��I_Ԙ�^M�X�4O�+�4T}}rHVq=Q�U�W�9�yjb�	p ۂP)?�G���.����XL���
�aF\�tR��<�~�lEȢ]��]����� M{����'|��A{��~�ƩE� �*l��Q�,N���vX���i���e�!��t��C��aL�U#�sk����]v��;���$��)>ɛ���+=9'�gG�l����Y ŵ�Q� +�^7I��ͯ2�6��������E��.�O�Y�~�J-��DvO�P��8�8̉�_�Ξm��*�h�y%Ig_6xMr�K4�(�*�楞�~��:��/s�"{D��A3�e�MH�!�8����M��R�*�&!�WD]�ELU��킲v��j��Aa��k��z2���KVH˒t�Au�h�!�3~^'%�����j}*�Η �4�@�H�d$p��,^;����tf����o��a�������O��jglM�@7�n�zǔXP�{Nr�p�<zk�[ON����9���t�ކv�NS9�k{��E�Ni��a�z ��𙿫>�\	Y���Jy�8� �}�H�i�Q�izk.�5���U��;��TX�ء�!0=�Җ6�s�*�O?�<n�5�kL��X:������O @I�uBe&4��9l���ږ��[�
S��V!�(S��j���&���ށ[O7�rK�����rTw�)������H�h&����5ۋg����(=���Ѱ�� Qf&)�XJ���� �Z�q�v-q���]�z��T<�)o%��9Bt������[:tk~Z,C/ߚ���^�:�%|�e�
��u���B�� ��6lL�V�0�gI�G�Ҩ�k���Ls��2>�s�>�Y�]E{�D�5l��s	�����Hb��� �:����`@�k�"��5	_��lm�W��r���[5|)�A�V}:D��.bw���o��G8���I-BMz�?f\�c�O�p��k�U�B��6.�� �a�ZV��^��$�t����a]+�0CH[s��>#�+�ݫFw�b�|/7��R�1B%M�QG���C�xm�������j`����Շ9�'b�F;n�y"�,7�Ǎm���T�T�I�cn9/�3��-�%�L�p����Z�֕X Q�0�~���`�u�Ì}$[�I�/cl�H�s��~����"��0˲̔pH����-70����B C�i�亾(��4|~tw@�����qw^����A�Wͤ�M ���=톭х=K뛰����'�G�d�����eX�e��vf�cW�5�N^�C�39ͱ�߄���AIՂ^|��99�Vr�X���]uG�3T�j���:X����+��^�(2EX�U���F`�h'�ҶG����<�a{&��Z/�.pI؏�{ 5BG�q�O�_P����x�)�]=o�XS�/�HK���$���rQ򿛁���T�S�-��*m7u���[u��a��d,H�3���!�D{��e�~Ƕ�D�F�=�G&4C����M�&c���cѼi���i��&}@+B�\�Ȫ�씧 Q˷Q� ��&l�������V_go�t:�d�kVYw�J�O�F��E���p���ihi�� I��4����%Ӎ.-�G�4L$�&!"C�Y^ʻ�,�����,�%O�k8#�j��p�� M��$J�#�Bi�9z�6
��L�m�3�''z�/�k=�gvL���s�{�G�iy�\%l/�'r�iO3��fr8�#ܖIlaĘ�m��?�h��L��{:f93zc�&ٌ_�Ҿ'��o7�%�5޺�`yj�����vuY�G�Y�
׵��;���4�V��*��a���
�E��w
����8u�?�߸#YW��/n c[�hO���N=с7��ܧ�<^��8���T�,Mo꼛��>Z�yCfּY��u����f�@Aa/�^P>G���!4����g�������� j��jg�rQ9A��d�' ��})Oy�y\�����	�h�U/D~K}'���hi _>��m�B�8��ܑ`b����ε��*��5=�x�<׵��8An&F:����u�O��(�i(uYF������͇}�~>�XȔ���/���5wMJV�1,�Q���`�*["��[#���FL�!�]�|��\B39�"��g����a�K�.�U
R��w��3p�X�?/���wl�&lU��+��g�j�m�+�"�,� ��&t���&&v;G(�?t�P)QT�F�:؈�'](� �P.��&@v���2>���DP�*o �>��~H{	�?9J�O�3�>�e)�EG����O��;4U��蔑_�xw'����@�˜��M�?��*��>@@_��ڱ�W��"%�{ۈ���r^�
���B��"D��F���[�ׁ=N��1I�+�(�/'�tmo���g,G��K�rB�3�8&���������^XK�:�֬�AH���fs�J�Ҳ_]����D�M��#w@w X�,�A��3�M3o�B��.��=�������&	ve�6�qZҶ�3����͂o��R�M��8���#B��bY�R$�����I�+Q�Q��i/|���ʆ�P�m�V-�7Ä�Mv�!��'��U留��'�ɞl�l�o�q�	�9�B�n�ϩ����?h�a����e������IA��L�dֱ����A�L¡G&�󪨥j�M�������G-4L-����z��A��ۢe�9�Y͇�/�qg���Q�M3*��a2n�|���:ɥ��2�(|x�'��z��|��|��|p8;-��p�vp,�5�v>Xd��]�I�X=`k�\��x2eH��)�����$V�����mE��Z�7p��������J�pM�o�z�Ѡ?w���t�qԢs�F�2����$/&wl�pf��M)ڻ쒰�T7N�Ib;k�!	�*�MF��;V�]H�~O��e*��"�M�)#+G�g�n�x���Q��.S�PI5�D�F��H	4�6Hx��"D�&�H�	L-yFOŹ�q�Q`T뚳�b�*";�)���>�k� b�3Xh'��x�FF���}*��f������*Y��e�{���Ӽ��uM����ŀ���2@z;��T���Ďtn����?���t+M���!Ŀ�8t	���!�4�y��[��m
8#A��u4��+N�uہ�ƣ�Ew��5�BH��+&]#��/�{�2��oK��5�m厘�p_�n�B:�.�������N���z�K��2��ӄ��'���z�}�vO�y�WN�Ⱥ�F�	��s��/��^y��7�Gc��2��.r�`�M_�$4����b�'���%t��$�'�8��<��k����� WAZ�z�]�M�n�Ю��$f�0>�����;��L�cT��8�C�流>��.�K�A�!\`��_�0J���95��9wj�Ӣv��;Z6~+��C�m�޶u��;�[�h�}O3;a*<D�ิ:{��O�Kcu���Kk2���/�yac8cq0� DT��߄hU�E�.;h��s���30�C�E�L���KX�t_ނ����ľ3�X�'K�	��^����{h'���p�}�s�\��ND۠�Y�N� �;r�v(�qN	��kv_�˵���+*Y��W|�]7>�oϭ��h��X�*as����1K0U��J���K���˙�0�Wz�2L�"���bQ�E�~a��"_��A(PhN�J�A�<�'��됎�7�+/>�����\bT���t�#S1��K�N�Ɓ�rٯ�@l<	I0S2�a[7/!,�9���t3(̀�GH��ԕ]ȿ�6��y��{(�Z��0;zK���G18J�~n}³��.6�_�����/ s��xYkJ������r���^1i	�`�4aJˁn�fL��Z�l���C�5p�&��i�eȅ�'�!��b_���<���N"�1'�D�(�(C�A��K1�S~[��l�|6:��i-�lx���s�.�I�+��ư2���l�����A�%s==�D" A�]m�|+uM2,csM'�#�[��������c9�-��Ƙ`>j����%L�,/�&	aU�������c��� 
���.�,�M�a'�㒠�/�d9����G�����3r���2*Ǜ(�n�JS�2�٨�.�ezS�m^S��[�L�9L��g��I�r�}��̆��>�L�e���TMσ��:୊"R�c�-Z��FG�l�w��M�k�WN�k��40�X���}skFQf`�=�	�Q������Mf�z4!��N(��8ߗd���bU��\Be:r#
bA)Ƙ)�A���� 9���CY�Z�������^��p�q��y�z�}Kt�غ������H���)�P��Q3a#e�E	c;�=$o�� k����wm�1,�()�
��S���mЈǯB�
�h�bѪ��TRJ��������>P�j5��3^�yb+(������Y�f��ʼH�b乊d�,��7�md��^����������a�"����}��! �H(_O!Ot���$�MŖ࿉�,��,*�Vi���V��w��Z����t�w?��W�Ϊ�ɀI}�3e��eP~�cLja��$�8N��x
;L�۩��?&#zjCmtQUW����e\�=�r+J�p�v6���Y��án�vY|�Ħ�n���R��t���7�S�W}CEs�����!]��o´�f*���i���p4���Ǝ.a������R�[�����֯��S\ki����ʍ���e����!K���ǌ����)vU;1
""�F�Y���	�Nq�k� ��v�"�{��4�17�����˾��ݝqV���^���'��,�qE�H3̅`�A�8z!�k,��3�)%FS���wמ�u��-�s�?�����k?k�4`��s�aȾ��"����
��|�󫲲W�AM^�b5��z4`|����@N���Ur�P{�,�^$v/�(U0z���Q��B�$��8.�{�2����t��Fו�[j�p�A�$���D�T���