��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�h+�yO��_6�o�7'/\/��I��K��vo	��L��o$n"�4�B��J��/k��ƅ���X��l-5�we��ڦ]0��F�X�%�-��P�E�s�X����ٷPڏ�ǕD��z�q8�M�3�zCvJ��H,�e
�*.�͈}�ak���պU�px��Y8Ӎ>��~�������)e*���-�4cg����ʽ=��1U�+���� `���N̓�a ��',�X���x�0�q��HZ���m���Âp2|zN�Ǹi5>qw��eU ��(z���w#�m4rci�.:���Ȭ�b���C�Y���D[BZ颺��S���y��Z��I�=/�n���@DwY<�5�;����@�����o�m�Y&�)�y���;��6QhN+��ؔ/}�jP��g�u�Q��\U�י����6�2H�z�Cz���gD�/S�5e��م����RV�Fl�������6lkF��!�)!H!���]�ѫ�I[]���པA^a�LO���/�0JK���vϻ���լR���q�9�Z��Q����۳@��+����z�i��v�إ	U�����WMy�r��K#��N����nwT��^�[X8������F��E/�[q�Z<F��I��#/Y���}9�������cøR�i������-�d��#�:=պ���(	1�K� �"&{�X�ܠ~�:��Y}>%�zA;!}��y�(2�M-�W��򝙷~�|j��l�Ǩ�	�V�ԙ�^�v�^�g(��؜�'c�;2_���⁛�P`�ӑY o�U��ʉM�.���a���j�� ��įYl���&�]��t<�g�?��s{�����-<�_�؂�9I1UW��_4l;px�j[�p#������xɍ@?"��,�$�}�~߉d�1lL��f��U��= ��Ǔ�bxle-�\�,�Y��C׉�o�heP 9wx$�a9��^�*��RX$��cB�1�E/h?z֣:,V4E����}֗�[S����������!�s19��<��~�B`�:�����ܢ$F�j��7�}�ѝ馑�M������@^__�4������1V��w	]Fc�R��������ӈS�ɴf`����I��]���JwB*Lwa��X��8Q�E�i"y/1�EĎ[���[dQ�D���H��a|Qk�!�C��̸+��r6�Ɇ��fD�dJ��2�FH���?VK���%M�CQii��7%�%�a��nx{u�Q�+ЛZ
hrf�	�d�N6�A��?l��������pl��<?��%�J�,Jx񄤺]�L�Ƶ��xZ�~y�1x-&���4��;[l��X��E"襏�"M�Ǧ"vIR����-'k�������9��!�yЪ���G��6��rf��|<��MOL��(��FI~���ڲ�h����i��)r�F���SCq5I�9���e  �����a��D�/P��5��m5m��l�տ/������/e�S���I�*7�˙so��V�]s���7�\՞�j��&�t�Yǂ'�p�ؚzIA���U�F��J`��5��
�����]��zK��)n	�5j��:�/}LtK����N��x�&���������Qb��6�2'�ʪ��������0�z��E����8w��G����0�o����b[�h3�� ݃-Fmk73�a]`C񔸪�5�^�]0r�qTI`�$Nlt���)��?���,�tM���igw��XDm�^)=�c�,��!T���-���0&�����%�W�w�pՖ�q���[��D|PQ����wL�Ģ`���#E�	�ߗB�\��jkƊ��o�����S�M*Y�s��_2�21����P�!�lG@�t�I���� �U��5�GO�95G�&�ʨ� Vqu�����NF����Se�$;�W'j�A\��>�te��e�%:G�׏a��������
%�}>y�a�3���2��{`9l��b��h����К�`�T�����������̒�]Yn�%���#`zv��=H���ToT{�1�L��-T#��
U��wEH�ron3�S�Z�xQ���/O=�x?7<�ц(y�d/4{q�v��CU݂|-8 ��(B��ȬQ}����w�*��
<�N��J�a,��U);�Op����>2Lp�L�<���<��ѝ}ut��+�5�2;��Xq�mb�vT��������ڟ�ӧ�q
�H%��(6+��6*��$�m�(
�}��dg� �d���>F�������rk�f��ԕ���k�������t�q8n�E(�Kz
��b�u&�X�%s�@����ba,h�~�1�u�{�/��z�ɐ�v_�bR�|�x[-q�0��2x���Z���a6ѵa)łO��͹��4�'^�c�M��π��J=>.�jN)�������U)���Ws�]o�Q2��/�Sq��S�I_M�9��5-����k�����E*�G��C0_�)B�e��� ��k���sT(?jB��gfI�@�C�r���!���b�������tqcw%��a��{7N/�R��\Sw���6��� tOr�q= ����ŗ��<��F�j}�t��j<�f�1l!~��ƐÂ4W�	@��[|�������US������}�OV�}D�JX�+N�kZ��Y��0+������)h	�����4������z���&ZGCtj0k����jЩKԼO@�	��0��O��d�$�e�kd��#{7��!]Z��!�V����lC
g_r�z3�k��-#�+i���P�c�n�D�:�8_S}��wA�Z	e��_��6��}f�ŘA��,��.���7�}�����&��K8Ii8�������I� �=Gk/�`�JԌ|��(���QTh����:��R��r��6l6�2��0�n��B���^6e
�~��"`��sc��P��#��z�ǚ����9��:��~F���L�v�����` r�/����>\�)!i��u8��)խ�1�>�H���$�٢ʹ�u?�Y��UN���s3�m_�0��NĨ��Z��ޒZ0���{9�W|^�����3 ��b���((�w�j`�p�M(��j��T��?
�3���2�[ڙ���ΕF��|ג���&[&��Z:g���rœ�U��S���%a�o"b���c�u95�K��М��
���rC��g��e���矋���������܋���A�pA��t�f������"����*�.F�_�(��膅����3,s�3�m�%�/��&lQs�6o5���T�A�l�7�'�