��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���d�P�0�W�4���Pvk�l�k�M{�uфL�8��R8K���YH�+�����:�)<� ��N���O�u���D��e�B
HQG]�X�	¢췜�FnV<�x����+����{�;����|��O���'��>U��%ӛ���U�nrw�G��1�8����er6��`��x��3��u��]ʚq�2�M��	�B�
�ĵ�ETGW��(���IB { �,���ϟ^������R�����s�q��E��4E�ا(�mKc�L8_M�E�P��5�i\ ��;JPLl�߿��ă9���q�l��1�6��=w��Wߝ'
)K`DG/�3���X�,�a�U)$y9�f�f���z4t=*�1г�b�QIm�C�>���ء�=S��͸�>k���)Gg�x�YU��s^�n-��H��(�!��-=��L��<�ш�9��|���a�7Y�$���͆�
�|��Rky����|�'4D�D�mǸ��yU}�e˓�W%')�ag�������S����Hё}"���h\B�=�t,�c�h�Cm���E�cI'��e����`����zE�ӕ%�v�z#�qC� ʺ%l�	�W�}&��J�+	�qeӺ�P=H����J�+9���	ò�v�w����&�)�#'1{��-�������7[����d�����^2,
���AQ�t@�z����E<��k 7*Z�l�n�f"�Ƭ]�k)U�3���T�l��kb�Aݼ:�i�7Ix{D�H��Տu��X@�N�d��7� �%�ٕ}��8���\�sA�Ow�K+r�>�P92��[h���JnƲ�2DJ^d�����fV(l"_q巻��*��)��#8-�3\�
���H���@Ρʆ�Fр�a�.4��tmvp8�#eBVAz��A�-��;׷,w�t�Ƿ[]��d�US,��oBA.~���x�t��7(C��L�O?�Rֹ�Q���y�$�WJ��u?�ll.���ts��%���$���+Y@�x&l]�t���^�p���0B�C�[9����Դn��zP��u|e�fՂY}�l�|�Tb�X:���{�s`'��c�|U�}�"����Z��t9�x�ն�q�mN�u�,"*]���V_�I@�ȴ���v��(Uf+t�gd��V��;�?-+$Zߥ�4Jh;+,R,{��p���Eɋz�����I�QI�����" ��F��:��aw�`�ƥ�OH׹�XX�^��lg�2&�:���$�G���C�O���q�>�D(�����y������$�;bE)�������]����G�-Z|_v|����|��22�`e�=�Ok����}��$��r]�����-)^�0���(O�ܜ,L�".�>7�Pt��)q��2
"�J_��5P��d�̚�R�)d&↑f)\�/���`��Q<���GZ$���^���&�o��
�r�f��Lꇡ�
�N��+�o �<��lkZ��\�r�F��#���yU��x��Fќ��lK+�e4lj:�E_43��zA{��b#b>�s%�^%A��T�9��]Jʺ�-�	Uǵj/��ۻ��L�_���[���s��4���s �7�ٻ�Q��R�s�i�+N���3�9�v��"J-s�Х�D�� �+ftpC=H����N�Ǝ�����R��g���}U���M{�+KR�6(au/j`�h-�S��w�=�nV�R��X$�tᒚ���Ë��*?��#�A�W3|Po�[�>m[!��}q���$�l*��obO�'Iݬ��cpm`u���Anƅ`\�o �ϕi��P�m�q)���5[Jmc��~r�l�ZL��~��
���3�e��� it�*��\-Eߙl�4H���-r�|�x�
9�_�tᚘ�և�w�GB(������$(z�N%�lSbX�Qf�\s�^��w���fCw5R��K �cP���5�sc���n�on�u��e�KJ-�C�R��A�3������k,��P0�d��t'fB4�j܋	9��Y�1`�w؟��Y1�� 1�TX�']1q�B%�ܼ����fyX���(�5�=m35��l�g��0е6>O�g�MN���] a�x��%��G��R���Y��CNIaH�L@/�s����iX����W�C��R�R���V֣��|\��c7��l8=n�X��:z2�v���"�٠?����&� �c)�"�vi�~(�������*O^��Q����[�Vl�<�|�p�u�4���hKY{��鱴��
9���o\�9Y$h�P-�0ps�"�~Ծs�g���B<�W�GQ����P(Y�b��P�%����C[0m����=����C,	�m����,�]��$Isn�~�_(�^���0��{O����7��5�7��J��v���@`&�HZEm�П�
�'�E�M�b����f��qV$F9y��y��C ����$R�q6���Q;B�������b��y�r�NS���1)�I]�ſtp�����V^+fq���v���
o;��?��*KF������B��}���䕔pz���Ci+u��r�,bn�[�*����gf�^�s�����ƷA'J-}~������n�D\/��,3�A�f����-I���-��k��>���|��`T�t�n�̭g_r���V(�o�_ >갦��`��"�0�ז��$���'SA���7��{��?[�E��t��㋄Jܛ]�#�i�I��.� ��~���n}�n.C��u�b�\2�q���j
�j�X��CK�7d��}x8y����!@'@����q���I�S�B-�&���5�tK���ƾ(�LS�e�N�G6v6�"@��I� �i��R�2y��+�=�rd1;s���ƾ���đ�Xi�5�bѪ��(�� ���x�)[��`i�-�u�@�U*VWQc�b�I*]v���{��b*blh[�G_"��Y�W��$ߘ�d�G�!a��)����M?kw.�j&��:�ź��hu�j�8oV�0�w��kF���0���`3��ς<a�j�f6:�Q�)�1����V��'#�����D�?d,]��C�(R�i�9P����m�\�k�ZrZ���s�k9}A7S�� (���0k|�x$�p)w%��l���]7:��9�݃�?K����D_=$%wo&�D��q��ٰ(��8�:�e�$щs��{%�8�