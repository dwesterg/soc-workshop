��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��tڐ�!��Q�����xZ�H��V�� �]d��� ��h�hQ�/���o�~�կ>?�5�z�+|��"D�[�!#��.J �SJ�Ҕ�5�Y7�0�f[秡3ڕ4�O�~�	����u�Q�Q�H��)*��V�o���}m�'_z�8�y�@� K$E�R�5^R�Ԇk2�vv�#�80����I��JI,3)e��	��	֢�	�W�k{1"^?����̚�3x}0�#��4څ�9�:������l�Ss�n�o��:��Ӻ�h�;��	⺿ob�46�����<�.���� ��Z��jAG=�
}���iW�Z=�)���-���;r�ƴ2�÷�%��������9�L86��v	*A�b#��Hveo�Sv}���6�&���d�/)<���XK{��aD=x`$V
�"��k�`*��P�I��VCc)NUN�_+�z�q��5�<^�1J�+˃*MH諲�p�:�ĬO�����t�T	�1�Q���lgj'JH��jL
�~�����餑�����YT{V�Smv��ػ)4�/[��`�2^�'(�!t_cv��Km�!!�n#Ŵ�Zh�Sv�2O���
����#Շs�c��O������Y���<���A�nǜa�r�0���8�?<6[{=����p[@�L��oɷ�[�z}&?b�4Y�h<���	��� ��<�x�QH��cC
u�?!�()���g��^+qdǣe�����/�״�v���^:p���\�����Y����%ɽ"،�e���>�'>�@�V���F�b�C*�\���DgT�N�����;Պ��w \�orlc�]>��=�=��/d)��̯�pzw��vbK���2о�k� ���ʏh�R_��8��Y�������o�5�?j�|��ڥ٭��D	z��Z���+G/;�j!R�l�~�� k�pc�ao/���1�/{����LK츚�|f]^ΛL�s�:�,�ks��-�Ԋ].���0e�����%U$e�X;H��@PY��靻$6�Mw|> *��X����>�����e7
���Fa� ��B*��
�6�,�~��`�����q���'��߿����;��4�%�>ߦ��7@GΖC�̆�HӐ9��3ŽGyf��\�Q12�V;�%���74|��Q喑T�?�1���_C���J�1x^�x�^!��~Q�+{�yńK�W՟豐Dq���v�K(�f}�U���uR�h���s�i�̢Q��p�f��@5fz7̶��{+#GK�������Ǘi���W��m�����㧬ʖ������l9��-uO�rf�q?Li�ʽ����Zt"��i�q,t��n�1(�zF�Ө�]��,�v�[��+�QxБk�����M��4���{󔩓�`��.��|6yڋV�݋�Jy#�+�93����!��#+�9���Vh��b~4G*B@��GU<v�]DZ� L�k��L��S� ����G+�
^.��I�>���0gY���,4���.��`�X+� D���"�؈��Ƴ
W��.D@�:E �B�YX���;�k����L�����A�Qb��Mr���]���5\����"�V���Q��tb���?�j7��j{"��tD\ѹ\� �紾OQ��^n��@�����
;e��؇�'76$z�Y-�zZ��蜃KV��B�=�q^�׉���"�JI����}�m�V�P3�6m�&D+�7�����RSu:ۛ�����eЬ�I� ���Fj��&��(뺿Q�M�Ga��G�F[��.��ˬ�����+ g�>�=c�x$Q�=�Z���	l�u�c�#Tڜ�ZDa�Hi�<@�8�<J)[�~2s��W��yB2Fԯ���4�����`	�:S�YQ��9#��fH�s2;q�G��,$rH��X���-����
�����{��|!�5�\���:X���i� ���X�9�C�����w@t���gU��';�܉p���I[�[�Nĭ��[`��}�q�s���9�j4�Ӎ�v��ؠU�f̵�WƐ�!��| 8���*}!v��`�H�_��J���T~��j%ܟ�y���ԡ��C!��yК�ߨK��BY�UM��ᖏC����xt
+�s������$2X8VZ&�#mW3�4�\Z�Z�.�9�q�ed�%{��NTt�r%�k��w9%�°���$^.s+��>}���;݃�97$o}���Od��秐���Yr��h��ʅ��IN�<kket]�+\v��7�T�A��f�*1��G�LS�	s)�r�C�g�~3oː=�6z[�7���5X�*�40�H�Gbe7˲/�~�'�}zy^^��i�\�܊�:� �pF�j���)`
�S4�P������F�#;�QI�#���Bε&��P's�(d�sŶ)��	K�OC���R/H�ʡ��,����y�S�� �$�D�'�qW��o��˚��DqrhL=Z�wv�Ǝ�a�.���T��BW�t��fz�ݘ��.�� �UT�$F �G����� ��}�����y�xoZj��
��B,�4�`����#�D��*J<��e!��e$���av�z�%�WN�=�q���pH$ɣ��=>Z(�Gse��ZË�W�󼪲��A6������J����k#J�Z�����IEX�k_p�n$Ջ�2W9?�4rv���yӒ