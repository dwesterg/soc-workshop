��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
'tHyx]�'��[������N|!�>7��'��5sA~E���fIx��V6�[y���L�*�bޔ���QT��,"��~�45P����#w��6ٴ�q����߹�B��Ն�W��Lc���h�2���ORb��Ѱ~�RU�Yg���p�m�}Y����H���UssV���a�`?���Ƒ�qj&���#k��vMq9�W����U��J�9́ӭ����Q/� ���N����A��b��	�i�d(��c�ZZ��\&��b1 �YG�6��N� � ������ŀ� �}��"i�����դ�/��5Lz��]�K�F��|��[��I"&ϕ٤�m"]�Kd�T+��a*Qnr��?�5��b���䲯w*C�
�tf���FƍZ��,`�jb��$m�e"W,Z2�Y}�����\����n��-�[�[wH�<��_���zV� ��%]���m�K�S gy)+�"�<F�sf,?1�_����;9�c��Uc�rr%>�h3�?\piN�P�)vP��*���5�?:�k�6D;�-K��*=��Z�2�I���p��ZV���Ҫ�ѻcSjd�Ц�O���EͿ��� ��.^J�_�b��6�y��_��̛���H{�[���7>ip��J9�s�GM����ӌ1�� .���f]��X�J[��f�hk�k���#Pd4BRFo������.D����"#��I�َ�"��B�?x���|ȥ�o�j�ͲފI�}z�l7�3y�ha0�g�]��&���5��b��CD��<n�o]����T>�]�$�c��M�)(\b��O�.�|9�U�2��$G�jػ=���2#�!Ĺ$-<Y�Ɏ�{a���6�%R�x��P�|P�^ys�&���A�i����B):t�"�<�0
_�b�h����9L���>���h�8���$�	�)GL1��5��u�)�������o��zϑ"u�}�O�n֋�d{Y�}��MB.���^��k��iw+��77�Ul��x����<\[Y�#1�^�Jw�*�JCÖ��=Z6��J�ze7䦏�[Ƹ�Q;A�F4��V��
�<�Jr �Ր�	���b�z���3� ��_ 0���������q%`��A��_G�
�1:��ҺւRq�:%�a:U'^X�_2l��@�u��vZ-���n��3���h�A�,w��&�8�Wޢ#��÷�۱��c&mo��Ώ^a�����y�֐u�;�oc̖��Uk�BU(8���u�&Io��9`�#j���d�"�����050qw~v��tr|��ڠ"��al��n㿘aAٿ�lx�v�Kx�]�+6W���t�>�r*����b�&�S����%)ȋ)wà��&��HO&�a�^�r ��c_��J�ke@�-��W�ڢOWM�l��լ�G��P:A�3C�ec >o}=����-p�Fnh�}=�Q:��Je�RG��`�*E�>����v���M���
l!�@=BOZ��hX�GKT�Uk�{[���}Z'Ϻ�=`�ı7�2���6F�)N�����f��K�pƐ�R�@7WAX2���?�����Z,�qؑ鎅�S��{�4-%ݔ��/���9��Ɨ��1��y��.p�
�8-�*?<ΛuE`�"�Mfܮ麐϶�w��z�\�S�-]�mH���wέ �2;�۵�zEb[���I�,7�Dx��Y�L�ֿB�O��Ux�j��~����ZO�`�u[C��B��v޷������u�ԗ���v\5���^d�=#V�o�,o�ņ�D����p��8SA�0Y�e��Y呋y�����//5p,��0�>�͂��U�c�g<����0㐝�q�R���e�ÿm^cO�߭��«��Y
����Vtޡ#X����s\�N�dyқJ�]�+D`8�ie�����-�>�{I /]��*�,��G����x=(O,�a�������c��ۡ�qHK�:��߮��4������krt�c�S�4_��=~Ϭ��Q���!=g�G�w��b��R;��+�X��*��^�oX�e^{pnI?�|A�l�#*-5�-B\䍁}�V���I�Ik�tt�2Q��+;�	#[��B�g��t�Ϊw(;5��� A6�l����"�i���mE��t��V6�����Կ%��"v���c���f �A1$�e^��$�6��t�׿�.O����&	�L:w�ڢ�����A���&M�%I�(���yV7��[#��R�zRg"jF�^Xr�y��q�
�� vX���AS�U�u�F@:H3l0A�ϒ�U��� �<rG;r���@��F�f�p�SJ4�hQ����W�lP����m@�-��੬\:n����q��7��������J�M+���?GSt)@0�������
DY���3� /��⢕�i��� ���j��+c��J�+q�l`]a�thbA���R.� ���5{�8C�c5��쀸]+Ku+���OO�ެ-�tN��K���$5��8�Yc��6G�oQ�\�:��o�%R#��7|��g���I��R��Jh��!���Ӳׅ��><%;�yy���n�H�4�Mb��BC{��	a �O&q��.c4����%)1�_���1�V*#�-)�-h��2qëc��@B�l���~K���3ڛ��U���P��	Xۏ����/L�pJ�������r�Σ}�}/���f%���m�L��Pp�,%۳� ��(��*2۩���T���1�Z� {J�WՑ� f�@݄����A�q�Jm�R�
,��):*Y�n�֑{J��i����^X'�[6�[{p��w�D�ƈ^>�#g��Z褭�&_��A*�(	��	�����
�ɸ���ֶ�*V=�;[v�}���pю`�Yધ��6ܰB�"ع�U�U�j��f��]�0#\����-���������.H�:2,%�q����l��J`�
�����p��O��lMf�r#(K���j�3�Qk���!@P/�1�Ud��j�L}cl\�E��o�rd9��o��*P$�j8�|?=*�p[�[~8{7��\���;�l����UƲ�6T5�L��4��]�t�͖�az�ec�f Cz��#�)��Ȁ94Dul����%���7��L@�C����+�#&KU���������2y|�c�@�<��R��
C�3���Ki��n�=,	�T�-mtC-���1� 3x���b���#O@ϛ��}��ZbE-ga��_���C�Β�{`W}�F�����^X�U�g1Է��ߑ,'�������
�F�䂣�`�Lh��5�-QK�^6�}g�.9�q!(\n����|8 �+^�~����(Η�42>���a v�ҭ��M�%H��(hL���8|ّ���3�2{�봡,��~�����s(�-S�gOQW�xj(f?�N����{��7tAQ_%t�~�R��D%�Y%Y���3S�~bZ��&W�"�s�� �����^�"�R�:/�h��g�c��4�Tg��#J�-~�Ѫ5��,��YY��㳅����#����>o��wӕz�1�^�5E0b)VJ��*ꖒ��QNJL���^s� �C��&�"�1�R��i��� ���
ܧv�d3�#�]�
6^]Ө�Gm��1mr	g�@���+Hkb�vU��	F�gW�U�=hR5����\B
T�G��;�
SZ�勃f<��29�4����(jb�w'G=�	&v|�b]�:�+�~3|�N2)��\zb�I8]�d��j��ɖS5%�N�n�7�f���]Q5���(Wht�����?{�t���t��z�I�<4���)���@�S|D/eb8���@��8��QL��� ��̻��֨%q���Hs�?�0!E��VHkE��>9�t���Gq^	����P��k�9��j|9�6��f�+)P�!IV�?����4������;R�� o{όO�r�q�N�]u���y�� r�9�����S����v�����H�~����i�<�;����b��K�[��������[���NL	���aw����"	��ȷ�;ZY<�H�m���J?V3Q^I*"��<	x���m�WJ'����rg14�+:�W�Gq�����kT��rN�s��r�k�}*2������2��ît��=�	�����χ����-v"�v�5o���`�y��,O��׽V􌐶U�=���7դ�#,���,΂<�?/�U@:uk~h��z!^���@R]��iF��K�څk�\6��֊z��&���*W������gz��a⇛w_W��s���YV����1	�x�y����i�~�o�K�k�-�\�;?��f~)�S%F��*�0�.f��c�����"d
��0!�#F�2�q�GlѢ�j"v��u���6�K^�Ef�)�M�����hsTȔ�K롚��;_�hX3IZ��WU�q���^�6��(~7��z^P��p;�G���+����)=��D�P��bN��� C��G�(����k�� 8o!�3�r���\КX!ll�v�K;�QG�+VKu j�"�I@��!���J��6��.V���A��ol04� $00�m��%)�nX�e��\`�F_&t��d���`7a�23"�~�Z��5�CAާ/������Ir��1T�����(\mL<���ۂ�e{��jY��
�F�z�'�k� ���jO3�*�Ш1�a�A=E��#��k�U{�c+P��Ȗ�4$�Ӵ$�6PLR�X�h��]�܌Ԋ�ߙ0��?XPB�!>���h��Z��{��ؓym͍�@���dL#2\�=�Ip4�ų��ۢ�y%�����7ˎ�2�^B�"`w��v�칸�đ�-ٿ�]�CQQ	7��WRt�N���_DbxDc\��f�"u����+�ܫr�1�q�#�.����MLﺜR'�<����l�N|�;����Y�O_�*�ؼ�=�n���F�m���~�ӂ7G�AN}�e�!}GKM���� �=W�23Q�!$}ʅU�8;�& ���Y�ıB���E��J�%����_"`��Q�X�r6h�A�0S=��\]-Γ�	�`����勭�)���kW2���1T�pS�Ԝľ{ts�^����̲�����
���͚Է��sF�i�� �N��H�I��?���E�8��f�v'�z�q��:�<�!l�G1��w�K=�M�a���A|2޸=��*��<o5�)��t�X泄�(�>S��oxM	J���5"�t����Q�50�۷,�D�A)��p����|�o��3�6ԆL��zKﻉ�n�}h���bU��Q`Y��b�*�2+��:yc�ʬϖ��y+�����2���et�NW3�`���_���'N�I���w�V��j�t�5K�@/	'˝д�ó�!�%�(p��D�wi"R����7�݄�=r�c��4&l�����}��R�]Y��A0�V*H���Lڱ@��5����
D�zE�8&02�}vg���E���-0H?b���)Cw�4����=�0J.�=�A�"���D�Z��'��QC?�r�*�_.'���I�_{P�N��) ��y&R�"�I��f��|����+P�2J�G����߸"Cq^�$�����:�F��t����� �e�Z凉���l,
�A�2��c`=�hs��d;�*�2.yqN�*�G�j�0}����ϺE�Pqw#7�)w����T
�寀v���ti����(�����>�O����9��h�2��W��s9n0{�R�!r��%��Twɡ���lw:&t�ׯњxl>�3p�K��	hQ��ȼ�j��Uz��$�z�\�?͖�v��ڬ	�^�2V��h-㝁,(�4m��'b-{T�͌�B�<���<�g3�rvG�hO�~��������xg����~uu�H�c�t#�oI���3[2G@���Pۅ�|�T��\���?��צ]��b�+&n���0˭H4><����z<�ݶ� @�a�p�a �Ak���P037z�s���(����� Ֆ�B�E��牒پ�3�A�R%�E��X3�&,M!�?��@L#8ntmO�viSV���$���:�>"���N����<�����X07f��g�	$)!Yx�p��zח�~�����'bZ�u������>�j=�.$V�:��>˕#3��͘=��,(WԘ��%���a.�͞�J���n`��T���E��D�(_������t���b��ߛ*�1�칈#���7m��0|��l����Kg R�m�J�
6�N@��0��❄�X���&�D%�fr�\�^̻;��C�dP ��p+<�ڷ�14�����N;��pX��^�'�u1��f������2a��p^��F�����@^6�↥N�Ϭ�~!+��b�\�1\f�����P�V/�F�p�ũ�Y��+�N�G�g�9�ԗe_�R��'�ppC���񋷞��4�[��k�-?VS��������&���(�B�ei��|aԽ�4� gʉ?1'Cߴ�O�{F(i�BTv�b�Ɲ��-����P�wA>�v�Eތ�{��Z���C��[I�'��J�W�u��u���2Dc|xѧ�q�V���_j'�ߝVPp4W�}���:������c��'V��	�/]��&���H&?������Z0)�^'�_@6:E��f�d˫��g�T����nCM���<9r�L���֛��m�������X��S�䬰V�! �d�m$�2����\�<pP�y]ǖ̟|�j��xc���NX��+W� MsBt�y��������H�R��S������mJh�;1��)�1��DB����rìX���8Ꜷ�l�PmgP~;�v�`�BW�Q��v�$J^��b�|�3_)4�N���nAza&l�z�$�A��9�{��Zo�V���ԦOv�G��WEo�16�Sp�P�^?=����uR�o�>�>�..���u�4��J�P��d�eqM;2�I������Aq�:����U_�O����E$x�=�K+w�X �M���
���6r�L}��UdȊ�kr���P(3�a��]��_GX�Ӳ�f�
C�K��88>uh<�K 4�.�B�x��ѯ*���� �\I*�k������;��s���d���U��ӫ1=\�l�.p��{+m�QJx�]��3閾;�������
W=�5��*bo�Q�ϰ�Ә=��;W10�֪@u¼ı�$w���^@p�p
֖D�w�X�o�aH��~��Ļ��q�$u��,s�ƙi�m,32r�aa����iN�7�ؚ�|���[)2�u��36�Iw�d�%�_����T���)�giڙ����wId�C�H���e��ӱ��$�u=�����@�`/(x��J���D,�f,��3�CY�;�<MQ�hH9�4*0�
ל��P�_�\"�s��9���)���Lo`m��Û m�+2��u
6?���q���x�&;fv3���o�fRB{ɽ{�����?&�D[�tQ��:�^��e���+��X!��VvM��"�wz[��s�R�_t
�y�y)��3a/w���:�MrY�n��e'l���N���m����ĝ�����d��22^�=�%͉N���`�m$�6?@g���#l���}�U:_Y���K�1�%L	~�(oVFL��|<��J4.6b���.�7�s�`W ˥I�,s������_���@�/ 
({��2�_=������P����Pe����G��7�ǚ�_�u�H8���3=^������-y������dfQI�Z�(�"	�M�:IN@��V��th�٨��jbs��+���#����@w���׃F_�t�/S\n�s����S�(��x@]�������;c%P�,@����F9(�)Z��W�}=�C��F0���9+ύ�旜�%0�A@��`��y��h1R� bF*�~��8S�&8D��,�cض7N���k��}����2�piζ�cB
C�&�dp;aE�Cv����j��0nj���Kc�[�����@byK@�!Z�L�j��6���C��@��ho���3���UҢ1��W��j�#�.�b���&I
x�8��œ�'��~ w/���*;a����J��=�L1�f�S"���<�����~�N��J
������Buy)�]@��$>af�ë=�L�oT��AX��ye0���lDN�������Y�g�Ѐ��&�����Z�Z�,�GuKg�^P���E�o�4�)�jj��Zm�!P�DU��[��S�mr5=n� ΣZF�n�Gs��ͺ`Ř�^�Mz�xrM���;R�H�[��ѥIp%B6�O�alt��pӎ�"4��(t~g��:I��Q/%��-��9���B$aw'{��1ы�s��^�:_Y坈�+@? ��׍9��ڝ g
q;�ދMԃV7RZ�o�y�62LQ����'�'[4�A�xA��X�ȠH@J	��NǨq���l{��v_N݊��H�Σ�ԯ��by�`�� �Y����iKZ�i>ݢH�X��%���<Ck��P�xb���(�}���V�8�׾~\,�{5(n�+�V�U�ᅳ��V/�����F���,G��_a�ʋ�У�c|2���*����,�s��8���]}F��	�W�ٮ��5�)G\��W��S�/I�Q| 7V(#uoM=��+@���U�|,�.V�n�I;~$AbmX�LB_��"n(>�[��](�*:��<�b4F;�C�٨�h����9.�Bwh�~��Ъ֦5�U��N_庤0��3��zߺ�MܟX<m�+@kH|\d�J����m`I��>��9F���Wm�z����F����b�^��o���L[,W>��t��4��*��:�X=�����kFg~�K��_��i��f���fr,H���q�ٷ���z����s*���LF(3he��>�k�uZ����g�_'P!L��;l7eq_pm8"��*"��@�\���0��b�>9����/X�ף�wj��a�Ģ���D�#'�& ���t >fR��V	��a��7)�\�=�Z\\b�����4`-�D: �^�m*�f��$`���h�
�A�+�I���a��7�|��߶-w��ٍ��̌�?j2D	�w�`�j�"�ܛ��@7�GN�m(��8�4�ؗ�8}�?BߕN�sV�d��Nr�-+bµ��f�x��vզ�'�ܒ"Ej���2�(��&�:,R���0�ZiH�ï+"U�e�q�K¼�I0�t��O���1;��lb��`OǇ-���?JO��:�<.X��dM��Cd�+�̩p���}Q�`��%���������}�N��X҉�#dj������H�1��4���JX�������<�mRӓN%q��6����g�C��,H�lc�(j���F��<�3?�j���h������Nu�,m�u6w�/$^Ib��:y1x����Ҕ6��-�=eZ�)|R�Q���x�f�@�i������7�>w&�i�����:z�X7��>-̤v��K8��1­o^HV~^FO%� ,]��?�e��?��+������(E�g�H<�~Z���g�{��c��`�w���Wp�?x�kT���V�f2��L�b���D���Q�Ūѫ-��p�O��K�'y݉�qb��iN�>�5߻B�~$"��d�/[�c�@��H��9( WU���}�~�/�1$1�_�{l��W�iV&L�~)i�?�ԯ���������a���}+vd/bk�@L�l����	�$x�f�%�|`4��� ����[�3.5M�}���f*r�f2��\T`h��Z�?�wW+@Ǟ�~�̚�b{�?^$���������_�(Z��[�����ї�x�$�X@�` �K���[@e����Gz?r&��@㽓��p͝EMM2���Q�.1�DQ��	{��m�K���8�p&�I�*V�1��W�-+������L����#�0
pK���͒28վR���8��^bP�Pn�!hϱY�O9�3�L�"0`���]1w���:SA>
����7þ�˯m���C�\�V]�Z��i��JN��o=>�U8��=�������ލ�"\���_��v4��S�	XT/�ȩ�����2���]zA7bV6�ġ�Iq���4`��-��q�xV� ��ˏ~��[�O\Ia�ĳ`8�.�lp�
�#�%�꺵qRP6[���bo��]��IyEzF�o� ��v��x��NU�r�5ބbzĦ⟦�= ,�c�o�c݇o��|�P�;8;�J:����gu��N�+8�B�����e��[}��r�N�V0$m�E�ф|���mȽ�a���"�;7�X �;�A��5oM�Y�9��� ��X�$/�~{ۢ?$�ndpq�/��O1'��8�qn��|����������ʇ��Wݙ1��Ad��e�n_�>�7
�`~��6�����f�1�����+0݉ș&O���:������rY��]f�� f�ݗ!Iv�(�}������C��b�iu�p5�`B/�WuuJ�Yo&
Z��]硕D�U���y�~e�w�2K ���i�af�\���Mbt�t�Rس1l���z���(�j)�`��#�4MQ���nY�����=�``���
٭=�DD%��FX��w�IVMBl@��.�
2r�'&�H�wQ����#%t`�z�]�3��'���{����تgm�l�D�D�xvr���Cq��9t<���� b�x�Lü��ժZ�& Y
��MhS��QP_�H*f�(�B����b���
�&ӅQ�A�l�g������[���yVP�loᱜC+�r0?\���!WB�s�,��Br�����i��Y�fq����єhJ�G���{̢S�c4Z��w�� �N�z���]�0t�D��%��RtIq���Z����E�.�H	g��b�T�U���q�����ok���rj�l(/��5͐�f��x���ȁ�s�$#X�h�p/!]�D���ŀG��+ށA���N��ix�Ո�?���B���s����³NE<[��'��	��b��d�hqT����S���-�c~�{�[9?����Q�b�zYm%�F/��U?��VG\x5H�p��������P�Xk`���Y�e�С�j��;�FyF���n�����K�
uB�g��pg��<B�	[͇A��+�i?��^�س�/%�.���ۉ{�a��P��IO[���� !���R���Oj�\�NEEzZ�ǆ�$ꆀ�E�6�>��Z�^�o䓧~����j">�|��T��tk&W�2w�5�ТE����ILo�W�拒��
���]���b#�hsP��¢�aՏ��s�g�H($Q[a����k��)�ց6p�֣���%�������%]qwIz�eG$��-�.iU1����C�|�>i�M�����y�Қx���O�%�ȶ,� �~s��	��
Z��5 b ؉�(80��>
��E��$�nL�p-�î��@�7p"������b��Ie	�;�����B���h�m�gA�@6���ُ'/����1Q��I�#�Y�b3_�7i��+�M�K6E+p�(��Zv��ܮm����"NB�ߗ�[A=�G_�|��p��K9Hg���n��SN��->�{���{���eJ��5}%ø�ZK���_�-��a�~��C�X�<eV����p� (Sݗ����*�b�(����
p������!ƚ�N��[�����;;�o{~O��iu���@����'�d�͢^*û�_�{뇁�!� ������	�V6--�[�lQ�_;�D6�!�-yF�"k�5�mR�r���vq�\�!_�O/h�^�<�.ٲ��$D=O�cE�rƝp`��>/��,^���Z
X
����[�Z��?a�Y�@�	�(m�N$���dͥui��)�<9�jv�H����ڃ�1��r���:)����5?��T��Ac2���A=�O�����*a��Mezw��2�(����_&���b}�����pp�U��3]S�!��:���S��XLQ�\�y�0�s]n���7�#q@���������a(IS��L�F�Y_ӄ��si[��qAٹ��/<��� kz��y	d?:L�����"|�h�����a��e�m�����
)��G]�c����>7�-����7�"��6���8�N|�Cn�+����4�8�Bn�W
Qɚ��3����!��9~Z�ɮ�ݙ|���=�R��X_�:��F��v��Б���e�F��B܈y��mŝ5�B<C�[R���9W�i�����}Bo�~�gq-zE��H��=���~���'�. M2�T���� ��B����W�1�M;=�����8O�2�O"�>�� )8�"�����}3�,X�5���"��Qc�k�R��܈���F�^ǃ^�x��;}p�>�� �d|�W�$�� x�[���-a�w�/f�����M��``��*s_��1��'�����q֛���T�6�������4��"8��r���K��f�[c,���?���m��}�����:�PC��m �d��a���Vq�/j�4�����u�h-��c2��};J��=o'��ߓ���>�L�P뭘�c=8v�b���ܽ�5W@)�eq����]��	�ކ
��:��{/%��[,W�l��Ga�N�A�z�nBЉ�5�\8ĥ͈N``��=px�7�����i�ïuU�_7An����n�T�˷�e�$��ShՆ��BY{�N��z�h���.� �{pU:.�1�;ī��b�m���#E��7���6�rWA�����nVc8�8O� G����aQH��h:{���>g���e�%�~���g:3���Դ�칮q[��M�������%P��J|�>ה��B6ڍ�a�E�K������-��D�_����۬���N }Γ��ћ�ô��Z{��7;j�|Xë,���=�܇��dS_n�;&ö>�.�Y=JQ�>�ac�"Y�e�}�����c��aA�HmF%�c�U��8�tԻ	�׺C��˵�͕@�hʳ�`+>��Q!L[.H~��2�M�ӆ�**�nT1�w����^����ڦq�H���h�Yߟ*�l� �>���h'=��O@�#jV�g��nv�SR�4+E]FE#����G$Vy�n^���G69��7E!D �IB�W ��c���Q醊 ��w�Ai��b"5M��z,�ښD��5���21V�ƛ��gBUK��Du+���qNw�l����M&���򥼦r'���w�a#մӄd�p��{a��t=��ԡ�qp��r�K'����N��{�;
<Y"�j�Ȍm-'�ɗ%|f'�9ڗ���'r���W%��8��\b�Ъ=��mȖ�0�W]Ymu>�|����ѱ���BhȄC)Fs03�6��>�x�9��~������w+�ءR���E����Y>m{�jL4c����R0���e ��Ju�	d!T �X� �?��+�4���K{�Y �q���᠋�)���29Z�����ma���o���� �n�V�,�+�z_c�r�T�@ö�Q��[1%���P���Ci"õ��#��c��t��1�&���|���ߜ�}b:����[���E��[ �AR #f�[Tq-�Ӡ�V��#D�&ȕ� ?���KY�7z*jgm�M������(�O㱂k��
Z,���<��En�o��DD6�z�Q�u2C5��0Cbˍ�yĦk-�<k�H��S�J��{ ͪM���V�7[@�0����y��Ք����H���G(4
�&o�����m������i������}�6�D!���D;��F��O����0\�ǟ8O��"����qGmx�f�v܉��n�_��UF��A'�k};`5���ļ��A5����L��d�a<����f%�J�O聋�����Cc�ج�����Le�瑾E�ep��n��wͤ��u!z5A�f׊& W(�+v�����L�֬�M���>��Q�F�|��܌/`�z���/��)"\�?���CVJŘ�W��ǁ_���*}�ln�� �3[��`��ue�D>��W:���F�ǭ�R���z�7J�ש�V��	Xp�:Q��[b�X���3���Dy*>�n<w"�-eH�)F��јT���)X��iMn�N1 ��6'
k�4e@y���xȴZ�0~�a3�N@,�PH}��e$�v��b���"���r���u2���AfF�	{V����U�Gr³B���?�m��n�?��T��$A�M��D�\��>�hXa�����ǡ R�߱0�Px��E[K� ��8]o�c��` �h�	�Ao������S�=m��^�b����_�r֛�K��A ����P�I|�������_k��j�QC �6� ��N	�N�e���<_ns��D�c&��;̱���'���C�����4®,"�6��[{1���~o���|i�l��mca����A��*�o�ʥ�Ut�NFY�O�2̎2`yO.
_*5C3/�(U!�p�Q՜��k4�Cdk<p�*�4�����6�e�N3�x�#'����Ts�a�0h�,���^�?�42<�S����m���=���Hݺ
�v4��hW���0�����h+�\3t��@}k�׼���E�|���ŝ*l?�Z�V(2��~����T��/`L���7Ku�CJ�%���4),��&l1�V���xl�Iہ2�(�h%[��5��t<<�)�(�sCc��i�6?	M�DcUj��%�������tY�v���_4��S� �˿�3�ެ�.�f����į������/�N�,��d	�Wc�4�U75(l9��u�f1�0?�
Iu�i�+�:�)��Z���)�3!< Z^q�)��~���:�	���m��V��xd�N�oM���tz�@��A���"mz�mg�g��6��ѹ�㺾�"��A}�M���
*)u�
P�O� �G�wd�XT�k�Z�*�HG=��P�T�Ij�cu���m9fk�t̿�kl������uZ�V����V9������]��pLZ�1�D�B�.>\���ɍ�M�v�uǕc�(��3�T����ڐ�,[�r�w�Խ���V��ET{�N�3��(�s��#��n�1�}�P==��A��Y���I�S������$0��3��x{�]AZ�ɶ�{��=`�`l~��o�R?�-�H�Be�~��ӟ5b�x�s��3�&a�o�bd�h%�����k~�2Z���vR����~B��TF�H��j׬γ]bgo���l��� r��,r�C�T���a���-�o:�HĲW ?S[yEÏ�`м'���9Aν8O-K	��k�g���{�'�i�ꌺ�)&ebIl���S-��I-���}>Ɨ��.Z�u���_X!��X&�3�@��Wa(b|,c�wJ��O���u��(R�l��ʅVN ^'/b�Z ^�w���6�H��j��_�K�7���pQ� �0�x�^��'�, ��ľ�v@����\X�c�g��2,�'t��٤���M؅n�a�R��"��<�����a���ٟ��S��*ɉqe�ϙXU�4r# l�B@&3�h!�7y,V�dE��i���"�s
�G^,�'K�p�jG�N���b��G 0��:�&db�����]#!1�-9k�?�������53�lߡ -��{��Q�����~�nc�2u�����ę�⦰Žl��A�<
k��	:n�F�-���k��Ӑ��Vn���F�}_MvsI�V�r��cN9VӰ�L��\�ݴ�(	�f��C�����X�R��ę���P�3lɹ���%���)1�Q������Dn~m?���Aڀt՟�gBc~����I�lc&�|�]�,}F�����#5��vra���>{UhB�aׂE,W�9�H(��މJ0w�t[R\A��\��@�VY�Y}�"P�i������v��f=�;�XPj��tx�X���y"`8���	A����q�b�%�Q���L:��
]�H4���0�2o�F	?�����q�x���ũ�9wdt�Zp�h8d����!�b.5{%�g��J�}�3RO��JA���h.�F%4.�"�ОC	q#�� ����=��y������{� �C����y��c���-�����w�q�ম%|H��0����Oz��5�lq5DΛn�:%Ʊ���?�R2ٸ$��ɸ�c@P�#��CVȓZ�-~�ͥ� ��}�SXt��x�2�p�d8�~��`�!�qF�����(\�A4cF+\�Iݳ؛m��Ӛ����B8�Ѕ�g8�?��}�yn�͛�%�j"��+�\����5k��9�,�����?
"�[���^:���P���)3�S�o����1��`��MkS���dJ�ħQ �Sm�͛��J6�l pOG�ig�:��uH�KL��������<�:~�j�q����
�V�,��mWڭ��	#^G��l��Z���
@<��eF��O��}�f�-� � ��1lǙGn�>*�ɤ����ӑ��-��wU
sŜ���<jl�J#ǒW��&���D�s 8/,:�����ۨ�}8։��֡u�������W�t�W_�:0�Gɓa�c����VƄZ�O9�?*�E�]֕��?j|1��ՕG�G
�VKq�B�|�l�u�������e��Q��~�c��i�U@h�h���
h7�����i_rI?�=�Zl�'>��ι�B ���ɿ���%ۅ�?�y�Y0��l�����_	������A�-����R8���0*��'�����\�����֤�� ǭ�g�\�.2�x�Z1^�E��<"Vc~@x@��5]Y���me�s��?�
|@Xތh/o'~+O��&�<*�ב��9ֲ�7`�G�9������O��_��3��#�`��/�ǌV񣙹�m��u�J�9���B��p|�rCp	�Gݐ�L��<�����l�t5����>�}L�XY��T꓍�ҫ��	WG�5�i"���֡;����[.�ْ"�{qL�Y�(5Q.�y�7��������?���t'-�x�->�=��`���g�zol�e���w��L��P�- �|��L�.&�G��ёfP�:��o6{��E�~P�u��"m�:���{c2`����SF�#��]5'��	�{baٜѝ�o,}i��K4�9��5>l�{�T�;�űazfuhq.��N-�!�����az�d�����c�.6w�#M�,oU�3�t�h���6����YR8��*`���Q�"�ieA��:�KtsLH��r���i	G��T��x��c-��C�C^����,�|V������Bͷ�֓0���+�8b�U�b�W�|U"ȳ��An|n�y��[��ms�����M�@Z�{k�� ��	��UCb��ܟ|���|k<k�Pp�+{��{ʢ'p}�^h�c�&�zRZ�U������e�[n��Cv�s..�U?�;'�Q@ �$��:&ϓ�а�e�o�����}!�
��1<�;إN�:���k
�b��ؕ{Y��uiQkO�L^�m���\���}=݃26JL7 P;WHCL��7q.�M���ۿ�釿>_Cs����i�� L?c�\�ϻ��Ðy�g��c8�)P4$����<@i����99��øPB���J���/�Ј�8?��Q�k\�Zꐜ9'pe��?|(Å���E7{��'oz����pn�5����2<)$�/���vӬ��;o�7a�e�\1܌T=6�������&�	Au������:צ��|	�����3�1BG�o���6܄���lk�(K����E�݂�n�0n�\�+c]<�o���|DU��oe�$�c5�����z�JJ�YK`ц������Qt��0���̪�}W���]��;|�1��!^γ��[ 
�q��2e[�+PR���P�.��9Ʋm(�'K���j���䍟>�����o�����J{_f��I�d���B`�V�$dO�7:Y[��L��S2[���N�@O.iu��1��H��[�DL��Ĩ)ޮ�N�zR�)�"�������=����ڃ�.��ih��Τ�*�!�l����� %�M�=�v0_w�v%���M�癷C#���f���w��wƿ���+���A;���n�C���5����Օ�L�H���%~���le<�9��
�nA�w�ݒmY���@�-�r�<�ɂ��n�%�z��\����߶�� �+^*���8�� �/s,9[���q�*-����v�#�����L:	rsQr5�s��/Z���/��������P���G71��^��b��2��(Jpy�d"Ak�LX�^+F�6t��h��Օ�Q��ݫ�/�I���nj�i�g�s@YSޢ�j䅶7|��T�)��~���3(L�}�<Kv���J�A�%��@�eb,�P.N�����^۪jϮM� }S��� w��tUd�#��x�xgI\�<Qد<׻�T½��/�C�<Y�\���J~<�&m���9���A}��+�2�^&�Je�A��Q��5l]�2T/�j��W-ݳp�O��8:h��3�mw��CdKr�3���>}T0I�	_�2Rx�Up(�@e����0!������ut6��� a���}}�\G�o�k���unժ�Ս98���6rx���ү6�@FHt[�S��Us0��tRTEd7�!k��zD���ƛ#�rF�x ���	!J^(5Ϫ�V�ۊf��Nt��f�J^�"v�N���.t����F͢�!��]'.��o	�GF�g�d�j�aVڎ#�&%t&c�Qbd�w=�}�w�K�PsAݜ&�j�Q�)�EM�W-2�$�'�$��$n�0@�}�s�u��j�u�Z�'��o��@�
}��tR���p�4)s�6�ĉb]x)�����rz��J!��D�w�5P�8��v�����8��C4�����),쓣`w��Q6y�i�O@,�?���L\H<���I���3�*g�i�>*8�l�G�}���E��D�|�kkٟ'���S(�D	3�u:��W��O�"^6�f�P܁(EDQء��:ΔDT6X�X	h�:Oj]#@t���Ԑ/�������F%�|f��֨�=�O�4js0�6����ޟ�|N�N���G;fH��z����]�Q�Y�X�m!��IB*"订��8��N)�"��<�(F��X��}��%0���f�	��y���n����9l�ʥѡ�&�A�m�oe�վ�
�JC�&!6���f��r��塤���Vdpk=��1}_�!B����O�E