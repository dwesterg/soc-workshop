��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd�G�'��"w�$���9���++�]
��>j�(��W7�q_���o���}�ghGz��@���ɃY=�����VÓqT/=�>�ނ��_��'��G$�P`:$��3�,(�w�w�R�\v�P������`����u�,�����~�׸���/cU����Ѐl�2��'�:� �A;�M;�S-3�6�\�	� ������ ���yް�h#�7b����*���$n-f�WCF�M}�)��i��ߏ0y�'aUG��{�6 nR�w��h� fm��}��D�'Fr���a��$X��߫��zR��}��fl�@��3�0U\9�m5�)Q+܅��	Z%W�5KC1q����
U����Y���Py\��İ(�į��Alr��L����H��}Y����1�r�G�4_ &�Þ������2������T�E�-{л��s��-�S:�C��(�\���I���z�Ll�/R�d95���J�@.!Z�`O��~]��T���5�@���W}S��|�p�����֪��,,(��~[��*^��rR	[D"��,�a�!�����7e��BO�����=C�J�f*���[�/�'�T7Uq�	D$� �Zy��&O�f(�IxiS�A$�y��X��V�%�;���nblm���r��1��ޛ-@f�:)�g(ZO�:^��]+���=��L}s_�-�����|�^����Pyg��s�$�$��Z�	�^��d4ʦQ�c)y������(�%�؋��SLvٍ�%����"�`{�.�a�-g��� u j�ph��vj�����~��H���r��p���H�����	+/��DX�4NN�?�E]*r.aq��o�:E^�E�:
o#D��)�_�8ĕ���?�:�2؁��"���楱���������E$��nK���7���D|��fq,j*���$W������í#�':�RׁKR@�?�^|g���^>��"�0�g�`D�p���y���!���N��=�����>_89�c�o)?iY�12,�6�CՑ�eT�!�d�1���%��?s��'vke8f�7'�j�O�J�DH{P�۟C��r��T@���ۇ���@��|�X0���T�9�׹oȬ,�|����H�K����2�kd"s�C�3�AB)���e�h��Xe��T�Yd���Hp�Hzr3/mC<o���J~KFo��?����>�l���5P0zw��:*)jb D��M�:2�����c��O㓘~����I��d�B�^e��ѥ�y���+x*�	TV(J�>���u�1���m�:^��� 2G��Y��t�UD+�9E4wC{�VD��x���m�A��dI�Sa���i60���!��k�G����x�r���l�QJ(m��$��B[+��Q�qF�?9�����A���*y0I<��� �j[�t�S�o�䖐�8�z?��Kϸ)�F��̸G�!}$\���2B%�
�Ϲ��}Q/�tW����
E QTx�6�1���pd�6荖.���j���_1_-�ߎD!�>�B%�|6	/>����=���k���Ե�)��n�0.�67�?��?�͍��
��=+�'a�U��Cl��ղ�a>��.�s ~�����*��q�o�|Y�kk��<YX̪t���ͩ�.N��0-�9pRC�>.AŢa�� �F���o��VA���fݒP�{�^c׬B�V$^��#�#E�N�Ԅ�*!�0�]Ѝ�Up��#��7�"a$ ;'�b�Qwk��3Z�q��������?�Ʃzj���<��=�H�θ%{ @�]ٞ�5h��f�r�OFi^щe���
-��M�⟌�ӷq�������q;;�X1�������\ݳY�1*!�/�,|���F
4��PM]\Vrm3�������m�T�$�h������ꎸ%Y[��0ϓ_�����tk�8jrk
�9�;�FZ�`�����Dˊ/�qj����w�k-�;���Gk��=籀���ҥ䨢E����cV0Z�6�]�t���q.��R�yS.K>`ŖT"�����@@�Y���kf�+	�i�CT�����S*�q�?���BR������+�4׶���d���C���#i4�(R��� �'��+?�Yh	��:�$�4�h�o	Y(��$�4�J��h��&�;��Z6��l����c��z�-�-ܸ��FfQ���}�`�H�l��R�S��;�y1��;wd�{�@��CJ�ƪ'�J��3ڱkK2L��馺�9�33\{\ǖ�2��JM%ҲD��/rE`�m5���	>�L����=+��WM��",��z��#v��m�"2�lA�s�1ZeGvӺj,ƣu]b�D.?~��ͷ��a���qԞ$`)css0Lw��srԮ=K� #Ш����yT���6ؖ�[x_���e���W���m������h�vSs4D����j�n�F��1QPR�^`�<��T�����g,�?^�A�b��`�f�J���{�+��tl�u��V�;�*��Y=��K�D)R�k����Ɨ�@e�^��yEo��UjK���.2��암��d0|X�S���Pi��p}�fUn��x�y'��A8��	�y;���EE�6�Sd��X���~�X��uQ_�1\RV��=Lvj�z�8����:)�+��wa� R��siTG�|��T"xJQ�͸b�ݷ�UG��:Dc�4������:�H�d�ۮ
�.������0��a��Ԛ�X�2\&-���:�����l�l.�/c���_	)a/sW�z}xFb� 97 ҏԈ�[�?���9���okvv�Q�؂���֚1�Q aݭ(ذ	A'y���6���p����B��;�nU�?"��� Ѿ���_�f�-�{�w�o�#�#���z)+kf�۩I)4C��λ�;�����m��`� L�oҭ4)��2ӓ?�ݩ�L���Y���e�`�
��C�Ƽ�l����-jk7q9�f��!���y!����zs8$R�z67D��ʓ0����$�S����F[n��N*�ۥ�y-�"�>��4�3_�R��BD2V� h���Э#)��uG.8���A\��a�� Y��o�lpZt�f��J=��`������ry�;e�p�*�3Dm9�����>`|�z1��5`�o������v_���2/�r����[�9�vl���/)G�j���jv��9��Nh~_�2eb��&��&�����V��-�u�=�(t����`�ɩ�C�Y�rD^�,�j�{�Zҳ��$C��4Y�8,#��0
l�G�����$���b�L'+:���Qp2��?����0J�����*����p��*�筮}�4Ә7�bH۹��W�10�%�Ο�U�DD5��bӬ������k�$�Ҡiwk�-�Z/�S���vK�X�3ihH��)�w�"��ܧ�_[0��۽�O[�����>����!nR(>{�_�o��	����j��2����ۡ����!�+b��T��|�VY�<���ȾqQNh�d�a$��D�ՙ�!��T�CBut�T����2�M�
r��U�^����琝<h�nXi��(���������FO�N�৵@��o5�MML�QvB\y���_C�}z��sl2o�����AV���ih��t:B#�:'�,6�� X
(�pH�93DH�Ш&�C�����p5��Li#��R\��'|2��޽"�Ӹ6�X�l�Z�뱞0c_�x4���������7�ZP%�q;���-so�9-���Z��w���`�N��4k�ǅ;��"���u8���W�%s���� ��v3q��b��mq�I�9�K�$&;��{,�H�Q�VD�!lꟆ�����]b$V�?A�J��&(���,֯�~��	��em,�ae;��(��e��B���(2��[��#��A�Wp�j�B��z
����玈�߅m�����2���>�=��	ug1�ݻ�*�a���8��MېnX���z��y��1� ���$)������tn�ځ�Ƒ�7fU����	G�'}B�E2���ܝ��$##�^�Ḫ}�o!�v�n��"�s����n=����!�Ӛ�zr��;�E$3�A��s3e��k�{���ӝ��)ȸt���4�MvhqF��,���{
݊� o��6�����0��l��e�q�QŎ}�X3�]ǡto�;�JkF"��*��1��.��d�&U^ٸʩ�yX2����~���J8R{���>���-�1�j�Q	p�r���j��1Ө�[@TV���������^�}���A�u�Ƽ��=Bq��}���3YZH]��f�p#����EU�a#�x>,��nv�e`��r�=u�������F�m�LP�U	Ϙ�O$�X�Q�gN4E�&X���9{�戕N�+ܹ�]��Vj ���( g(�b���lS`��O&95\�hVj3U>�T��r�/M8�k�K��)hϝ����KA����dӤzxv0�z�h�-��0�@:�Q��P�bҍ�J�N!�Z�/���7m�c��c��h�$��!�uZ�_[�A��]�%r92��Ɯ1s�Y�z����?tT�|_��?�+� 1��a   >��"����!�w18p
�`�x�j�h�ȶN��U@[���fRt
�g�q�t�Y	`��A:�t�=�˚�ӟ�{Ѷ@yG�"kHPd�K�|����(Pg�'J]�F���H�r:$�U��U�[�W�_iXU����i��,�ո3�]��|�=s���!�x��٣|����$�b��~71��gL�;5�Y�`���-���[�
�+eX��5;�\��Ҽ�Ej5�<N�Јf?֧���xUP[��l{.���h���D�|vd(��C�vژֵ׆q��k�Y|�Յի�wW�xМ �,�g�,��o���s!�cc'A9���TR�&�u��:�@��1!�Wx@��:�M�`0����\ɻ�y3��&"���*CY��)s٪���+�S����R�����>;��������C�O�Qu�v��������jG|�U,ˉ���|�[Z{s���p8�h�O�84eTs�d��z����'fD@RO�𺡞���)*3��G�G䡉xR�k����s�Ү��̑Y�+�2�nV���J&���ZEr�|�e��`���fDW6�X�!�/��;0J�S�F�	��� �F���7$��,�X�lyq&C���S�����ze�ɞ��)�������������ш�N�<Pʧ�#��=���rS豅�+^o�����@t���m5'~������)��0���(3��	�ܛZ�p�p�Uz���P̳��	�m.Bܣc� C6�K�����Z.�^��C�@�{MI�wa��,�h�|��w�8�v2�0�L,3��W���x�4�>ד��a`x�$�o���a:�r�l����+,ߍ�!"@��ԛh1ڧ:�V�I�n�ѥ^:�c���4��	�,���v&�c1��gM�C�8��o�J,x?3PF�-�M�"�̎:�H�Ѓkj\�H)�����jb�2�Y�~�����CN��@���"��JF��4��: �N��Jm\�V-�/|���Ü�[��m�m��^!�W�)i�|3[q��f��~>�RQ���fv�����4��
Qh{0���:�2,�4�C$�t�f�R'f�8��wo�Ie���!�h��N���r��w<z��f2	#�-�!�ӫ�8��R�����`>���E��,�����1a�n=�+��z?�9�i6�XA��v��±�3�<��;�rZճuJ�D��V4��?���]�m�T�u�@\`�d�%]�H�a1>��<H��A)"��_-C$�P�'���.�Q���Bd���!��K��,��	 ;;�Z�*���Y������N7ʳݔ�åY��C���4��yy
�$���?}�r�+�ϝ�&��ѵ��Kp묙;�K����y�r��ɕ�?�o�����=�S�A�o�e��0XJ�HA�Riտ`��T��q���l"���<h�����x��x��}Lu�$�T��݋��|��T�'�
��K�i�-`�ac�����gh~���a�L^�]@������|g&p���frg&k�m�@�vuښ��^�]��9�1��ːe��xK��Pڎ)��
j86t�����RL��eZ �
���qaܳ�W�M��w�h�\;k����Q�-4���-���V��(��(v���5H���؈��<�&�z�7lSSH4*i�D雤?��#v���g�L��?�q��:��00 =4��E;�$t{�ݭ�^��U��Bmjh�xoat�0r�@E��ó���4~h�w�4iEo�S�����07�S��ǟD�,�7�7N;InZ�{�*�QxB&��RB�)�yٯ.b�.۳����K<����6�Bôu�neV���"5��+��fC�n�x�̒-4c���jU�����W�~(��{Jm~c5� P�U��曇��d�1��7�4�i��BVtUjo<:��	�	5_��U9��Њ�;�iu�[���w>��Ǝ�a�E�G��7٭#�~R����RC	T&�;��6��ąKI�K%TP��sԤ�h}ۻt\���{��I_��v)�]��m��[�R�|���0�O���MÍ�%��\Vm@״� .��&�/�W�mǹ)��W�T�}�Mӈ�\Ԧm�D�t3�K��B���5b�����~m�2�X7�