��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��˲�|U�eu2���P�1����J�2�@y=܆��X�n��t���+-1#Հ�B�H�b�~"�{����;GH��Y9�QR��c��ׯ�b�i�j��Ñ"(Y y�AG��) lW;#��2��rn n�c��n����dӻ��4q���狙e};�e�h����ήr���[�̉���Y~
�-�ʙ�d`�d�Y��8���N����j�B��M��tI na��#B�`��f�v����+�~X�<�V���~�����p��ӕ�i�:[�<!n$
������˰?��<R�$fjA!*�,�gH�ihRxpBLJ��w�kS�n'�����fcCjD��͹��[��,[SuZ &苒����1_���1�Kx����tb0�PP�������9�{l� 2��@��ZTS6Ӣ�(*L�ě���cr�3T�- It��j�f-f�!W!}5�?T}2�<���`��?!�"ُ|��I��a
>q�Z��y��K�����f�Ϝۣ2���Vg�+�UK4�)(Z�����a59�l�����lˊ�g�VP\/^~�7�W���֙�PMD���D�B�WL��km;1���K5���#�n���W�i�#0���Ӊ�Q/Jd���:IYl�r�P�*i̦֦���ry'��ϪZ�1�ǃ�j>xW
���	����_�w������ԟ�ќW��~Lf柟5�XaU�f���^�SƸ��].L8�.9o/�A�7���W�E�����Ԕ�@��<�{��
$nZ���O��EN��˓�={�=��D�"��}s&7��l���W�Y��Zd��g��鼦8�`9��~'�����ۊ�p\ma�Y�����7��Em��&�E��[��MV1ؙ�z���4����Z*�uƱ�e\��l�{cc���yЈ�Nj�F�b*�?�:X5uY���A��c8X�3Q���Nꟷ,���4�6c��8/��n�7S��M�ߗ[���C�s���0��8�}�e�춳��uwp��|�Gc�x_bx^z��NB��������Z6&�S=x�wׂYAU"��V�<:܈�C(��$�
e����Lؗ��]�C	w�yD��R�+�g��/g�Z�~a|������@�<�)������[��$L�oy�r��y�dDb�-�kTE���E�fK���k��V��iӣ��}%Ut��1?z�ϳ��DP4�1=e��NGp�����$g�P����c���q4#�/�[�����5T���%c�;�/vY�ɱh+�Q~=��(��j���킈<�I߁i���W��t�����);�����էl��"���Etq���GV�}t�7GKJr'+�2�I7*L�/�e�D݂�Ȣ�����*{�@���>g&��
����}��Ļp�z� �r&j���`�/V��*�$i����:�p"�y,���C��EJ�ޙ����gIy^��jɪ�Omg�wD��������"����O�GB��+�o`��WF�%�f��:���JZ��g!U(jkmf�2WN���w.bAN^!���5;R�E���R�Sl�g>���O�0T<�^7�'�'u�Nںmy���4��dW$��s�]��f���覇���1Tgli�+ �y�5`m���Q<��ތ+�/��h�Ƨ9�h�t�����9�i���{�Vr�h_��ŭ�}>�5Kʸ�������4h�sC�I�"ݠʢPQI�Ї�5���'�_��L+
/�Ig�2�@s^F��J���#�+�%��ݷ޴�{_F���N����h� �;௉#y�ُw�|�dU�CА�%�[��.	�Z(�I��~iPh�0�r9pgI�Xi̽��%|���$�~��v��s�%P]���z��	+��8m�r���^��tB-i�����N�.�ܱ��>m_J��sk��Xm'�{��0%.�Y�[�vTE�d7�m��R������.��N�^�rD��>��ٱ���3[�čNnX��Q���Z�$�T���J�k�wMщd���� kQJi���W�O��aR�GlFMd�ʧӊ��Ō���`�6�[U(�N?M "̙�.��ƚ~~��ź.A��F��S$Нs��o��Z�)k'�y��sl��n P3��ަz�,+ntB��\8��`~��,�TL�t��Ixޕ�7�a�N�>���� �Ԝ�M6�>�2b]�?�7�W���ZӺ����kf3|^�Ť[J���֮2lc�S/*�s��"��c�1O0D�ޝ0w�Gos��e����ݤn �d6�Q�+se��V(��ch�h�6L4XG����S�GYxt����(�TzH���iM��<�^���2�r�U
�|���q3�]�v�-�nM��0_���(���~,Y�C�.��Q#}��4�D�/�ݖ�ݥ�����Qq�f=\Ί]8��E�Ӫ%e���Ae��9���aT�~3���զ��	�M��D��hm�N�m�'���4�C:{H��s���FN�,�B���=��T8/3jRq܇m�ۭ�%נs�	�!��i*u�7Gr0N#7�u�l�;�)�!�]{��wi�ֱ�tW&�|���4Ǡh��S)�D��wa�W @�MLHY�k���S����g����iO�m(Ͽ��c�xƜ��wYad>��W*�/	��K�>5[�����59�
+�M�7r�^$�΂�#�����2�Ty,������N����0΢&�az�:�HEZ'�S�-���ݫ~�������5<8j���^s@���Ԍ�k0�P����>���I*h�&��nu����3��6�&Ia`_A��zj�n�/5��b:�!������kr�8$ƯJ�a��5��hqo�`�W�[��c����̟�~���A�T4N_>֑����AL����F�� ��M/��'�m�6
�rܹ��l�A��eOZ��Ȕ�ϓ��o���a���<w?!+�)�,m2E޲>�ˢx��m�9֗N�pܵ����?h���8G��^�����e�'G�/6�{�ڿ�py?0�� ��R��5C�]�G:�Y:2J|��JX�����訧[Պ��9L���� *;��k#hN���Y�7�-x�o"'=��iZ� �Zdq���Re���/��qh�e������Y>�A����>h�-�r�I�#�t�¦\�)����2�Sap�^|bm�I���]���AGRqZ��PW�oa�Q���Ca�K��A�HGէ��J���*�_I[5��T�38KrC��܋�g�,�й
q�'�XnR�2�a��0z�&���Vf�5N6�t���`����5�c�
���ierj�Y)a�����f�!6I�W�%r��X�t��v/Es�.�^�ޫͮ$�� %��-Ҳ��6�K#L9��g[(�4#u�V�$����@Ҕ��:*�:QPL������ŷ�h;F�$�C�������tR�m��5��>!L�qJ߫D�pql�-l+�������Aއ�z��e}�	��s�?�º<��d���E���?��|�z<&+�]�IOȥ�c��
�1`�zr0�9������n�o��d+���%�^�A��0�� �����|��d�p"'%�G-b�͡��JVzm��:lA!�P�uB����a[�q9��7��&�ϥyg1��;2ӓ��������Ֆ�W
`� =o���P�y�T��9q�u��+�&���J�֡�3�gfLD�x?��to�h�ZG珄����w%R�V#W��AFn�<�A99���D�=@_ VaҔ��R�J��������o�>!�46�����d@��J�J�;�<��d�{���[)+� �Yj4NY3I�@� �/��tA����s�6�|�3s.e��Ͳ�;K5�:�G�_(�s�y�<�Yg&)���dM�thZ*}�/���<%
���"T���hR3�E<�j(<�"�!!�Y�z��Ж藺�4�Be������ši��`��7Ip�;����~��c����O ��x��,�`�DAB�ExBޅ�ኄ=4�A�4=��M�������{R5a�aRԭ|�̊�:������24Qɍ�4ȌzN���n�z�lw#�pf��U��@�Ȏ@�K���Rn\T/��X1�ǓvCgY�t�2
*�������֫�� ��0��@ß��p�ko����a����g�= 6���	m$f�JJ��9����֢�+�F�i9�O�&(�.��g�k�����hgY�j����(I�a*7�I���X,�n��W��u3=S�Uct��&���7��.CX��6^L��ι$�v��ը��Iܳ'b��k��яB72ֲ�0~��H��${�g��'30�<������&	=�d�H�x��!�/�2��Df�c�/�Bk���d��WD憍�
�s
,iښ�U���xi_Xk0rO�IR��N�#���s���nq��1��ZY3e��&�6��J�\��J�O���	r*A�4lb����]r2��,cc��X�8oᛆ��/Ҝ�/��X��˝��u�O�BC|f<�퀤 	"y�t��EW�3/��#���Eٛ_xoO^\��7���b8Q�^8���ߏ���cx%Nos�\�Eh{K=����*嫝���9���0���֎����&�(�p��aQh�b��!�H��Hk��۩G^�mB��1KL���?�:���k����帾1���/��(�	��>Ǔ\Lyd�!��/�g>�k1�b%j���=T�v�C�W��i��$>���C70��V�,$+*S�p�ɢ� ;S�d�$f��Y�b����Tc
Zi����KKr�7" &V�K�GaÃq�kޓ7��_��[(v�mi<����glp���U��3<D�A�S��a���}��� �s��"n[���������E�c��C�!�'�M�,2\P�[|������-��0Y��w��PM:��F�ᴶ	��M��u��@z-����{��L�����ЭV+ÑE�Y�^*)X����N�XU�~�XC?H�-�c�<
���B���C�g3����X5mP�l)�7�r����3�>��w��d�J�=֤Iƃ�p5 �e���:��0�i��1{�\��Lǜ3q6-�V���4�������cĈsA�Z�O��OW�qG阽�R�t�I8�F�ȇ���[��&?A�zv���5)�e�	��p�	=��)fh�G�WQ�m�+��EJ�n��vC#د��	/�_���O����4���4&d3�t��X�d�Y^ʅ)Nv�J���� y��-���&]cm� ]�`���<�_����f���N#�s�̂���j���E��L�7��y@vo�h�l�&���a����~A^{p='E���z��$�8�`V6�AOƵ� �^~��u1Rϯ�lP%�3Kl�;Y74w��B�:��;�ƴ��s��ke�AVg���!��+J&����3�7*�t8����j��ɿ#~a]+�,�g#]��3<NY���L*�|�W��k`��Yk�� ��^����-^���y�f���4n�.+�Hcv�|��ò�t�x/g�g�^�ry��`���tw	���Ǩ�������6�O�:+�H��B5�G#�5�b�i�t68��U�\I��y�W������
Hi�)#B~Ӻ�Ys>�(�uu��� �B�wW���Ζ����
/�l!��_��A�6������X�U��VE�fN�
�l�ua=i�qU�V�;��t*fO����`'���C>d����4@�Rn�;1�b��e�?�.�IG�2��}-#�&+������I�?=����5	��I�~)��UjRIoPT��>�ѻ'nI��|�C�Qq��nz���hі���o�l���'%=A��bɛ-�m�@cQ?1M:�G3.-2Vq���7�&���5��H�%��flRv��(p�z�2w���$"V++U�_ (�Sș��4�����C��6å�Üʫ�w�����$�Ɛlx��55�h�֖���#�+�qHe=�ƞ���2фU7Mxn�4�+j�C�*�Y�!�?T
L˺9��`�Mb����ˠ�F\G��İ��zA�G(�0��/�������gc| ;�^�,����b�XV��wM�idtG��gF���wJ:�:{
:�*����2��{�	.wDU�P�6$�{�p\b?��t�i6���1�|(��ȩ�܍S^�==c�eR�wR��rJS�8,HT�$Lw"<�Q��+�5�>B;J��ߛ�����@�ry�`�8l58�F����F��O��v�~6;
�a�{AP|e�6�pM\ X}s�co0�[u;,�W���@ _��=�}�����׼hL&��}$:��eڜM%]q�d3�A|�8���@C�0p����ґ��"pq�Z������<�j���z�;��޴<��$1Ҳ�*�Z@0����k�+_7�}��7��;.���$��4i�C�4��i2�q��^MU'��0sc!��~��׌�/M����s�F�$��#7H���7�r"kS������!��#�Nv{9tt��H�`�%�F%��s��w�ۯؚC����lR�8Itr�M�OMz!�-� �B�A(�@����b�pZ��?��V�����;߃�5�S�)��1pb��Zd#��w�E,��N�D!Vy2��,dd�J ��Z5\�D�B���Ny+�� *���>�_�z#ҙ�T�g�0L����<�m����D:�	{0�n�k�_O9	�"9$P�w�8P�@�u�K"_ҟ�vn��(�X=1rː~wy�Kq�eg5o��� �ǜ�
�����"��v��Pf2\5���$4���?�
\fV���<r�ڳ��s���@�ȱCь*���,�֜��6Q���α1|���Wp�$�H���ӥ�/�h汏�Jr"��%�!�!3p,E��xa��|��H޲N����>�X���p�⼾�@|���SA��ƚ�@
`�t��������x~#�O�ޒ�	��n�c��}}�4K��i|��[�)r�YXa�#Zf�P�JPIM��S�w��x�����u�{2ߒ��N[V������[ �NiI�r60�|�(�\Zp� K6�k�N�E��Sv�tB��~���[�ˆJh��m��y �+5��I܎K��G��\����Z�вr���M��+/T���v��Ԁ^K�*�ȟ��~���4ߏ����S��ϵ�
sC��;�H1��j�G��s�����4&�:e�0��)M�n఍��Z�����9��&��}�V��f-�)���}�
u��3
*�Kl�0�cwl9k�QT���*�zC��r��,���2���4ЫI�f��ȑzo���n��ٌ�J���b�ʺ��,B����X��7{ �����w��f� ��sd5	9���w9�j����r��p-⨱]{��{�pxP�Te�n�v���R��V �(��ͫ��0��J�8��8�`�{��H�c7�WB��I�8ܹ�y��Sd%�D��x=*TiM��X���^�ȱY͢H�ϩC�k�dM^/��k�������n�c�-�zMԇ��a�;�@�"6�����%���KvS��NAʛ	��xQ�`o��BԨƏ �6�W4/��|.,֦�n�$�5���?�}5/'}�
�n8�N,��քcn��7�<v��ٻ���э��-�����Ѝ� F����n��&q�4|u���g�k�����\����MO�)�sM�]Ny��7��b9��r��������g�e��S�?�"��x�o�>�5�a꜇Oye�����ߐ�s��h�Ӵwc�l��kʼe�U������'�l�g*0�aKH�N��.��S���Zw>_Ǿ����[Ūl�r�T�˧��UĴ3���|�Y��(��!H9xi�'5)��^KԶ��#g�-�D�&�E-6�߮�᠚�+#F�w�o�e�ت
���8��"_38M�CD!�����c�2�~�>d�XhmK����j�;
_��9��)b��W��]��EMj�p�A�����#Z�.�
��_cǆg�M���#R�A�˒�-�?��Q{,j����f�!��h�uk���8E�+b��t���tS�(T�UFJly��x��^-�)��q>�t��0�������a��e��1��SJ}̢��dUI^�"i}�}�<F��T���` ���L1�}����'� Ohi�Ec�A=1�~�%#GA͡N�&���^�Ht�*u��, 2�گ�
�m�1��x����	�?\ ��32�x8thV=�K��r9\y>L���)����SA9Ł���g��͛Z
W�'��ʺ�O���3���K�Vǒ���y�-&ҟ�W��Buv��eb2!���i��gC��n�d#Z0e�\JF����j=J3Q�>C)�s��Ų�\������.t�2��Z�L��{m�+�\�
W5�y�"�<���p��N��S�������D���}ӿ]��[oH��5���,\��@1��|�����$5�3���8�X��/���2p�+٤�"0Yj���7����<u����i���0�K.��L��^mg�B���Z�9?,���5�
hk
;����[���E�Z�f�I�x�l��;V��DS�a9�R�׵�ΰ�o4�&Z����R� ^��v�K�qdhm�xn�|�C�so�S���O'����pN�cZ)P��Ѫ�Cw��H��y�C(^�z���t�m��g��^žF�d��q(������+"���K�H/(�=�=�g�}��XE�Q��a�لl�W�'���9d���!KB��~�7uܑmՐi=P�^z��@y`�D�S��'/x7���\�Υ��&�I �Rm|���8�&�����<��N�(��_�R�E5�$WP��B�����4�޳��̿3��]A�WP���'|���OaC!�r�'T�M��=����)�.^�<�0�&�dޛ��dsx���쎄6�=a�z�j����j+�p�#ᚋQo\8�:��E��a����ٝ�&@�}�D���E�����X�������E3(���(s�r�r�W��$�:{u �ox�\��6g]$�d�T[�[��	xp+�0�k��74�l~�`��-J�	�@�3\�0n�^�T���-2v(�A����92�f�fZ��.�О@�������etl��ګ�$:����2�������˞2�>Lz�&��O��ݰ�0�'"��8�=��>������	�����[�S���J%�N��	X�c�������#���%nOj��7�w�d�RN���O��S���&���n�@}���(u��(I��0	�-�G�s��聂�=�E��!�낞��#*��K�WՅy3�+��!Q7B�vS�PM��f�/�w,%�R:�m�?��TG�r�l����7�*ZZ?��KC4(kͦ��h2���[�>[;3��*�g�@3�7�>�)�#�l*��A����{ԝ��J˶g��Љ\�-,��<?�N\�-ݪ<B�XE����Y�Y!��#���r�)� ;��ߨ����;��Ƀ�}Ծj��!���0Va�8l���G#�2�p4.�(��fJ��Xま�2^���;���f2�`�>�B)���V �����|hf_?��k�T�+Q�s�i��zP�H���N���끕9�xNt�ѓ�ɷ�[��O��znB�
�23����AP���Z�0�fs�j<�4�?Dd�s�?$)���{z�u�I��I܃`yޕ�w��2�6�UQ%~=�#cgh~qh%aƃR��M����{�3��LO��X�4��LV�k�����L](�HO�ԣu�#�vB��o���nU-.g_2�)b
�LH����/ap����X�[/ ���r@��q%��Z%H;���8��5�C�9y[�����~7�F��o� �l��/l|�����|��f�c�b�G�#�_Yf���	�\��وw�6r����L!�7#gM��jG�7o���:�+��w�m�<��������6���l	ަj�-�EW��кl���f���J�f4��`��!㨋��cE���佮+b�����"a"|��*�u�ك��B�����PzP�ϺJ91V������~�c���(;-�����2S
 ��+_"g��9���J�����5hCQ%�� v�L��h/ I_	Vs�>m=:�˘��e�Ӧ��H!1���`�H(�!�M�}���l�S6l���Ă��YlI�U��A.o\��H���\؆�vTl�\����N<<��[��~��pd��l�,l�G�}.��=��CI��X~\���>ҳ�����;9d�T��Ry���n/Ty�V�Ʃ���S����v��TMǊ3�|���U��Rs,�iRq�k�x���gJ�؏Z�4P[�K5Y�r�����U��+$l2�H�H☬�o�oI<�5�`���M��E�#�v��yӆ�J���Q�;q;�!/���Zj��3��+��h��;���_�c7U\��9�� �������v8��	;I�&H{A�����6x�O��x�ѯ�a�����'�o�0��~�B�U��c#H�6�		���|��Fqq�(nx,n�|�~�V����9+4���pNP}7�щH�m�f�] rO#�%�77�o9��)����G2�9�ɑ'��(�'��#�V�<�eq�u7 4��Bog���KC�1��k�P"P�J�9��hRL]����֞`��x?�����q���aFut�����K�#�Zܞ�p~"�[�+ɖ󽰢���+�T=#.� �s�ۏ[]�����,64�!��\a��S�<�rTq��>R1<��'tԎ㜮�fϺ2.H�X�X2��.��8�-��ݷ�*��paN��~���C�?$����r�m�M���V0�}�'�հ����c*�7����Q&��^�2��g��Kg�
�|����<3�#ށ�D��mo�E�p��ܼ]����p�9s��/�1;Kt�׺��q��9F��K�����S�n�R�n��N�p��g����l����t�[�t��J���;,ՕJ�*��mu:�L�;v�BCE��?�^���k���Pz��5	��x���B�nўOA7�MK����M��륤e1�qU�����ε�W<� ��>F�.��=�g��!��S"�vq{Kn�z�Sq�,�5�W��mbzV�y!45Y��	}'@�&$���p��1���c�:�uBk����&�r���O��x�r� ��,&{Å�i��<����R�Ԡ�� �o'��nW���lCJ�:VB&�L�tùsH�xu�0&��@�{X;ax���8��o !z���J������O��2�AlN�H�QK�NI������.��oIr�;��d|
�w���
a� �B�ux�jI�/Y(vm��
5Fr��;% L���ΥJ��vEtl��[�a�Mt��n�ڵ��j�/�f]��j��k/^�r`���FL��l�p����)�*�UV�9v*�p�	��;L�̂a���UH+
��H���E�nܧ�/�f
R��e���^g?ue��]��8)��KP4��j�y�YS<���jg�gQ��a 3C1]����B����~��O����i�����[���2���G����grq�8� �G�b^]�j -�9`O�	)���Ȓ����i���a��[&����ң�*���e"e|^�(j1��?������#\kFCr��bB���N���i�_g�`�	�m��.}lh;���,�&�
��S�d�+�R�`�=����W'&�̮��u�Z�"�Xv���lv`ģ"G����#$�����tz\'hI����_���B��|�yb�޾���^q ˝�:�*c��=>��|�-+�徨��}��l�*��0�	���%i�L�FYF��F�c̣����l���E��V�z3}��jv��u����aP�_�m��q8����o��\�f���
��h�ͯ_�;��i=��q�P��`#��q�����n?5� _9��~�y�E��+�k�C�X����cjk�+��u�*�=����&أ䔕���x)��E"�x��->���*���Rh���Yy3��>��=E��>Q�(��T��Ĩ�t:�G���Ra��\T��k�-��8Rw����9u.RL�(��l�����<@�)����Xy�QC��֏�	��,Y��F����{��F��W[ħp�-�1:��t�$צ^�S�C� �w���e2X7��cO��o�ǖ��vQf\}��(	����Y�u]��Tcl�Q�*��l�{�U��Iqs�yn;�K�O^�t���Y6n�F�<Xu'�^Q^4[�����������9�Q��f@Һ.Jގ�����R�80��/[��n�)p����ԶPb��Q`�by�:���	P��d�����8��p3v#�a�B���|�bn`l?F �ڞ��Q`m��@D,y;n}�/Ƞ�e�ae��k̡��O�\�d�\�1���z��D�T�~⛆Hl���8�u/]�0:ʢ�jT�)��Rv�s$���<d����K��r*b$`ul�,� �)
%�E�vyY|wp
[C�:0k�$&eH�r���i���vRa�UZ�i	:�zc�IQp,ԃ.p�"���66�Նe��]��s���U� C�-E���_�I�����,0��s��`X��~\0�xm�������A�����?���p�z�R��tz1ۗ[8����R�I!@jZ��ʴ[�|��7���\1ٕ���4%<���Oc�Fr���]�!:�����TY����"�՗�"�Z�����~�Y�q�)"ğ�����B���G�8��u��[��C�4�ԙ)�����J��y���fE٢�]\n^�fng�֘$�vL&(ܵ��8FZe.Dftg���mޥ��>Tr�3WxZ�J�?��m�d�^g񶜜� ��%�e�APѳ��C����u:�i��+q�����?w�B�SL�-��-ٵ��u?�F���<��7@L�J�9s:���Zc�>��x���k�=�|8�`����"��{9��H�v���a�1
(�ʈ5�a(�$b}=��� bKie�#=�+?�8�"�?���Ș��O��E�a�8M'ވy�\i�	�@w5jEXޕX�.�-Df�v����׆��$�:�p�]�WX�\!N]D���%��*}���,�p{�q`V��҈g[�Fb�S��j���Y��|�Ϡj
�PB*:s2'K�1����>����QXn1��ڦ
7R��%�r�}��h�j��?��.f��[o@�a��;1�o�!�	�L��䝊�.Y�����A �����sջQ�%s��%(���^��%��/*�Ls��+M͏�������b��HV�a�����V���9N��x�5���Rzr�T� �Cǩ�D����o�Fe��\��c�{($�i��R��l�6�>W�yLvb�!�9q�?iIj,�#���ӥ���%��CR Q����j8z"�bc��c�� �	.GL�ֆT���,�}�vm:m�����RGV�G|&�|xm]#����P�j#\��Rc���q���bs����G£z]7���9+���n��6s2|�y< (���Cn����90��[V����ɫ������LPmm��< �8�����)��9��n��Y��$����d���-�u -9ԥ�~�Ҭ�e���u��`�GPHJ	4��N x�a+B�����R����g��'@��Yk���G�z�61C'o:�	��~��҉��_�:;"хQjh�Tl�o�;<���*��%�f��"vt�+o��T�u{t�޸ӹ[�k��_��uk�����_��U�U�/%x�y�;��˳X��E�z�:�s�4OҘ^S�{��Ԓ�#g�S�{��C)s_r�Z	�>�Er���b��_��PU������l{�vR�{�<¶'*^�ˈ�+���EQ�k�n��VxQSVo�+�g��O���F���{P���X>���d���2Q"�G�F��z�sǖ��"���	����L�S���Q����+"R��9=šY ��E]���$Ւ�("$M�'VK�J�D�B�.<����@|�=٠A�t��6�$])��~zW+�q@i&�%�J?��5��	�;;6��Hm��۫X~5�Н	�U`#�؝�7��0J�ރ~��E;L3�y2�_�O&����%���������8�B�>����{��|��6��d���Ǜ���_�ڀjn��H����ũ� ͝��v.��J�_���
��l��Ց;����mu"H���zf�ا��C���<��I�~ʄ�nF���M�xX��W�>{�t�*7��x,�
���@|m'��̇&i$]���x�j�^�ٗ6M��P�(�̓����R.�<!������l�� �r{9	���*EYD��"rHTC��,�l�݂VZ��]c���ZH�J�Q	�#lQ?+�1��)yX�Q�_9��s�$��yVL��6��}���[���#�6_jQv�PV��Ѱ��C!y���2�2��`�=��M�d�7�����D�����1.��ܑ9"���%+�*c<�)�ԏ6�j+���q�B��Ŭ��Z���9��4k�Aؿ#�^��l`*wU�&AQ�禋�E٨nιA�7.r呂{�9��(���
��U���Y�lf��X�Oqǎ���{��~R�ā�\�����cCpϳ�]םr��q6��"yߓ��ܘ���;x�]��h�{oG��P�4E	#g|^+'�vA�CI��qXC_��@��QE�ŝc$����&���Y��C�_���uSH�D��;Aa(R������9T�^�3g�������{���h�|yy�)�z$x�<�3O�����K����Ti�@�(am5]�] F�d.��bp��@�9G|'��8���2�������UAiQk�Ç�U���Ft05FGk�%�s�(,�,�s�1�=�m�F�J��0��1н����:�7��s�����~md���1UY>���,�z�*Q_i�!y���ݻ�q��"|C��ޯm���?y�"?Ma�΅o���� N��Y��0��^��N-;�x�섟Y��[ǭ�g�m��H��o|c��E�P�T=j���e`?��J�p+�)g��VX��ǜ @�����/�VX���|4Um�|>38p:�L��؁���o�.���P���9��nx�V�oc�
1�O���]h,p������$Ps�*p6F���$=�A��S��U��b���ph!��~��ӂ'�X����C�PH�]^��������Ȳr<~r��=f����C�>ַK3*i'~����o3u���*[:o+=�g�-R�o���I\j!E�{�Lk������%;�o�@�K�a �F�X6n�=�(~���F���_}EQ����c��s*�#�T�}��)K��	Y�k~�5]����Ͷ���Bȡ~�m?N���Fg����a�Y����@��]�T�;ם�0PM�Re� �����"W�g����lᶩ5�sE��:�œyV�����R\�o��F������(y;������?�m����e;Ѕ#�SR9[h�ɿ���Z���UdĴȟ�ZhF��h7�.tVA�[tU���F�{ϫ�h��ٜ���>Ҵ�۝���m��.�"�?s<�Dd���#E�ȇ�����޼w����R�# �X�a���K)NBYEÏ���*S	�ҡ����ե��B�0�Ftه�D6��X��ˉ�<i	$e$�\�߅�:fŚ��5�8�YDyk?�Ժ�)��Z|�L������<���
���3�N�ު�*��c�������r�Ʉ�/��"���	S
�4f�,h �\�Fa��-Y�2���_a��=��ژLЩ�B\{��ު�����'��4U�ITu����m����>�g'�>%�@]�ˎ�<�Ňf��<���TlQu�!b��)	���F]��'�1���|�FV�<ʗ7M�T����ϣJ�̐71?R���^N.��	��Ф$$��v��D��tߴ�4�Ys ���l�A�$+�(ː������]8�dX	}[9�`:�v����B�vQ>�h�~-������A��L2%��4�{��b���`� �w�*�T�Q-_g��.s֞��J����."iO�}�_�Fŀ`�+��ǔ �B��Mv�oz�e�"յ/�'t��;�L,��SP��
�n���J����� �%*#k`[/�y���.��"p���o>��kEA@��p��<^�*i.[M4m�E�f��l�([;1[)l(	$Q��.��C�&u��#'��z������I�&Y���A$�����ّ���0[�ǂ�!��+uI���zb��w�R�ǳٷ�J�c1�jG����ۊ&���ߍ�R�B�w`y#8���v�:gwQkoe���L� �Z��k����x\1Y>9�F�ˢ9�(�O��I�u�~�x���T5�X�^�i�e�4�(bӛ���'-���i$9��}�Z����SPO�찁�n���=�i�/dLQ[��k���`V��ڵ?T�R��Vdd^o�A	��V�� ^= &_��F�u8ahm������¦�H���Tc�.�RxP˗� ����c`��h��&����a�pU���.Q�PQ��w�+�}�������|8�i<dH��g`ZX̆�g�JE{D�H;�_�󄛒Y��'�w�����7��h1�M����Rfy6�g��H��en���a�;�p����~�ŶO��X���w`{6�oT���jgc�
d���ܦ����a$B����>�H�ر�7��ܽ>��H2�!{H4B�C���	i--�(X]�%�Х-d���'�H5���_Pd�5l�j�a����.S����C
Ie�A�ٴL�*��|9k���\���
I�#���0	F�Dd�	H
|��k>��1�6�?����ˣk=d$��� �������/�9/]{�����/FeiD����"g,B�μ(��t>$Æԡr%���#Ŀ�uP�T��޺{=�͞3~s!8�0!�%f������{d�VwaD����Zݒ�r�m�����U��Pd�{.��U�_x�$"�h��r�h����&����b��a�Y��x��(��'!=F��~�P�8!�3�\�Pwl� ?>]�Haҕ��.�ˈ��D|���C!|�O3��_�%h��q�6rg�xQ妇�h�u ��ʏ��a�~�~=F��ğ�:lOr��X��V�^]�ޜ��6m���p����,�S�1Sb���כB�Q�$+���7��w�E�jf����;rw�\��ܝ>_�Kc�Њb��v$J6z����w��Y���<������5�ۏ�C]�;�`V*�Y�ۻ��%�_V"d�g��MϘ]x^�M8,��H���W߭���Ǐ��	1/:�¢�-Q ����HwК8����lw�(,e=Uib��*�D�m���Z�bj�9H�� ����G��^�޲ ���x6WCO��y$�k�|�Ŧ���!��4���(J�qzY-�B��w���-sV��gx:_l��
� ��n�����|���B{�l����;Yaܼǫt�p"��c��a�H�L�-t���.�=۪s����`�ɨ�eN5�o�<o�
�G�sa��k�����լ]U��~�G�I�&Y�'ֿŮ�_C5�A�&2����m�����?p+�:Ō������,ŵ���K�{ۺP��H���%ۚ�}��V�߳Z��3W �J�zޅ���k��s;�t+�ཤ�c��I����| ��o������@ZY��4�9�l��k��ӻ�jYT14Iؗ�J��7}�B%���v,ǁPʈa���T\��}���E:(!M�����ղ���o��^k�����_$)1���wس2Z���=��
��BCত�����O�5mi�bM_�LI88�k�������jk�hޅ���)�繽�@nY�л-����8Y�K�����ᇴ7�{���dD�x����l<>ŎԱ��e�qj0%b�AB}A��nrĔ�mm��~3��C�\L���;YU�j�K���,��ו��n��!p�8����|d ���/nd?<��ٖ*������լ�� 
�A�8n��E�����ƃ�7-/aB.�\Twkba�Y�$HF���Ȭ�M`�{9�"ZIs��WN��S�ƹ��>F�i��]��!������̢������,��ޱ�
T�wZ �Cϥ�:`�52�|<����o�Xt^T�#R�K�u#��{���r�W
dQJ#��!U5��V|�Y��Io�^��;Ξ.n;yT��.	��ה��_�s��$�O� �2m2ܘ�7Y���e�I^'wN�MC���Bn�g��J�p�vr=����p֩�ȭK�s�ι���aY'�ʈX����7����B�Ż�)}Q� �]\�h��J
%0� �?l�ź��������S��l/���
[��>�K{k��?�3��nb8<�4ug�)�Ie��Gq�Wz�8ĕO���d���%�V�H��彲��#=+@��ę�厶�,��t�v�}�8�ϕ�3Cd�[�I�g��Nk��CvL������dVZ�S�k<����Y�̆J.��?��S�X7�O�<�Y{K�\_����k�.�]�5�;M�MѫU��
,dl�o�Z��,�`���ū�Ϊb�Q��CHGG�P"�T|��u�+���������l�h_��aS�b�Ņ��!�;�]�S����k���<jXU{"NFxk����CrZe5_�1���Xbn~��1��l[lt��0T��0g�V$w\ib�7� �K/�S��C�'<������ڂ֙�&�ȱ�9��E8��-�B�XM��Omtw7���x��>�"3R�F�8Z'�~规3/&��\���4SR>�I�T@U�A]�gv�w�_�3�֎��w�T��� �N˭�fr_&�9���>Z��~N����0_C{ �k�����ᗽ(&�<��W��R9��r'�3^Ϡ?�R�:O~fk���u��跎ʉ��D.���So��ܒ�R62����/�{ҡ��8kfv;(j��M��