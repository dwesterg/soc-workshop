��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E��KU87�שsLF(�y�Ơ�m[��ܐ�Ċ��4�� l�h�q�.�w����3`���� ��P�ɊZ�L�jY<�2zY&�!2C݀�b��U���cpA�p&�|�M�b�_*��d�D���OT�*j#��]��g��n5�����)���)������D�i8_���gaz1~4�jUx���4�HɈR=.�R�<O���O g#NUW�=$V�D�^�c$C�z"[�l����Db�k,K���d#�z+8�W<�/��bQ�^��A��`��aUU������~�Ka�n��Ap������q��]	����H\��d��[��^��=�̥��aCD4\hFn;vlA�������VS���H�-�'k e����g�TPy	U��#��I��U�~Ee������"h0C���&�RI�AJ�PѶ&�@�O��n 1�<�٦_Ѽ��D�������ة���n�IV�;�[*�A])�A��M;�Y���nA)3gL.HS�e��3;��S9�3jOA#���y��7�݁����!c �/
O����@���	��`�����m�;o�(ћ�bd�d���X~H<��7& ݢY˒��} dA��΍9�>���0<9z�L��� �U$���B��F�&�t)���E�xUk��e�
^���u��K2���3*�B�$.'� x�ӚI�� R�X�-6j�j5 �=#ἀ����P�Q���	^�zC*���z����@� ���c3����Ɣ�<^ �+`7մU�0���o��{�p��Z0(@=iU k�^��"�o��Z�P�Ă�w9����?7JA�y��Xm�D��'MkY�˧N� ���=4�M�?�F��C��_�u���p����0�W�M"m6縠BEH�7��t���~+g��p���F�l/n��y�<�8�$���̋� ���d�.��7S�p睨p�+��0N	H@fx�ڄk2��"������+%P8K<&N�A��OD�&�ң��F�S+{��F�省��w���~�6�v%<z ���(9�}ڝp��`��k�������7���a�[|�$GbQ��}U��F��JNٹ�ϝ���mq����E�{y��O�ԏg�	v���Jc���E�L�`9@�f������H��n�	�sڠ�l@�&/��7��eHg@53W��BRF	��p�PZyF(��K����6P�GŸR:�������4�êx+.����P�S��3Q�ڦ8 �\�5Qdg�9:���o#�'P�d"��P��2Є�1�V^mU��1�dI$!8���
ڠjmB��N]�¾�d������ϼ��4�u�kh#0h>���,S�&� ��c��8wc:":̕+���H�<��[�y��COC�liӕ��{���L�����X3�_���T��|�P�P<τ�	Ĕ㒪WgJ�!Ng�ud>4�8����/��᝶o���ʺ,t� �t��^O�K����(1'�f���N>ᗨ	v���.I
_<�i�8�IB����H����xH�f	�q�+S���gI'T��\]2D�EI;ʇ�����o��S���)�"�T"�W��%��6�~U1��^�&�i?��O^�3-ج���LA:]�+�8Gtݿ�6�M]��g`��ď���W�)rv��{�)��Ń]ġ7z�ަ�dP:C{�=8?Ov��.ITyB~޿�B�uvg�Т�v/x7�tѾk��z���\��DĪ���B�DB�ٌ/Cl&f���n���j��N�6��:*�`>Z�'U��5>i (5Ĭ����Т"nY�.8�MKK

n�g�3�^.���Gԣ�{�j��7�$-�xW�������c�I՟�Py��{l���%K�aU6q<����m,�ws�u^�x��|yA����f�2��/�e�#[�L��B[�X۲��b����P��2��mٯ��%��bxZ���_	ǿ�p���7���e&mj	�;�/��C~ۖ�=E��HZ�|�]��='~'���b�5�
pI��qU	������V���9p�P�o��b�I�>�[h=`��ɷ��Hl�����PR���:}|�6�U����&AW⋐��|��:�%W=+��Z"����Q���3Xn������Hj5*m҈~S?>�U��.#G���������gX�z��Z|�E�<ܼ�Y{��q�
f�ljrj�DpE�ݙ�2%̹��CU�t��?v6�m���/d� ��Ka��z%΅�@ Ŋ��c���E��k��tp��_��r��Q��#!vfy/0o����&ӯZ�Xbr�5��{j��&���j����U0j)6_�,��ƀ����T$}�
Z�8_i%�� ����n��NV5���~=���y!I����w(�[p��"��$3GY����a��Y^�ꖾ�׏vk%���a1���b�*��=�f� hD@G ��$lx����$�PY�7�&<��*�k�)"غ]?�$���.œd��A@"XV̕I�8���q��h"�/�j+��w8E���3?P&��cv��`�z���]wT���O�m�RFf���ٮfeHP+��e"gt�����bX�l0���𸙡���Q��BJ:<��48���g�-��k�>e�`JuY"2�rH�^k)�C`�cm�����j��ߌ����n��L�Gb8��[opP�8ܹ=��|n\��~�U%�����@�b*ce�>k��O���fk�)�|�#H2l�$
Ć�ndxA� ����d6��y7�	#���{�ݑ���Z �.��5���� ��RtzT�s��j��C���V�a3h�� tDk)5����SBT��eW&�a� ��H��i�Wޥ�\v�0� +�o��LH�� �	ŏM�57�OѼ��/ו��7M�qG��P����!��Ϣ�O�����>>m�&��W�WRYK��_�@o4��$-O*Ҿі�6n,���D��.�- �\ X�j������:�j�l-���қbK'N����%��68,P�ƍ��}!�?
o�v�10Rk�]�bW��\��S�����o��� "�I�i#��ߴޡ�b4:�<�:g��G~�Q��Jwϳr�MAN�[@V�
��C�����n�"�Y����vP���\��	��g9�g�L�I��#L��b��P�-z�Ԋ�}�Sw��\��#���-��y�K����RĖ~��<%ws��H��_�2������w�+��\<[�AwE:@�����,sCB��GF���!��&*�7Q��#�/�:�{(v�1��y�/�z/���m�Q����\D$#����n�'I�1�Y*l��@-�Z,�f�%����Nm�We��y�߫p0u�z�3�ta���9��㟜�&+�v�ɧ��!�#�R|ݷ+i{Vl5����u�j7e�\�����8.珈�0ҧ���Z����m)l��W�3��<hn�Wg$�3()�_��QQf��I#�)|0G�#����h�s�0��9�K\��:���[�KG%@�����sT� ��k�Z�H���|a<;k�C(�`��)�<�9�=U�?�z�	@�'7��!�W+C�lu�Tߌ��{�â�� 7&��N���Dt�R�.+�_��Y�����O!Bib���tM3ɶ���{c>�9�:�������͢,�������Yo��lTj,��j �H�H�������n�A���g*K[A�LZy,����L���%�{�?V�(3�<��bAбP����{?��X�;g�J(���_t Q��Ic�.�_.���!����ҩ��&)������Y�~��O�[�	:��������T'$�>��XC\�ƪjӧ��`O�슬N�I0��q�uT;t�X1i%�kG^��W�ЊM�c�W��ci5W!�s��zp�$�
p�"Ճ�vĶ�R�&~�f��Ja���c�+�Mh��J^NBw�������*=�sˁ�w��E�\[��vA�N�_=b����E�yЅ%-z�p��Eei$�>
��;����L�T���>]��tuq%(�7d�,�G��I6��$��ϥ�'���-A���Ƞ5Ɯㆵ.���)���U�&�}��U�p��� IЉv�7�)I��GĈU����i��oK�,��2��-�[��f�o�~K;uǽ�-j��g`z]ہ�D}��Ȑ��r�*W�	Q�j��t���@���x�V��O��Ɍ�	�]4ǈ�"�;�o�]`�����;��/�����m?f��,��S�:�TS���3�zmQT�c��/bļ���[Vغ��}��ǀ��T\90�E��l�/�*�Y��ũ�S�;��!o���XۢP���*o���m�dJ�%a�m@�4Ǹ�[u;�|m��S���3���'#ɡuR`h�@]�#�v�_�_�T����Y�(%�g++ty�\�g^,���5:�O���|eV����n��3����MO&������e�6*=����eY���D5�}I.��#���,^Ŕ0T\&o�3�r�+�ZD6�N
�y'SGRo"_�V����MX��W�Z^��	�9�f�˻���+��(C$b����>"��"e�c��5�ˎ���fZ��IƄى�{ʣ�mE;}��9�W�&�0iؘۂ�Ƀ'k�6�Z#�UB {�R��L� �����G����ƈmʛ���JE��|]X�6o�1�P�U�t��a�˃&N/o�s����O�%�N���lH�b��|=\�o����+n�+D��]��[����\�W���+�]��Ow]�P�I����˿;��aM��k�D��ǧx�APCH�Z�1[6�t�oHH��?5#�]����yv����U��k$c��݈�q�u��]�1�+�dS�%AI��x�<��「u�f�ʘ_M>��@�R��ӆrR���؁V?~�^
���>�Lg@H����,^'�"z�8tl�t6�[J]�S,u?��UE=��x(��2��AF�(�>�x�JaK�UB�R�/�S.���\���}�[ �,R˒�xہ���2�#����,��C5�{��`�{�VRZ+Ó�
�vE�3A ��W�VU��:y`�67����LO�4�j�]�17hf�^��F&�h����˅�X( C���~��Y�d���vM�o+����C�}��B�X�����v�B<�!�IBBTt�����;�zt��< =4�I��V�}w~2OWڢ)p7/�it:�moA�%��������*"���O<t�6!���o3Zr�MR#�uR�:^��G���I�Q����/�6V������@ͣ�	`M�a�t$U��dO�����x�6cv㍤�{l��eoYn�ʐc b̐�T8n*�#%uո��*�6�YU{���撫i��)-��o����x���s�g�+�\�Ж�l���y���H���B�G2���� �ڛ���:ڶo��0�f���ղ^]���B����(���]5����S|6-C-��RH�@�U��M��Qa��,b�nG(V���7��𳢁^;��X6r���؜��J��l���; �αq�%�+����rw�\���6<��0��< Z�����^٨3�Ӯ{_^+^�&�J
��m2�:X;��d����y��p c}9\7ޭ���OT�P�f�8N"�Vd<�����|8��C��IK����M	�����5�E�Ň9��i�-?�9W�����;��S̖�%>f�>G���6��/,��c�kloDh2�o>�ZyL%�pD�LW @{��j�f0\6�1�Đ��Q��V���<�@uݰ����\�R��[�����d�<"qR�>�K�WQ�T1�_�P�.B���+;��m�O��0�Đ��%��>��r����(TP6s+����PvSB�у��G�ڣ�z�$�
)�M�.��a�:�ڋ�f��ϱ�3��Gm��^[���5������H`�y����`��^��8n495�v��/>RY�Q`�R�E�3YTD2H�"s���k��V۩�jN\��\:�usܞ���'��3�E1�-�T�z���g6|<�x�2�Fv��9��/ދ$�=���i ���}$�����x��w�8;���~z�h�~x�j��M��A}��%�X3�F�8B���������dN�&-4���ǝ�y��>��7��b�����3� �S�#�ѻ�"m��o�+����8�����c��=C�Dהfo�.��H{o6�ފ���IrM��F�m�Xᩮ��,l������|�c����X�ʮ�{^(�y��F��~�v7a��7�Y�mI���g����C��ᆍ�%7?V��'��Ah ��ڴI���q�wA��*�1yK�%p��rt6:W��g����e8B׷fe��Դ{w�e�˟R��Cy�	wl�E/�/8sL@ffd7��$��dS��6DW`7���H�_��1b����lB��o[$�ik��Z��m`� _�����hL�ȡ��S��'̑��<����3m�/�!X�֞�,kb�s��>�½)p�,��O���)%}+u�%�u�q�G�m���>$���o�����`p$����O[|��<��}Y��zyς4�'�d�V��ϬF�:��Mw�y"��MnJ�@:s�G֖��T3�\$W���������ywԁ����X�1���{"Ft��t<qa���c~��ͨ%0h��C��_l+�0�k�-�.Y;]e7-�FW�
�8'�5/�6&��A���y�����d�ak3vh���չ����B��/�D���<'Tć��yU���wes"�Ϗ�QGQ8���K;�0D#���տ�?S�5���+#@�+K��?���c�9 2O�J�j��2j6�]����}
�K}�,����tN�`I�T��H�l�e��
>b����L�V���r��s7�xRm�����	(�̕<��o�Ž���S0"r��p���P%�����7��♳m�2O��WU���=�4�&���΋:f�$ b>���.
�c%����&��S`��l[�����s�6�m|ƽ6#+�Tb0��JI������՗��=������ a���z����1M��msm@�fؼ,F!Z����8fQ�2�3H���;7.�0����apm׍��'���50�LM^18TaA�\���:���5�D 
���.	<::�c�5�*�B�.�o~��<WDId��0�N?��m����^�c����5�<Nn�0��^��Z�^�-�dɅ���\�8���q���J��&�;u+|���8��Ξ	J��Ul>��}(/���xf��+�c=���|�s�AH�>i�p�ga��W�������84W��4&�w���&od���i��>������p*�}�2���v�ց;�=}%�4N a��誒��`�PԊ��|��j���Ȓ�݂)~F�M����I�4�����z�a�#��c�-��N����!޹cD ݺ꽷�<�i���Jq����y�$����; �	臇�f��fx���q���̅�0
��9Pn�K��_s��r+����z�D0���/'�|)^M-uyN'�
{&��r\��P[�xȧ��Ԡ&y�=�k"��cT3��iO���kz��� u���������B�����3����D
�r�D,��U��!�]Hv���+��ꡗ�/)�>�$�d���
i��]�3��>��A�z8b;97Ca�*�b+���$����o�%)�_�./j8+k!7;��X2j�T�T~+/����RnEYl[نZ.�}��O]�g�#+ ���Aw�/j��ȃ�ԧ �@�w'�Yb6��p��C������:�x�$��`�֛
TBl����;sW	%ݭ>M��b�a����7)��&�{�ӂ)VԊcr1�Wy�*��PVכ�u݄Y��TK���`�L!��������R?^Z�J[U�u���y�O��|�U3��CU��ΓxĖ�:6�f �e�늊��?�G���6_җD�v�7���������;�Uq�-F��6���;o��6N.:\��d -�&�7_f0���޵�yᏩ:��^Uv�r��5���B&�����$��(h�����MR,�㣦P�S���5;�+]f����'�������ե!Sx������.5����������w�U���.lDj��z�Hrw�_X��SL�ƴD�Ҩ��YK�V��`���!�߫��m1 ��f���L4Y�F��;ԟ��3�2߱��1��74�{�y�kJ����^�`d슓�~�EVZJ���oi��j����%:KF^{��^]Mq����cXd�`-2���yk'r���jn�_�s ��j�E�wz�N�|�'b��tO�����㚚k�8�o�+k#
�!vnS�aupB>x�\��А�}�C���AH*���"w�ntO{���u��{��F�;&����g�M�O�$��G��/9f�lLd�p2/ō\���џ���Ɣ�p>%[�p�e�����m�\1�T)$��&�������[ ��G�S��?Q[�R���w���E�,�}��'F꾸�O�:�0���PC���L���!���ᓏ����=�J�t���h���m^P��Gh+J����q�ƛ��%�w/N�ˣ���H?w��r��1'zq��c�=�zV&����C��J�́ULʙ��ܤ|�����R�ءO٨��L[j�:���@�׭.�6�0;�ȍљ��K�j�c��F��l��lʘ���HaWˏJsv6��#H��s�8���ݭ�صNJ_�>'1$W��"I��<l�A�3�Y3���ڼ�F�?��LD���B=;Q�t&���릮�xGt�ྟP�hC�1�����r�ח�-�4��"�-�\��6)Pn�ۀչ�ݰ�u\�%^o/��.�%5� Z��ޖ�ೇ�E0�?8	������!�;Q�l��o�)y�M�$b\Kno�"�N����Gt�2�k��MJE��n0V�i4�넱4Ԏ�/��4���8g#��p���&;\��:�t?K��u2���P�6">����Nu4N�6=�uګS����|�2�M�:�?r17�2��g� Bs�U>�s7�9	J1��;4FI	�=�5t�6���6���cM`�L��[�h�o�.�؊ֲ"\R	���Gl\p�?�2+��w��f�۰�H�^=�Gm
�t�=J�t��"��8�ǀ$�J�M��,�ɐX�'y��N嫙d���	�7�ME3��-j���O�����(^=y��l�N��N
�D+�¦ê��{���4�s������bD�v!�f]6}���u���|��D��t�8�޵�z�+��_�಼4j)�]�:o�Mz��tYz&,e�{D���R���N��6ͷjH��f�U*<(rk����aiW=z|���s �T��pƑi$��ޚ�
�p�o�h��{AI��B�4�P�p��ܯ�`��P��V�����H�z����7+"����bW8M͵�h�*� ���{6�U��6Z,e�6��p۩q�i3-��.m�D����`�pۃ�'���-z�MX�-��s��y�_neT�0r��a�Y}99g4n-�T^&MZ�!�U��*�P����L�o���}#�~Q �䎽�V8����T��qՅ}�O�u���?�}��x ���ұ�Jh����4��3Z������l�/�����:�Vk�t'*.ﴯ4���P_uh���u?#�0���"��s���
��nNSnE���r�F&5�����w��J������_�����8Ј��͸��F�,����ى.@B}��B��G�E[Rz��9��տ(�j�_:������o��(_�����O#�����!�%�h�pt (�Gݏ�\x�?r����t��X����A�n ;��2����ǯQc-���-x�G6s������8~�/�ky�}qr��QJٺ�M����r_3�M��;=1�z�Ɍ��@�Z����oi%T���pN>p��RA�y��?\ig�*'?r�%�:J��uV�j
����<�m���'h�������>����w���D���ݩ������\%����u�`�R>_��Z]�C�Ahj�`�[ރ�:������&�ePf�����t1�� ����v#z��S��͚��K����Y�r��5�LzP뭩��Ĭ���2�/��ƃq�@X�$J��<�T�DV܁�3	�Lw:�1�7k���ZP�<��x���P�hG�y�Ui+;��W9��=	<�-î���bK(��8I�A��]���;1�Z����dǎŰ���q΄��)��2IZ�_Ʋv6y�km����������0?{�M��OU�I�݋���M%]=y�-�ANWo4��\7��f��;���8ň;�9�8'�g y���i�i��>�շ��[ �be���r�/�9�z���Evp)��Oe�j�cr���uK��&��;���*��ʐ�'�ݥx�w����&U�G�qM��|��k,�%s+�>� ȊO��M����m��.���d��F}\"�74&?.M�4��ޢT$0�8O:�	D��j�俥n'����U_p�l�j��43Kq���{�!>��/���D�HnՂ�j@���R�5ȥKoCs���[��CJ�;A��y��^U��}�(�^�dH�����̾�{zT�^��[XM�6���jdyz�����v��]���g*"q7�T�=�(�&�t?�
S��d�kK���$�pP+Q�U�IJ
�����Z��""
BǨ��,�ܜD�Zc��y�8�Ê�:���l/G�m2�Al�Ev��`'"X���<݈U�h���"�O��պ.� ���Ncw�8A�A 	��s��x�_"DX�h	��`�SZ�z�xE4A��/�T�~ka?v���6)����Ц (��ܙ�Ϣy80�0V���|/xє�y�jb�Je˜iD�8Pn�k��>D:��#m&P:0wo��g�+�+;,9M��.eva��R��N�_�82�:�2��8
?a1U�(k�8�ṃ����Y���Q
B�ɐ���eU|��3	Q+�6�c�L�B��t87��r�/�D�%��'�Jg�~e�>�\a���XזG�w��?� �)XҨR�-�xE�O)�B�g$K�rTZ�UJjfE�a0�W]���Ί5|�G��Jf^!��Bf���M�Uei�P19F7w��ͻ}Ra���J���3�1���-;}�'�?��dn��}���%���c��(�0%�Y5H�c�F�+G�}�!O�I�����2�5ٓi��
vwy��K�؆O�i�:���>�[�ͣ|p4�u#R���n�o:���.��m"36xA
(�KǟS$��	�ţ��+�Fη����K0�|@b�qȎK��ZM��jdPy�Gƪ�T����Z��F2��7��Y���G+�};���xRI5}cu��#`���h����Xu��@�~J��Ó��}�7L6E�I�'�'�Zd|�@��Mcpv6�ʝ��،�����B6�^Kf��pѥ�oLՃ�M�B��`��y���c����G��}�`q?9��y74k�lZw��E����1�.�'�z�Lu�� Eg1���Wg� ��^k���Y��-�t�m���c�1���BG��v�a9+n��$pa��I�f�͸t3#lvU����$�d�t�\+rށ��<���??s���z+�2�9ќZZ 䡧ɣӀ\��~��sy=\[Y)��Jہ%��"�8��j�z	�(��n�()�S�nKRܳƻ:-[�.y����p�(�qͭR���X�q��wșh��▛�p'v蜿�������=�ɊQ���Y�#���Ǻ����G��b��Q&�̷�{�,d���i��^B�C�O����lN�7�1�N���y�O�M�%�f�l�js>Z#j���NO<���md\�@
�S~מ&ͨ��(8�Xf�+(�G��^��d�Q����߫t�4h����<���&&�?Z�@I������o���P�þ�GIn�ܾ�)�k����Gvr����20�.d?<�i�/���c^+�l	
?�t�!j��Xx a��a�yB�f+��Mm��.��� ����
����~3Q�"pm2$1���1("��~�*�:��/��LT��a&�ͺ�<- ER.60
<s��;���Q$��ew6ɉp�u���dȱ)�K��P���Q���C;k���E��i�������H�%^��3�P.|�^�+<����G�wq�����=!AB�ŠX8蛖��)=�?#�z�X��'�V�4ol�α�1*���ꂀ��Zj�goVܥE�d{(���ѧ�K\L���b���{�j�`�Ț}@m�� ���a2X/,���e��#�tGsj�-#�1���1�� I����t�3�J�NR���b��l%�,�K�����Y`���?BE-|�Ճ�H�if}?t��Y0�*�D{����U5;�Q-.��.�\���5f�~M�C�5잸��aR!I�h���Ҧ��C�!�`|M�a�0�eV�z�q���~pj�2�1��ّ����E��ktz�>��q�z<�s���"2d�_(�)��9��s����t�Pv^���X��e��W�M5io�}������W�K�A�r��Gê6��R���7�N#�g��I]�||2P�!�m���Ѿ:���ǫ5�ޱʥ�ufS���(�Y��vu��7��Zܲ"�<���Z ŧ�PZ|�`��&%� l�y�4�C�٦R��ø�[��7:��h-�Gہ��Rg� 9�	���'��9JEn�c���ԃi�԰~�I?�qeL�C���o1)��e�-��x�N��EB|�ޜ���U4� �^&^���;P�&J[G��~yx��+q?י#0.S�E�hO�m��p�!8�#Rn;�(�{A%���
���p}"hzO�Q�k�%hX��r��f��=���q��A$N7Vf��_�O�R�����\��w*��L3ڔ'��?3�"B�A,�u7m��2��;�sb�.����c���hNe�:�d	<-�S�XY(+k�H�5u�u��i�(��Q��'�����Dx=�ɿ��A�O��XO�����0-F��Wc�a�Y��ܳ4å�-� '���^ ��B�ҵvor���<��E�Sh�*���,����l��P���,�q��=2��T�N�J	�(�(��6��C�%� ��^����N���w`;)��>�y	1	XX��sk�C�Qڑ��H�r����a?���\P�3qQ����Z�e��͹��(F���B+����쾘k�^+O��ڋ�x.�⫑N�(�}鞼����!��X�!�͡���,ل��v�ʛ��:5�;��Kn��cR�Ӝ~?���!�uj��Ȳ��BDg���5��>�B���-� �8�t�};�U��e8V	�#aF���C�ԃ�Zt%R2<h�X
���G@�㸷�W���g�݌x�	�]�Ļ�����n�)�!j&��W�U�,��[y��Gݓq3a��o�Q�U�o�S@�5"�p����x�k���;��^��QH������J�Z]�����W�(M���=&�rx=����2�1p����Oo׺gӊ�[*Qΰ��=�5駗���us~�4��r%SMc���u"V�2�����]�Ҡ�$7�c;�f1�k7~�ԇ��Y3$��yK�t.3�2�Ȧ�S��gu���vb=����0c�_5f���:�	����*c��î�Ic���_�9�����Cx+�9dR5�U���U���~�_^,����A�&d��*�m2W���voJ1�}��n���Ӊu2G��9���"��ls� �a��B��<��f*6�kFv�J7#��#]<�/�iR�rQ7�9�
��p����Gv�f%'����P��'��|��>�.w�W�J��Č�I�.��X�\fö�]à���c���F|5����Z�-lW�S�*�z�d��T��t/�d��+�j�Z��u��&c���Zg�H-S_n��K��6�R�Ł���Rf=�,DA�6�p�+p���B��T��/�L��o#ާ�W�G�Z R0�ڱ	n�J�S0��,�K����}7��J��O�ыSml���I$��A�4��%~�+��J{蒑,d��񆆑l����;��f�t؉J��	->]�vU�:p�n/+�d�����InO��/	�Pp��1��B���v���o6y��	4�w�C���n�TW�p8ǤF�Q�Ϩr�䌎f�-̲m)�K��xCj��¾�·��f����/=�`k����i�T����%��n"��������B���T���qƴ=�.Sv�z=:߯�@%�:�r�O,m�I��orTӅ-�)�u�<����i�J�<�w�`��eF�}V�*J0��E3��W�x�;nx�u�Ef���� oׁ�?�I3� #��c˱XK$���>S1$^�3�E�13�[B���~7@��#�\\�����b�KK��wGd4��6��Z:��ޒFW`qp���r��SǢ��T���s
c�z%�%.��C���Zwi�(��f%F��\���v�&��'#5U}xޔ�������c�"G,#���bT?�8[�A�q��I�wdI����Q
��X�	��t �W����=�OC�}8t�f����,��o���쥏�&K�WM�,����&�n���@;��e���^p$�#v-�R�/��f�e��Z��կ!��Dd�$wCM�艕���8�����'�]k�Tc���p�-�u�vz#�S���Snt��_�=�����V�aj2)��U\��F%�:il6=����3�O36=&�B���A`�����Y�� "KrF����`W�X��6� ���1WO�L���tד#Mq�0s_<��6!����#S&�.9�]2��gZ<����?h��myo�y�B��q$����Y��S,��_��xΐN'<�/OQ�~�O#�J#��p��nX��ɐ�I��2�|`�8��Hj�r���W���"�e�[�pI��Y1P��4��	�#c�a
	�u��C���2��A�5��雇�v;G��s<KwB>�e��������2V��q�>�Q/
V|�����8��J}}$�lJz�3�o��ߋqM�d(g��+�zw�����t���숩E��
�@�ЄX/F@j�,�	�Y�
x8�3}�R�XP�"�rA�a�߸߈�kj�{0�����W���QWaDv�;�Xpt��o-X�b�����;�;!�P���X@#ſ�Uy��АҨ��LS��i��b��Y_i;>���x=[;å�/�(f����n��K�*��B�cG�6諂vP<̊Od���?���}������%��~��Mv20��o{8��4�~�6�7���%eG��Ge�n ���zL�5"�_�}�<;����$-�M��L��%z���b?$I�*�=W��M�E{�g������Sl�9����Bյ��svʦi`�m2�I��K����dM��R�@@��"�7���ʄ�5�^hW��7�i&�kNXl�<��Fk��=I	#�4B�(�[�Y8�5YZ��#MA����$����U�;)ָGl��Np����Cd�.���L��e<��|�]�X�ԳlwuV�Ɣť� ���l��NExk�|L���*#<�'eU~����}Qq��(�^bɐ4O�R/tE�j=�Ƥ��oh�niU�D�T�. 2��p&Db�����:4��ڪ㥙pd����|�
c>�����+�c���^!~����t��h���<عnd�@�{>5MR	��a_X�=�<'�TzO�/������R9k�!��٩$[�8s�3u�d�\PkpE�n�����Sb\׳�T��=̾_n[�dr�<&��$���v������4A_�5���j�yn�&�ez|��_�A��5s��]��Q�.p+~����꿌_�f�]\� ��=թ�<�"[\(�ȇ6e�P7j�NI���O{��J��kY��8�"�p9�-�'%��<O�=��]>��hi$���"����M<}h_���qF}��{gΦ3��B�$]~V��:�z�K����;�}9�����"B]�`����΀ �J����6ZNfp+������F���9�	\M��ĮR���D0��	�\>1��<�+��GL;��š����k��y�����ጄg��p�k	���l4�m/;@B�2`n'��;*22v�~#������
��`�7���5����|ޫǂ���{P�UҪO�0E3���^��Ά�fkXq�U2^�%��pk@j� M��¿�?�`�o�e��yLJ���YD�W"�G��&Xz�� ^����vQ�\��ȓ�#�1:z�X�K1*����Rʢm�Tb�0�NS� �;��|�J:���>����|��DB�1`wɸR�0�g�u���uC��sU�����V_��Gh��f�����T�`�P�+%� �$
 �=Z`���
��H���^� d@�i��~����Lҳ��&�D����1���+V=����Go�^c1LU��c �`Œ����մ`�ڼͳ�a����K@��-	B3��3�BDܦ�Ԋ��>�M�w����D4����2^���]�06:�B�<�#<����.�Z���R�6J�l}�%�4V�E�/��ִ�
i'Hy��*���s��o�����.>�4fFW5���
vs���)���;��V�u/�t[^/t�H�	e洯���Ћm��[޳I��UrM��/Fʆ��m�p�b̆M끾4)戏1��vݯ>ɛ}��fHb�9S���s�Z9)b���>�ǆ+e`�������W��^p�ޔ�sҁu���
��D�ȷ`8�oFZp˷��_�k #�����;O
8�����~��h؍�׻��{Z��N��1(d´J"~h��е���%C���P�B�i�@����L��=jgA/y�[�s$/ǌ�%����(�P�ڗ�m�n��4N����6J�|
�B�)dE������LA������	����?	��E)��9N}#�&��U(�y��M���c\l��J�t�(��*"�+ZOcx�H/q���p{��2�ȩ]ɼ��u�Cq���϶c�"-�Ơ->�K[ܖ���B��5y���$=����� ����D�bO Z�?�@L��p�n2f��=^�э�eב���VR��E�&M�w�8��\�%>�Sb�W��9V���ؒ})iO�h��'2?/Û5S\��+uu���(=}�f���ޠZ������iu_�T�M��k����ު��-�<���-�U�E�	�f���d��ߑ̒"����A�E��Zl*��O�b.�h|�z,8�]F�7��(�9�6ɗ2*!u�@�d�մ^c��Om8��W_h㜂�b��k�ߞK�g%}K;),��{^*z��0�����Qb�}9�d~)�;��E�g*�	����ަ�^��rPEx���W��O����B��C��F<��}Z��(l w�*�>cąK诙`���N�@��d��f�Q}UjJWf����2Y�n̐�{�^�g}�Y*L7'ao�UyA4lL��-g���j5֑�(JÂ�TDE_��g��*.��[5a*�呻�p
6=��c��|5<�W5@�D%���6�t8^	�#��}a`�B^:i�p>��MNߕ;��T:wl<��$�
��y��`��SfN@���>��"�w����PU����`��Yxxuv�[��C�Ⱥ=��6Ys�	�wX���mh���	&�t���5�9G��H�㢴�3t�ǳ��~�M�a��4BY�!��9D�l�oA�Z	�����^f��cрe�+8J�g[c���"��kz�
�z�2x2}������{t���s~�оV���
�tp����#���6�,P�[3Vڄ���m����0�F��dU3c��7��5�����;eHB<K�JP���g�ܦ�������+j7Dԭ
*0�
G���p��J�L� QY��a����#�W�峩']3�v]��9�%���X�˞�!���o�&5^#��3`)����)�����!O�6pC���y�5�8N�����KϮ*5d}ԗ��QB8���7�h�1�A�/�7۳�����3<�ō��]��{b�Jq�׆b����� �!�p~D.�"6s�%5�6D}ύ1��i�J��#���at�*ze����X���l�_�4Cu/��3��j�9��տ`�|�wq�=�O�|����Ss���*���Z8r�2�bMQQ=G�p��i�.�[NQe̓�dԍ���~�e�h�6�Tv|/�8:0EA=�nb��e�L���6��S����c� �!=�sHߥ+ͱ�H9u�#��^Ͼ��#s�]w!�*���CU�F0�.`��8���D�B& Ɍ���2.t��p#.j��?C4`��]5������u˗Q>Z��.��ф۪�����tÞ����dr�S댷���$��L��:�[b��a[�|Ŷ�Ty �`Z�>}�!ۮ5Z/r�L��}�K���1�a�ʴ5tC�yݲIc�W���u�P��G(6䁔ۇMI�4Y��n�~�x/'8��|o��>��H�֡flk$���U�HrJwoS(�a�yB?�s�2�;�]�G����9-"�+� с�x��:������yRaQ�?듊[_�-o �[gj���C��I�[�t�̮�ء5�6A�d>^rZ&ˍ�W2�G<�7�z���F��& w"�E;V�bPQ#H�:B�!i��  ����jr��h?��L��\�8,"m�����M���;L���4 )sk��rʽ�ao3."V�lˑg�Pȏz��� �m����Վ9H�X:��ڱ�KE�uu�b�������$��z���1\o���}�<����C��N�4�I����0�]{s�Ov��*��A)Օ�Wǳ��7t/�̷�-���ti�t�o�s��G��Ќdq��+Q!a���!�L�L�'0/#�܂{��X�L��B���v�_��P� �{��_m�S�u�ӧ%�d�s�z��U����
���;�%�+r��*9�[�G��gD�1��n�����sMfb��W"��L@��O|��v{��Nn��ԧ�C�I�51�d��J��S�jh%40�⹲P9�F#�G%1,�T����G���I�}��k�lK�/a�p���0 ���D��e�_�s�R_�i$�@+g<��5��%�EUfPsYz߁_���_	����t&9U�L���ͬg͜�r��؟�Z:�n�N��6󑅲l��Ψ289a܆�ѻ���ۙ��C>+c�s�n v|��H�"�y���ޒY�ܙ���+q�̇LO�CӲE�0�Vi�/m|����Y�g>��V/�{Ze�x S�	�7u6�)S"�A�d�7jjh51���o�H�JE���ԣ���%~�p]�;c�Vx�I�;t���Nij0.N��_l���aI� ���Y�#M)��e�ܡ�T��r�D��)����,�-x,�H��PW��$13�EQ���	�(f���]^í��Y&^ɿ�]�0��g��=_҃��l9��p��+c��n-�|�&G*��Is^�8����;���v�*�~�G��`���ru���	 �S��=ȳ������!��{:P�ϐ쥧��#>��Ibo	ZJ�̢IXq��՚�6R��M�)�X�DJv���>�����7*�;@������(���{£V̹0����[.(�!H�[Z�sr��ZN�R+�O���1�?�wMQ�kݹ2ܮ31��Iw�r�~��ѐ�`Uk�R�ܸ��F�=����O�O
��dW�:y�j�ٷ��N��hg�������F�O��]�|��O�['9��x�t*>��m/!�Ӟ��s������ҫ��Z�|�����=�1x�( $%n�lf�r^�_�aq_�b�"��Z ���o���Zmx*ܲ�Ed��p�9�0d�� �7���X������k��n��k�;S^���i������:*M.���rq{���N�k�p>��q���T�@;Q�A����-Y��ta���dIK�Sa�qXd:^H��&tA��Q�m��rV�!!%�Ҕ"�vC�������\��m�K��K��gB��#��'j���T�T��s�"�����73�(�ʇf���	��uL�o�
s>�
��tq��1\=0=�X�Ĭ����=(Y�z��&QI�?)GR�>��0.�#$u����3]�'�r՞�����w��(����J뿏O.71:{k�J��w֏B2���3�/T�q@x;�����Q_���(�2��s�.�w���D]Ot���X�k���|�h߰A��>D#�3���+q�a<���oB��cǧ3=ɪ<����֧��v�B4�����/Ry^	7Hsfs��dW/�N���kμ���>��ǷA���Z�+3]���<Cu�f���>"�5����:hU+X�&���@��V�i��!���d�4�A�ߴ5_p\�����d���܉��i���vL��#:@�cꡞ�C��f
sM�8��n�2�N+��qA��NH^�d�{�Ty�S"���kB���+�bэJ��yJ�F.��=hK�$1� ��ԑ�Ϩ:$�m=�rQτVIX�B�ߴ�6�Ď���ǼNVweJ17`�`$ܺ��Io�r�E��E�i'���VԼ��A�St�٪�����NA|B�%l�1�+�ϐ8K�
�*�
��g7��x�x��Z{##(B����
)��0�!,�eC29�H̚�PaZ��V^f�|�'{�ҳ"ڐ��,J�d`�S�ɷ�����.TW{y\��ROtb.��"��	o}��5��W��K������E=���C�⥣����ყ
p2N����
��ު<�j��|t�A�����ؒ@��ט�� �V�'�q�u�R��*�M_P:���#�3Z�dA�WL�1)S��w-��kS�V��pϐ�����fI��V�3����ȵZY�ex����l>���^�������v��&#���k3/�Ry�9S%D�I,^G�c�.?�Ɋ��,�m�A��ֻt�k�вeoJ��a�V�.����0j���_��3�Y�t
.��Ϊ��?�qqGtó̳ٱ��K������h�9o���k��֑���m��٢���/��l���/d��y�#���S�C#���!��`�C�`��Qr-ПmL�����w��<�h��VeFՎ�.���C/��"b�=�� )d]��no�t-<0�g�-�ktɑ�c��0,���p#˒����_B��!�h��߆ ��~(d�Ť����ѸU=�(���+�&s����He}\�u���7r�FGz��Z���.�q�g�����s�Ni�k^iE&n�������R���2�5�)8"��O�����Z'��w�QF#*�������|FA����8s㾱�.���Ex��A2��CxY}i�#��B���@�h�����*4;���N�;;baM3���q�AuG���%]װ�d�~���/P>]�D88��WEp)Ҡוb���7��;�m�0�@�IV�b��'v��;��V(�$h7��g�&R�H�&`�W4
S�)���b��{�D\c������#�}�k�u;Z��O���S���i��rL��1P}��L�o�[��z� ho>c����>Bx���c��0�k�c���c����oy)~�_��V�("1��ݰ��ߚ������%�̏B����{O��t�H76"��~�|v�t����R�@ ?eo-.��D3l:S�ҧ����V��m��%T[1�E�^�C��"�c��q?51B�Z�?�o)!�;����4}��um���7��y�҈��D:�V����}������̿�T��4upSs=��0�ۚ�%AX�I�2"!����#d�X�gr䥦B�v�^���({��jx���YlM�z4Xה�t���׶$&C��ҡz�#��||n7Sl����#96[�t��;w[U�(�������!_�D�f�� �1�����nU-{w�uԣr��Z�X
Zj|E�3s�a�K�WW;y���"~��c�

��������k&|���P���j��y� c Z��� �i'C�P��$�Ȥ��C1��"��#� �^4��s`,zI[�R�Wc�5]g#FN=[� tZۆGK�g��zN<���^�:��3�Z�R�rD�CK�Nߖ��u�lN@�����u�~8�:ֹdn'�`�mog��O�����e����+4�
�L���L�޵�i��x�$È_�Zh �	3�>w�d����, �?`��Ǿ��hJ���<���N7�B�}���їZ��Lj�6g��X��W]����Uj`�;���B�y[�����&�$�����I4`�c�%£��-P��*b:�|̔��CI\�VK��}H����]t�͜1�#h��X+��L��\L�{R�601B��sb	!��e�i�һ�jD(��Q��6[]v̧��h$���Y6b�����pӎ_E{����Kx{!�V����dp�8Y�������p��P��ɽ��ht��S\� 1��,1}2�U�~�����|^1�8��h���&L0�4��kz���;��5���J�ˠ�T"\R6]�z�8u��_���9C�(kF��soh(?��8������ׯ�r%�P@N��l7]cu���{���9�@�{sYbR~E>� q)���)щJ}��}Y��Ra?Єq좶�1�s���ML2�DI��|�.����~�p�ӣc�9���z�5%����FKt7H�H� �$͓����<R�`�J_��޳t.�q4u9]a�(���8@���a
n-1�N���S�3�%��׏\'M�E�6]y��vZ���ִ\
�Qll��q���iV'�NL��b�<�	��J��Ղ�S�67A�6R��B���;w�k��[l�&���5�6YH~���}4G�r����9ύ#�ama�s6R��w��DR�Bu5���Q��R�U���T�:��<?���K�#[,�֔��NT}�oT
]�o����o池a�Zaܶ���N�-��0��Dl��0����$�do��Hg$�S���Ƥ΀�:������!N��/��eW�w
��P�?�� l�!�=��Dh\�h�	�0�W,#暪���f忚�K���f�$MRvƜ��)�k
P��E98��]\��<�F3n\����=H�~F�mif��`�nVm�%a^	A	X�$���E���8	 R�}w�X�Q���yz�פ6�S�׀γ�Ev�_�44�2��p���ُ�:z��e����[�,1A�-��UpBx3\���R�ܽW����RO���3�<������/��<C���q�:��ދ�w�����%�Ë�~�C�ǄMQ�CM�6OS�L^�^p[�S^�е�d~�6��;U�RuF!8���B���K
���$="`U^`Y�����+ˁL'0��{�
G�?��SA��	���Y�f�8��^o���j\��K(�w�	����8��^r�'�HI<�{BV�~�ۺF���F}�+$�,/V���N�g�_nj������qE������� �ӪVmh�{�p�ԫ\���)R�W��$ ߙ���%���p��w�?�m�p�Zc�S✅���ш�P�BbGP��B�
Qޙ�p���3�m�D�:?�9��hOSA::Q�$Kk��� C�6MB*EX���N�/�{�ͷ�+�4�5���LCԇ����QU�h8�m�~:q�� �d�	���^�/� �=�{���d�p�_�<r� ����`A�m�3�L+��߇I���m�K�[�A/02�$
5��� �3i7��ԑ~i�Rm�_�L�骅`m�{08lr�,"�˞mkA��kv�J��,<�@wL�y3�+��	�z�8K�|	ҷ����W��}����+2�����f������6��Ӂ<G��9o�������4oo��?������D�U��i�T�ǅ�?�>����_o�ӻ�0��¸�Nn)-TH��I�T��ٿ�$n�4߯UdpY�m���(��"�R�]a�ӂ�;�����Yf.�a��3B��w���B�V���@໩^��D��#p�F�i�dc�v;ҷv�N��� .���������&=�aW�`<>f(`�ϩ�_��	�(w�Bz�}���0
 �"
��2�/ �,ђqh�2o�I���u:��Y�~���xδ�ɶړ.���X�q旱��~�v12gc�)?d##�F)86u���5���P�o[�%g������Ԃ�V���Xq��qC��uL"2^U���;��scafA�/�H���j.���مY>������S=� 񚦪��5�QAq�ݮ���>ȭ��/����Á|���oz8�w�;�@m#d F�ɺ9�w���'�y��vݯ��`9���.)5jΔƐ��^���7�)G�W])�miCZ��Xe��oT
� =/�d1��u3Z	fc���s̫��TnӅ���q������&������V�3��1܁@�+��9w��i��/⢇s"<�n��ȋn<�g�K<�Ӯ�=�[#SA\p5
I��5D��"�'Z�.([z�A_/�M$Z~�"��w8�	���vV�c~����g�#:J��j�.���c� h9�$KS��z���5�=��K��P��{�B��kĤUQ��\uP���5��o�<��V���uj�1E�t��䵯(z&���X�@FTf4����3ѷ��6�
���s|/�J���zY?��E5�|��E�����~֝���	d�������� ��t�8��b��抏�����n\��U3[���������V���E��ª��j�Z���؍�M%����3���]z�$�kxޯ8�S\
���R�����rw	˕,8n�X�e9}^`�O3�U�T/���b����l��O��Q Z+%W�>u�nZ3�O����W�3���=8\|��;6���6E�7��&�.�=������K�C�p�L����]Be��6SK�tɆkǰ��0?5�σ�r�lĦ� �I,���-0�p���a��g{�D����Q7��9yoI�B�\?��B�5��m"a�(�IԊ ��ž��	xf������{��0���ņx�i��ηauBV�oG=Mxa�(�]�g�h��A���W��l�2}�Z@\�)��kfvA�8�١No��܄H�:Y��ٷ&��L���c��I�c�/:]�j�eN��|C�:$�g �B���۴�3���2;	Z�[/�Te������D�ڦ�3�3�4ȯؐT��k��Dn��J}����v�<WU/F9��\5<�E�H;�<7�{m~�	f+��Du!UЅ9엺x{���E)3𕊴���G��>ˠ>\�m<��9�n2���u=�ܙ�/\ワ��$~�}�)d��1�4��YJ4�mO6�V��JG�u�^�p��KD$���0S�p� }�@�pծ��o�Z��7���l
`F�Vh�w}����dvpB��!�o�Q�A\��p�2U;=��ѵ������vf�LҰ�7m�.�$�]8�Lǭ�����v��}�#�K!"g��^8AN����ttr-�Q��v���LʗP�h�K��r��ŨԇĢd��	Y ��7����|��zZ���V`d~ �ln�����k��f�:u��w��G��͟�F��ק;O<��T��
�}����wB}\\?9-��H�qC��𓭡X����XY+ C���DL̊R
�2��)��/N�݌<XO�R�n�T�vַ���צ�K��"	����"�z, @=���e�-d�s�|Q��W
c�l����ۅ�Vm���-�㽚��/^�ݠ�1_�����,sP��,4z�v��)P��H�`7�B��J@��(�T����z�ݰ�i�$�|E�h���v����9"�i�T�J�K۹���\��%
�s��c�m��vl��KhT�����U�y������~Z����?�B����pm��:�'�71 w����mi���^rE-0�{w{t����M�)ؗ�koe-���T�l�6�}5zF��-�
%6S�8"ԫ�B�Dۜ�br��`�����K?y��m��s�&A�O�57�^�7]YVu��S�Xx��ȈL�0|$�I�T0����T__*b�G�~���Ǹe.MR�9�dD;f�e�f6��:�p��A��./�Q^lm$��QBQ�:��aUHfx�s��E�NY�&�)RBiT!�������1��S�,�^*y����./͎��i,F�Y���h�V��͞m�=��W7Z˧��$�n�u���>&v��+4��C �a������{*�v3�9"���t�4'�����BM��gE�w��҄������Э��O ��F<������Ǚa���x�Ϊ |�5���P��PR	�R\{�R�x��+x����ھ��(C�p�pa�P�.�W�?\���#q	`ſ6�j#�^I�.���?F��'�S�PZ���ܘ�Y�@S�af`���!bF2&�~ss�!�p��Ǖ�а��#�4�,�J,�OpO�WrKc�9~�z��E{� ���A�5օv���#�l��Xu�m�����-��.�Ñz�&:�������I���\���
|���:�Ӆj�F����?��h���)�-� �(��gD:x� }�<}+M]�G�}h�t{��������Q��-3�0�Ġ�O=F�j6l�dۻ`�p�s��i\�GAB�	m���	��1;���<����1���U(��!`b�.5�]Qn�ݯS��9hT�bw�����s��̽�bv�m���"" sAvu��ZEN<	fI�8�`uXqi)��\vRF�J
�L��Η�9����I�P�5{����;�,$��)�zZ
&["�ٚC���b�qO$�q�z��=,E+���Ѓp����bY��. ^_b�MW�_���qϠY��_s��9E%�m���$�5-}�Tϲ�M�d���F�U�|�k��M�L��ݏ�0ɶ�&���y��.7���iFk�-;��W:��F�r[a���{k߉��%̬�Ҹ�_J�?��}�F��۞�����J�3��z# `��_-Lӏ��'���HY:2�0�9Τ�g]{݁���`#��ue�2x	c�1n����(5�i*�b�����b+��J�2�ܢ��{��	�5/=��O�4{��m�)�arޑ߇��xb�6�(�H��˓f6�f����"�{����q��:)a:�?p�ֈ1�6jm�̘8������ӵ�����&��߀R��ZTYv�n����WhҸ�PH���	i�Ky�BKz�5���64��Y�W[c2Pi��=�~0�/瞺��BCz�����dK\��S.jJr�-���uQ:�ɕ����0�}Ӵ���4&5pΙ��X��i�t<)�|^��^B�Wa����Y����,���Ƀ�[i���ʾ�ǯ{~x�
��|-�tԎ'Hy�.OzFW1�)�J՞ӓ�@6�;o����c�F<��?�=-X�7�p�YT�w�4�	U�� Yuu��%���(>T���i)�秷z�ɦ���_����&A�_霻0@q��㜜���$�u��Z�V��� ΀\h����m��2*ʥO�o%@�'Z/��BqI+5x�7�M2�ؠ�x�����*�,x�	Hr����{VX9�A���Pu���`��~��ņ��($\��N��J�;����,4|eU���
�*�Z8PaZD8x+��#�LnA�ƒ��g�'�>�O;��?�7���Ђ�^O~K9M�X_1N��41)� �6%a�D��(*b��J�%�t�W���תr	�C�Ub���r�Sh��-�Z�O*iK��a<���y�vS��E
��Z���c������U�,�����?�*>>�G����
&���[t��M:ʟ,� 9�4�ф�UƧ����r���quiEVr�:;K�d"��iC�Ɏ?�KԇxfR�jS4i�3u���"#������=�%���"��+_m�)�b��b����.���M�~�xXq�Vc�]�bz'��<����^x���4lۡ�������b�¿�2o���x�edg��˔����%O�!�a({�%QN3�¦eo��x O��gAj;��*b��#ZR79�Z�z9��7E�G'�&k?>g\�<K�+:b�����=�OT���<�៷�a(�п�t��]*���6�����I�w� �9�m��K�>
��ջRJ���R�d*�f射���щ��TI~=Ā��O�?�f[_�峁��~�v���S9E���h����c��=C3�h
pd{U��⎗*:1�en�RnH�r��ct�0xw>Ag5�
�#��!��-��E�쇴u4B+�u��PNtCaLi�T���~[�2��#q`8�,��y&�/].�;<]��1�_2��`9��1ƁUm��i�~��t�`�I��i�	/�Ҷ^�ҝ�$��$8$�j��է˓����Q��9�X��wX�d@�35j�E����j�����QmfqҘ4P����I]���`�p��xK(�<T��£G�$@��w�P\���$�F���2�G���c"m�0 ���Eϒˈevy.P��O�jo��0ϱf�1��d�]�ַ�rn��p���l��<pG��?�����=Ga��x����3��ݙ��1E�e;�$�>aX��-��:純&�ɨ�w�>���,����ś�}>�ʺ<���9�Ծ6 ��K�_����kX\�O�{Y�uP��(���Ε�?j}q����#�H���W���-�7LYlD�z�k�C��bم�9_��pjO1�ݳ��A�i����Nە� [%~W�pTv^�@i~��I���Xe�VI�}�,%��tl��`'��5:8� ����Fu㸚MZ�	�W�tJ��[U��\zR�h)_�6�A�+�����P�Pʢ��XО��gy�,{Tz6��	hU(4b{$qjg-��$�a��[EO)��=����<��`���^w�R�e;G��ƇF=RF'\�{B(+;�|2fq������NLm�'�D`�'���F�]��7��S���Wg�H�g��s�mςs����hy֌�䡟��I������ưa�>��>\Ȝ�.9P��Z�k`S�n'�>�	�vF��9V�l��W^�1t�����h�k/g��l�T��w:��H���6Q;��ѐ��t�Cխ�����W��Xeh��(�X0��A?�JMˎ��>L�JEX��Ж�3��	Z��c'�p�����s�f�p�g�Z�p)^,ـ�ʗiE�Vq[�`�SۀHW�G�s{���%����H�*�MSxӂo��T����\&jg�o�2��w�@��x���G��d���)������z9o�1)X��3����x=�(>�[c>,J