��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*{r#Jz�v�O,�X�F[prG>��AG�����+z��T�ͺ ������*PX���
�6U�8i��Q��-��8O�=%��)3�]̒d�|f�S$�J���lՇ���6���6����?��m��2�Un��؅��z�d7�c�a����'t���v�S������������zzȑ>��D����3���Xk�}���'���:^��˻'h��͒�Sw��(K�� ݿ�*�O�V�:j���	�CY�M�C�c�"���B�0l�9ݜ�`pL����OEL�A+N���A�K�UN����UMޚUW��*��$��b�����185�M�g-�B�{���AN��u�-�����uK�y�	$�%Z�ߺ�Ω�Ǎ�d�}��:�3 �|]�iH��ѝ1mR��G�ԧj�\@)$�F�=A�r��S��N�Z;�x�&�k�^;%���<[�l��逻���4�F��l��r�F0����='��0Ibϙ'��u��fm�����Bf�xI�N�������"Rc�s���|�c����9?�I�ƨq���ܵ��a��M��t���������+Φ���m�O���CP�s �������q(�)�F:U�J��^0�o��P�9�Զ+Af?`��Ĭ�2bf���k�d�T�X.�eKһ�7Q��hL�3矉���F~���:�.��4��/�ly�3�槖9�2�C�佳v��݌|�ј[Nx���i�н�?4�>_0���~,j,��	�[�p�O�1��2��w{B8P�Fa�rN�w$>}Եs��G��˚���J�,J�kX�>�;I�c��c]�&9kb�R���Q*���TJ߶����W�X�rs$���R�������@s��+"[���x<���%�8��9z6�ټ{Z[O�}�������Q+y��1.��d��UՃ�mF�U	���n���������=5��'�L^S���}Q� "�k���5�i�gZ	Dr\`���{��
����=b9>O��ģ��9�Վ=f:��%�X^ί�V9n�(d|ҲʗTA�	o��	�&�Uk����H3�v"�����\2�\�|�����&�6��7���c3v�ȋ�F�Jy���w:ƚ�ɋ-S�5�N��(��v�Y޸9����2
9
EQ���A%H�#l�Z���`]?eo����-���!��6��|�ӳ1j���:�q��­P$N}c.��W� ����($jc�F����ǹ@��Q���[��R�!�u�����Z8p��3��⣡��_�$�w�}�v"]�m���-�ʄ���x�d懞1��i_��)�"*��6jE����	��O{��5P᠑R���Ŕ�xъ��������=4�d_�%#���F�VPc�P�^����/S���m�p&��EPwXP��|�z;���-�*%��M8"��V ꘏�^�H���ZV�֊�g�Rt��Z�H�*9�u�v!HQ�J������!I�~�����׬�l�'�S4����C��%����Q6M����Q ���]T�N��~��]Iha�,#�-Hs�����ݥ)V(j_E'^������=׃��,�Hz������.�H85v�_@���Pd7G�ӗ��,y��Xރ����������~^����Q�ˠ7��H_��r(ҫ��=6�=��D6����R���D�j9A�y�ͦ�y�������P���`1���=Y��֔�@PX����.¯��3�{Q��x�,n|]&����N�e'f�r�{ў��C�2J?�Nr`t>��OkEHW��� r�"_��������?��E+>��#f)h�/��pֲo:p�ɪN�Mx>� �}5�L,����M��[�b���z���ae�?ʈ�h=�hs�Q�;'S��3���UW�i=�s'rzL����z��a�4Eex�[��8���v��Q��-������Z��_^��o���8��,����湝
3�-�$�.G�?��@�a��)��#����,����$v#�"�>���*�U���B|�װ�[9��Bc�5	������X;���n��y�����3�`��Oy�,���]�S�U���9��:ؽ. �E�fwL)S��N?�Vɲ����ܴ趾1N*tS�g:�Wۏ�2X)�9����|� [i<�2�=6yA�4�#<�#�1-ى~��� U�o��'Q��NOS��ɾ~����L8G�1
�y�� �䮙;���TM�&��
KX�#T�H�y�Ft��&3*��c�ޗ�cM�x�̨�,�r�3:��I�^�i�S�L|C���_���R'Z�v����L�e�]��VG�m��c�;h��{����w�?�]�>�9��"��4��G� 6{�sԙ���|o�Q���[���������Xx�هX���8�PZ+L��\�|�6c �gEh������VJ%�}�@�MV|���W��j�:�̢�W}j8^�xp�y�=7ϼ���!Wf��#�i���K7�Ҋ$� GX��Df o���Q�ji��F��澘䑂4�]��[��[�*M��g�z����+���b�to�T��JPj]����ޙ �9Pф4݉ڛ��c�<�Sx�lKcxU��K���>��G�-�$��]bI���x	��M��~5P1{��"Y��%�B]@���D�:�KT�j�k���`�?�,�)�>��J��F��q!l�� /�Hݚ �(e�m�rUi�J��3"��6p�����p������gBr{�P�1~Qd�~뾨@À�0�%G3����)�JT�*9���Ts�gG��c B��q4��7���0��ܥ��+�>�!v��t�8@%d;�%��^c��N~:�Yv`S"��6w~_�A��7�m�ْ+C&�b(&�9�����m*֙W9ڢ��ց��H��F��ü��E�6�{6�)��+��aC���.X`h���´�ڦ�xC���S���j�X뭬Dk	����8s��F��qa��9�v�"�[ɝ�
ܣp��C�Fw�W�}���<�}�h�J�^�d�D�-�񀟳���I�J���Y~Ր�g�6����<]��^H�>�4��O<�a�6%� ����Ų?��ꣵ�^�ܯC��	��MpU��Rl~��%b����d����VÓb�9�0!V'�Yj)�V��`wdy�I���:]�4�|nu��]@7&çR��e �	ġRM�@D�vv�n���1���^c2�V߫I�����7,@)��ƘΛ�*m���꼏��X3����u"��l���p�����x���S_N}�����^��'�b̳?$UC�BR6J�SɎ ��Mp~=/�HyuLB���� l�Ve�� q� :BԲ%~.���sU*�'�C���g(�X�i=�l:EW�T#�����N���WFqcn������:��!�?��D�q[�&v*ǅ?x������f��H�jV@�&��L���̱��V��KP��{�V8�7t��iu��r�"�IA�=37,�.؟�s��x��.I1����Tyc1%����YN�=6�.��f��A:��P�#`c��A�f��4��O�]�����z=X)Z��� �3�d�"�r6�?�=��%w(g��5�۬mV�ح����a��R�|��*��(��k��~����A0� �n�_������ż,=��+�
��NY�^�?�uD`8�;-'�Ak2��HNBT�>6�'�$����+�Ħ��Fznv��'��N�~S�Z\�W�c��S��U��5�`����A|x�#��5OLQx�]��NˬH�N�4a�:z�ﰐB�N�(�|�_���R�8�JOm�~lɰ�4P C�A���>�?�8��Qc�7.W�[�1�".���Pe�\S��@&�}�r��0��=��[$^V�_��^�M=yޞ|�{���������,�+��6w�wc����su�9�0�^��I�1߹մ��Aj`�Y�\�wHT�L�0���l�k;�O���c�����|�B���j	�p��J,5F�YM~���,�a��<�:�"�|L(y./��斦�E��ʰ{����P��F}#����4V��U�ނ���.F�.�`q�(�������]g|Zn/3��t�`}����S��2MЍZ�C��g�ʇ���+e���6�J�NUAe�g���iu��U'\����ӱ�+H�&�Y�TNgsy�������<\�O.���rQ�����f��|��b��,hM����w��op~�ә��)���D(�̱p*������J[��m?s���o�i���
����l�d)4W9]�G�M�z��WiH���nF����)����y���U:>e���L'�E���j^��5��C*���0�1nQ��͉^++�`Ƈ�|��3y-%Ӽ��mX�%�b}&�x��ۖ_�w�L�.��a�jWD���Z������!��+	�WI^��9�3�R>n��h!��j,�]��j�-�3�J�=��V�����B�Ync�ێ߬�6�C��ԈjU�,�c�:N�=�D��U<zN��c�F(�+`8��RTx-���~��{ݻo@� Y���G��6Sd4/^v��s�SW!����kx�D�@�v�5�L7a>C�]�V%5öW�$���_�
A�?���.�y���шE�j�#�{����HI���+���B�z E�p�"�H�OJ˙H��Z��A�Q9��~`�QyR\�2m^&9��Hv�ͳS=0�:O����,� �j�I�꟬avS�9��uA8Z��x%i᠓g(��J���%����=#�xɶ"�Y��]vco�wJ�<p�D�^��g���s��0�ךˀ�F;���۪�
�	J��t\͟"O���oD����!r눠P�@*M�y��(�1tn����3��v���uE�
���eKۥvVp��+4ot�&�Zݛ>���>��!Ռ�q�R����� @5�JN<���~Ώd���l�I!���Iq����\ϾƸf1.��(y�!i�>�o���X�4D�:U�Zw�E�R �+j�'�e��V�sV_^�(%�E�1�~y�����B<�& �Au�ɰX!MO��z�VP���}~x�S9���!���F"gSu^�j5b��$��}�Vc���!�_��؇�c>M0�f`�M#Ҷ���;ΰd�����%s�,v��T6�c�P#��r�uez�(��\R�|��~���r$���cc
�(���]����oJ�O��*p��o2r��Q�Ҧy"�"�ԟ��bZ�nZ���o$L��Nj���
�a�q;x����:�NN �N���~3\�i���Ƿ�F3E�b��gZm�ҟӾ �q���S��qr��ͻ�[�Pz�D�ލ��ļ�h4�f��_e(�DҒ'���3D�S	��Ө�9��#w��]�Ȓܰ��b�9�#�
h�����%��(:O�V��:��=�t±�}\ޤ_�aLg���
~�(b4&�i:��]Oz,X�Y��&���a)�tL��nU��?���D8�Ĭg�!v���8k*�B�Vin����J���g���I篛�i
(���U 6guo��芰c��@_7� |�[Y���(�t:�elAԮIG �S���g7D-EI�S/��N�����*�V�~���5�˓RHj&�؀;�?�Qq,�A��xqq/���=���r�+�� ��!�'(�cY��PU��P����dF�=G��Ba^������J�ah:��95G:�9�uL��[ה6�ǥ�IcO��17d"/��TWo�?H��glNaZ���^E��i�9ko{�n�,�'��K`W����VbVki��) z.wH{w�]������nd�ӗ6�1�1A/t6�&z�0Jz�q= �D�WB�t[.��n������� xG6rQܷ�A�%HN��-q�pte��"-�=u�k���]�l]��J`��G��Z�Ӯء�y��^�r������6^8�*���%��Z8*�@�� %��
�P��웚䀥�ط�0ƨ���$`�2 >8�n���n�>������$��4Q�>ʡ�m����9�؎�PM�IhF�Pk�wh��{�{>��uΖ��yލ۾�uh�����H%ï�?���"j���ba����OM��ܥ	��UK��Cu���e��;���x�%��c�q<1��3,P%���N |6���>�L��$��UI��9a�W�Y�@�1�Vt�'�rD�=)K����$ �/�+!���)���~��0
��9U�h�"�2�8�Ẅ́��}�W�Z�t�J���t�Űg��4bhNM�>��xQ*�]{�zXޯ��
S��4ȟ5�=sh�I��׋Ove.�w�JD#@�1�`�Z��!Օ$�&��\��c��ɝ�>!ꖦ���5�p8y-U��CS�!���I�����IL��a��OQ���%f˂�#e7��y��.��pkGr2�X��.������D�����t�V��2�a����M%�'ꍬ�����dĳF�΍Q�a�B�|Ÿ�Q`p�͖aUsl�A[��0�ߧԆ�Q�� ���hӯ����P@0uf��ciQ"�'�H��2������<�S��|�0}\�^���
��m��/��都���>���%/W���G(�:�ás}��y�i��5m�0�D��٠����0�@�5�"0F�PP=�/��Y;T�m�s����mt�N�f���9,���WQ��E�џ�_�)g��r��vY/0�L�_&�ӛ�_{�����پdS���%�T�#� ��#F_�Z���j@V{��*�Ul��Z�v={��,D�3V�>�8��5}Ӷ3h���O��_�
3LXmHbw�m٢��+,�,4f�c�rQ�GO�=!?*v�"�A�ؙ�6,$�g�v�;��� �}Æ���3 �3��(v�e�~37���g�<�a2_�8nd>,����B	Xq5�h�ܟ>�@�[���]~b2N��{@٫%��bi�E5���1�6ݚ�\/�U�i�|��]�ց��m$�w)}礨�ɹ՚��P9d�W3���=�G
�H��>��.D���W�_��'D����a=��mO���b��<���V2Տ��Q�oj-Q��T��@�5L)����@��\d��b�-u�`��j�8��NQF�����Y�a�
qK�U*�X�@�V�NVMT�hh{/��x��K�~6�5�.�;Gi��&�F2�.�� `�m�	�upJ]*�b���\|EFtצ�g:,�i�Kh��8�.^5�h� �	�o�V̝�iD���c�95`'������M=�/l���@m�8B@D|/J� �����S7���ڛӏ[���B!x��_�ض)���KW�#E0R�C�ORd�j�-���p�c�D��������l����-E��C�g�����ޙKh�*�"p��vYMM�JJp:e�k�Y�
�$�؋�[�����*���hCK�-X3��`�\�����%����[�� �H0�a�Ra��m�wd�_	I�]?�΁���'R�u%U��{���=��Důa�iy'������ �h*d�?ۮ�PG�(]Y���v�U�u|�h�l�.�)�6ȱ�~/��8p�xi���
��T��|R�O�oe'Y&|0�&��u�e˒A�|b��]���G�X�</=@p߯K 9�8�g e2e���rCL���A��a�qYQ���~u]�d�T"��.����adr���B����	{:�t4�p�`���'����g$�������P�Q�T��X+�./��4�B���o�V#Y������E� <�IXѫ�#����%"+�w��4s#��-�[;�K��ĚD/_8��~+���h�V0ur��qtE>l7N[+u��D��G^%B ���>�q���]	5�]2��/phź �~�[[�ɻ�lR|p��@_�	���&�⡛1��pH�uX=���fi����Ш�'=P���]6�R�!�A��t���C��e��Lf�I�?G�2�\�&sqy��rRq	�HD�Q{�(=��������p
�D"&���-eXz7�w��_���g(@ɂ�8v�=T���hM��/5@�WKUȡ\c� 0���!@�_���F!��CG������W���:I���"�T��]��nҖzW�fFn]�����tW��4����j��5�ش�BL �o�a�b� �)ts�p5ɋ3�SS�~Q���*ƿBJ�5�QJ
�t~u]Nj0�<5�ۂez_(���'W���ȫ%G�HxItZ8*����h��9�-
d'����`�A�v��
�cv�TI3�F�N�XD}�<ؑI3.jh��L�o��Lg�ٯ̷Ɣ��-���"sF� �a�`x���Ͳ�?���u��WV� ��A�����w�>
9!vQ����.yD벜���,���n8/��)�"62�����1Dk*#Ƽ� �G�oun��-�6C�U/�4�(߹���W�0(�5\ �P�}u��aO�I����	3d.�ދ$$�l��8�Ҝ5R�(��9��'�>�	�=���aY�3n�;I'�y$�Sw��Q���ӵ�J1<_�<����?å|��Վ=���G~�����Ui~�v�����K�?�X'd���77K��.��-���0�MleW%�Z��?i��G\j�o{|������������#Rj=�E�|^[�)��Wy�u��6�E-^x�bf{�:)�^�չf�D̗�UN=��kA�������3���6J��\p�k�o)/��.�p�*�1�Y#���/�=�j�|:����l�GB%�ʃ�W��Ύ�|9��Z����.���d��
��xm�w��2��c�4�
W�ݓţjz�ܝ&9�T�������Y�w<58va��n���{Gm�f4������Hbh�ҟ��lD�8Be�ݚ�����
���; �ZGrb�n�E�D_���Q8���C7F\	����=b ;»�%�΁�ŕ����7�� ʎ1m'��Y��"��/<p1�x��*��$�`T���%��s��R��[�ܻsJ����4��-�uyqf�p�H��⍘����u�b1�xW���i�#^<:��B�����&���C/�����Җ��p�Ơ_W����N��A"�	#�
UbSY[G
5��7]��$��ӷ9N��W�%|�iF��2��u�ڮ��w��)��q�z涋��Q"G-4��'��qnz���\U���mb�į�H����Y'�����L��gOq�%Y6�[�r	�A�e�I!�Q�
$Y��J�vLt%�y��p�,�� !�ـ���K;껝�?�U�9R�g��t�kk���/�GH�|�@G�q�����59���W�_$|��1��k�V��9ĩ<N<P%s]���:�.�i��KF,��K�n��y���5�7�9��)@影S�E� �0q�!��K����ߍ��ti�6�""�4Y�]=��k����r�2��V�x^5�8��b�'���h���G᫐��O7B<�b�G�JT��b=9��}9Z�JW�Q����%��}����nS����D�(�=>}�H=���2>q���߸\�uQ�:*ʚz�1)2����h�xs�	PK���� ��*}_�Xlm���5�*���t	�6�|ǲ�!u�Y���K�pƱU��#����)�:ܡ��/N#�����e����c�Q�ە�)�2z�
s���mw`O�dA.ї7��օ��ۧ>�x������ԙ�����)��v�G���~ffAP�E5�+�o�Qo6�.�se�=)����~2Si�����A���y;?7�)jc��C�3_+#h���yY�K�r8'��6�Gex�e}�龚��-�z��-R����,w�IМ�Wx�N�n;���G#���+K=�W5�
:	|����;�����������{!���h�0���c�aԛ��a�)+/��d��P��Ud�U��B00$�1O�I�!�
�\�ȅS�}Z�� �T�����Pcp:X�!��؋�`�CZ��M}E��/��\�ٍ$R#A]OV��@�6i[����J+I�ݴ�s})�q�[GiM��\H2*�C��%�����cS=3���h�D I��I�[q��n�L`k�ʎ��y 7���CXݬ���I �Xz�1Fu���ԺD��V������ֱ�?{n=�>ju:�M���Ԍב\mG�jH��.	]��Ah	S���:��mM�m�$���i��'}'�1��E%3���wP�2�M�L�+0�66h�¡�?�={Y*M+������H����Vz]T��0Ä�Z|r��`,��E�@���VY�oW��h�P�4Ã��K>��L�OTn�Arf��«��e��RH���hU��s3Z!���"�ّ��3@F96�9�@�*�l�;�B�w:�0a���f���4ٖ��]��u�ILV�$d﩮'<������ZX$�����* \%Q̾u�xTv�|�a�LJ�+!�<���U֑|��Qmv�]U��l�C���z�_y�*q�^�H�.��p�οNg��Y>E��]Cqx�M����p��_4�Z��@h�F�����ɫ��������K�p[5����|`�5`�w����t��z�t	��*}T���R����W���Hm7$�^��I��Hw}լ���]hw]NӖb�3�8C�}���@�??3�|?p��]�����W�g��5M���.��AG/���*ZE��u �ټp�yԫ�i��0�xH��?J���D��f� �*��⅙���!c����6jS6�%JK$�E��?����#)� +4ڦ*���jC��[�n��fx\�0��h�sq�ȹf,�{<l�á�ɛ�d.E���'YJ'	#^Y)k��ⴅ3�G��ۨ�&l/F>ۋ�� ��fI���g'/�)W��f��Μ=���ClƵq���N|`�3�[��6W
�V�Fێ�ǾU�2�w�G�99G?�}C��'/0�UV�����[R� vO}�Er���.6ƨ�U[P'>�s[�M)���;�Y3[�W�����3z9*����'��V��5ؓ���Ҋ&��0]��$�)�x�0�<���e �I#Ӏ�_�G�
o�?�I錪U��q��p����i�ʤ���q����A@)�g��$�3�uL����Fy�a�e��m\�QUP/;1n�����{��D~a�� ,���)~��tQ���X$�|�׊��T8�bp���u�XV�F�E߂�v-I¿��!aD,�D�0İ�ClQ�<�,�E�~$2��e�r��N�5W��[,9�>��H�� ��~����p���Uw��x)>� q�=|��#��kh!�,ʽD���BJڱK��zs9*L�<��I��0#�2��mcM�P-�I����78�l������ .^����ۛ�e��e� v6�Nm���\�'��`�N+\�T
�*�ͮv>����T?��=ϋGJ'x��4K3��V� \X�,^Q�l�9 �V�(���,� �%7�/ᴳ���Kc쎴�Ʀ�p��/�	�Eu!��a�x�K?{�m40}y�t����w�	��o�s~V�M��I�R�aJ齓�$���-�(��x��fJ6�w>�>��Pw+�_����P��&�&��j?����īJ_����B��0�6�%7�}��0c��˱��7	��1�`J@���&�
 rx��h>N.�騂l�/>��/�(:���J��o��y�g�ֲ� ku����F�� �d��9�B��&�/W����Dk~+)V�.��QG�oc0{k�N��P�[L8����� �����DA�FHp�qe�W�t�w�䂊
�W��c�)����`���2@���O�/m]��}���T�\������ₗ�k�=�E"Q�̩5�C0E���2+j.�b���̩4\����A�j����׻�y��i�՘q��av���/.���Ѳ֊V���0I�Q��?�Z$d]�a��9	2K.}�B� �)]�6�f��nB=
0�:ی��v�9��K/Bn+J�ְ�����]�z`T�%��ܯ��E�Z��)�U0�����G��>�W{9ᦇ%�44��B��
�
r�J���5�a60��8ܷ����8�0<+A�,?��q�m�k�f��ڪ�y��� ���y��DnOub�ټ)�?��f���]��O9-H�:Q"����
K�!���q3�4��2zl��G�t9�Ŗ��͋(��X����h��/`zu�C��R46 ���Ë+�pjf�v[��2 *�*���R� 7N%�b�s�>׏u���L([��	����h��})���C�$��y�U�/�������Q"(B5�#��!��\���	?�?�@��}#au]�/Z4��},����"y1�i�3ҊTHn!;'{V�� E������e�o;�J'LJy��Dt(�*ס��{s�v�i�w����b�r���f����E�Ӌ�)�o6z�in��N��p�j���YA�~��2�~~vZP�^}��h\�ǆ�+�I�[�m�S��*И���P&�x���40�(�~�Q�i�P�u``F'��0|��6+u5���T����-}w�h<�<�_�C7�8���}=DF�I%;y����*~M�a�c��-�������u�}F8�m�%r�s�㹜߈m�Or���Gs,:��W65o#\�� ŏ#d�U����<�=3zM�6�Hbo7��K����/�a��p+�JYY0Gy�P�������f��^��//.�9�21���H���<'-��"�
	2� �̄�*4[R/xߞ��(HXC� �����E])c�s��M�c+��O���i�L��ӿ���Cќm ��;�!_�d?\�|�8���, ��vi=n�N��e��N���'�Ⱥ�֨�`�M�a�*�aze���Q�m�ͼ��D�@�C<K�b�6���8�sJ��O�c��s���2F^y��	x��^�C/���=x�NSь�ߧG�S������!-@�5�Y�x�S��7�4`�h��W���@�����IVF�dhȪ�9b�	�'���9�����_B��7Y�0%�*���oX����H�1h;������n.,�e��qa%:I�"[%��LC��\�|�S�|2�"3f�`U[���m���BR^P��*� �,��&�����D�ݙ�`H`.����%}�
#�B1��X��I6{�O/���c�O�*Ȫt��K1P$��-4P� º�j�V,O�˼������p��,`=�׭z	p�8���i��w�Ѯ�����T<2Ϗ*4D��5�R��'x=zV��2�G�KFZPBǚ*���Te����Y��}����Iň���=��*FRU_�I�H�^���Y�.й��L/S��ҷ�F������aͦ�n!OZ�,s�U�֨5G�f��C�����q�M��B���Y��0 vmѱ�E ��K�8�	�*v�r���)����ͫ����b�6+J�{Ss�]�=���_W��dGfS�s����� �����s������c���nt@� �C�~���i����0�@!ۇ��<�6b�?��>I;i\��]!���P������ ��bI�����>�.�����g��/�StI��^�O�M(�Z"�����DXԕ�:E�;�#�Cך����b�;��ά��]�f���r6/cwǙ&�4��R>l'ܶ����n���Ee��j~���y���5�8|�V�ݙE��� -`v�<��=� ӫ��H[!ވzK�J_ҵ�!��Q���I�m��J';"ӻA��0VrB�F7VT�R��<���ụ�p1�C�[(}$�k�Zѯ6%.�Q�l&п�~��ްd(�&��p{�>��:1>��r������.9#c�ɉx��s���J�g��6,@v�N��:3�}e����Lه�\��
�jXx��"�g��:&��wġ��H�*P�ö�b�(Q,w�,0��W�Ev*.)�����E��W��&�[րR������u��wBk|j���>��-�KQzc������tm��u�E��#��!�	�g  t����k�#7�y��֐��6�rʧ��w��_�
q��g��o�;�\U[�y�|׉1�P����%��g��K�u^i�C.כE}̹�;�}߅����J��i�5ᦙ�@�W�nV�<�=;c�d�$�.*�������b�.��1���-���*Ze��Z~y-�#F0fP���y�?v��מ�qS���KhE��L�o�1�n:e?���� gj���t+����uDR�A(�0�I�-�$�L��0x��G��Y'q��P�G���m+�ͯþ��3��a�.Dޗ9�����!!Y�$x	 
%ƣ�c4��}:�����{_� vh�&@�p�9oҧ�Xe$,)MG�a� ���EIE���:8d%#V}�;��NT8����5cO�q$� ������iQt{@�Wq�C Ǆ0� �(����Ѯ؀�gG���u��G�_��n!0b��k��o^������88�b`�na~�#H5Zl��R�?�4h��q�L�M,`T�]|bK�����;�٣��'��e)i(�F�Ay7���,�hp�塣Aޖ��RO+WJ$*��e��KGTk��֫�ԝ�/Cȿu�v��S[�
�j�	I�Lq1������e�I�	�*�'��F3iQ�m6�|0� �w�<\yL�i1��HÏg����+.7?-���i\����n�[
N����GEz��Gx��͵u��Z���3�b�^R ��d%�V�w�J����k�W�8�ŮOf���4�^����տpkl�5��<2�`�S��@f{�a'D�qi!e���������_2�/$�&�WG9F5�^:g�h�͕j�q��N�v�9�#8��9g^��O��T!W�5��v۠TV����CI��w�ȴ���d|{���3��R�_�^U_h���Wߕ[����&�������K3s��zh�����5�8C7PS�6�'�9������������}{�}ki��h:����L�1=!�9Jw�o2��*�F�\k:�7O����K�ӻt����b>~�!���3�=��6UӖ�����"�ej��[ka�����N��Y��i]�1l^&>�����}���F?�Hl51_?v�)��L�f�?��Z��Lc%�1�f��N�t��Kq��g����.Z_ϼ-A�<X:z���:�4J%$n�r�쒳�\Gy*��E����/�	grһ�uN���Df6A������c�[v��q�;;j�{bm�f�/z����s\��S�� �ן������z%Ζ�;�%���I�0j5 =��}B]�3q(�.+1���'�]t�bu���
�Q<(��u��?l�~pg�w~���Q:2�&r@�X�ƒ;�|�HG���D��%x%Fʢ	Q)�A�O���^0�@�UY��M�m��^*�%������r94g-JM��
:B����Ut���W��%S����c".��1`[-wd�1%g*G�n+C�~�T��k�n
$k����O.Iu]
r�Yo;��&�5��zc�}�2t�d���_	w��얟q�t��
��T/�:�eD8Q�0���l<�����e��j����*D��q�%*�����}m��O�[+zA��d7}�*F��iԯ`[��kN�qQ�&�L�i�v�I7B#L���}�p31�?OYΤ��'8I��s�y���������5�<����m���l�%�n��{�d�'s�|ha6�u�%V#�Q+��7�>r�=*�G����h�t]���7n�7�9�J�N���^�U�v�5�zJ�ze�.���о����Lk[�J�9��hv�CqxN�/f���͗������S�˛�9J7O������D�G�� 5�s��ݮ ��> ��m
�DN7�^�nd<���5�\ed�tņ�i��`�wTXD��ư��Ԧ��h0��C��8-��	��~���/�G�g4q��̽�l�֫i[	�f&ܫ���lf@[�|��V����m��R����hk_"��lߢi�S���
(����L�Jiuťn�2򑝚Q��h溽��vO������7T/B�ӯ��!e�2��#���uq�m&��BS��EȦ֢�ſ���;��}�#5[���S�?��f��o�>��`r2Q���6,������#8Y�������گ
[�D��&c��=Fd�����-$�C��E��p5s�I*���]C<�~�⩤.�Nruդ�R����������m����`����}���Z�Ca�¡�
��Z���M~~g�)(2�-��ױ�H�2�,��L�$�M��8�6�!#F�.\_I���g`���-��K�62��	�\2��ɔĀƪc<��4یOC����#�*�öy��Kh��jgj��r���˅5|`i�eo�R�/�g��	�p�K��I���.��.�{+hy�a�Q�:����`�I�P$Ocg��8" �3ZH��d׻,:xA����VS3���5����I*�'��ܥ�`��]���"#)��Yo9�.�f���,m�Fu��o�|#.s*��d���N��.ڀ��`�G+N��=J��KlV�{+����WH��y��W��d�_5�|��F�4�ɽd��b��(CFM�4Ζ��]���?}&��(؊�g�|���7ݾ��4�:Թ�:=?�P\>�����ҁU��񳯚q��e�|cSB~]�E��l�akNԔA�u���)�r�w��n)O�X�1�\ ��;�;�Be���u�J���"	�v~r��Z;X�cf���ԧlv�wQZL���3=��%������L��(v��K�:��z�5=>�Y�M���M��gX٣�x�ZMƌ�XG(?`��%F����k���+ F4iF[+�S�o�l�O�}BA�u�⏥�ao �*sΎ��<�q�����%�`����}�?d-��GT!{"̋-�g@J�@�o��$�����mۄ�T�w�?YE��{w��	��/����_�*��vt�?^���vI����d�a��[Ρ���-����,|O��?M	��G�|�C~�ّ���ʨK|��5l��P5+-&$6��\��~L9��p޻f�v�p6��%�F7rr����ͧ���G����X����:���vʚ��6�G3���������I��{����5v�:1F�n��V�Ӱ<<"_ؖ\e�kOKh�����:Tv�1�bVf1��'�	H��+L��|v��W;�*���K�3�Bv{!�4г��,� �?�.�7-�CO�/2C���cl���=�U��_&J^���=�8�߫��i���(�~:!�۟%dv�rp�4�/�&���0b�O��ocg�׮g�R=^�G��"�O�!F�i����M���_t�R"��ω�~�`C�t�v����hM�J�@T�(Mk�)d�-�
�gی���+���	��F�;V�KC>��u^��HX�28Wǵ�^����qiQ*pCiN� M=,�n��$$�4s �DQqrX�z �w�t�7q��Iߖ���;.�M�2C���S��EOP-?a9��爐�K��gW�_�+�!D��2cZA}ׅ���y� X'P(��`ų"d����pλA͑L>�l>���Oꈔ ��e��$_s�̭���LDi��@���u*Ӌ!^A��p�~(��T~�bK+�hn�w d2�c��^z��c	�b	�m�gB���a[⼦��D���]'D{�k$�@��1�n�Ng?Ψ
1q����NCu�˦;6q�-rM�?�]�(�3�fx �i�����%G�z��M�t
z׹�n�_r\�Tk`-q}ճQ�G*�`v�E>���Z�mw�%����_���h�i� y�%u���>�l�p�Ҽ+��D=dI���1D���
N��{O���5)���m�Pn��x�^6=i�L�/�Z]�F�v���t���E+���
C��M^H�Mԁi�J��/�c6pm�(F��Vc���=e�D��lS��`{NV��=I��
�����F��>��m(�
 ���aB_sG�l��!fLA�ɝ�^g����g�ݗ���u}I�Y�1 �B�Gy����д���ʪ��deНpO��O���،�p=�~�D�* �0���q�n���{��$�<�����9�.@��_��Ͻ�߹qe�t<����E(Rs�dGg,&bd-}F$Ә�!^䃟�r��&R��>��Z�w�m� ��0^���D,?��V�3�K�~]b�y \����<�d�G�:�_  澌X�A�2t�����{
6R`�:���,:�ZD���xҖ���X����=)��)�+�X�r��0K���*�޼Pr4�<��.�����;�&!�U�[OF�������S����O�b�!��GX�\����a�J��9�؝��Oy(�QƂ��+�8��l�]�J�c{-�=q	�]�`�ѭp�w��nR�2�,��'��L�� ���#(&�f�� ��^8_GPs��!CsN�˲M��m<��!��/
;P=,�~um�f�L�������T�2RtT�O���<�N�B���Qr.jA�L.kJ�	�Ϸ3���B�VЏ�H�OQ#�D�H=.��e���-��źH����V��|���P������H��Ԋ���vu����U�������Bє��a{��ؼ�Ĥ=�h=�s�F�ʌ�&v�U
���mH�ϖx��!A�(�G����|�ڳo��5 ���$�$��Ӂ/;R3I�%�v�+XO�Uࠌ�%���J�<�ZV�%m���)�H��<�ƾ#��d�D�6$�y�Ѧ85�'i��0�U���؍S,�5�Z!�0K�`��������L�&.1w���|��Ba�4k�`~��m.}��=mEFy��M�t���3��'�s��������;#�/�!#���>��M0`oq(�ߋ9�R�!�@��U�(A}��?��:Œ)���_/�m/M��4���E�����_/�4f�y�-��A�b��Ar�A[)���(qw��X�6���M/�R����%��]a��%B�}��舻���Q����b"�a�9$��Kf��j���˟����4��٘��<�����e6�\T/0.����Wקi����
M]Vo1:����M �<'�S>W�Eb�i���o���\ lrY�э%�h�Ru�c�a�/C���'ԣ�-JM�m��Sm:Ⱥ�!׷y���6�lJ���N��V+���;h<H�5�s,�����!'�0|B�ra%Ӣ�������%�;�<@��#��7�7O�������H��׋��7�fd�yfO���::]�I&ﴍ��?@,2���f.<R��J�4}�� )���X0X�dL�4N���]3�ݧr�η�?���O�������[8�ƵuUH9�FTy�	Ic׭z�(�6��<��'4�m�6~�� I�o1�7M�$Ie��p+ǂ�J���g>�Y:�jӖ������k��Z�$p�`��22�Β��T#o?{;1�bL@�� ���# ��u9�M=4R�?h�JM�Bm)�e���R���rЊ��:����1f�ik��������U�t��Aba����L W�VZ{��r��&�Q �F�L��_�'�����`��W6���zo�`$O?}Ӿ!.GI������T\U=^J��ӽ��jR��}�&���q&߾a��	\�eus�~ ��{��/�'�W�9�K���pם�Zz`��6�5he��w�xǩ0d�0��"l�NLғ��5.��LɘB�n*H����m�-����M9�ء�grs��n[�(����)��4#��yu�#���-�q���~��[wBT��`oN7橗�I�ep3�UO�r�0���
�����C���⭘J+~V�d�* S�ʟd�����w}�q������D��拨<��+rܼ|�Ed^3�Չ9ѵ^�CE|b�!u�e���Y ���kk���/)��X6�;��@���U����Ȼ*��a��aH[E�/Az�py�{?6�9�8���O�@�!uP ��ф�g�U�����o�SH�\������zU�����w^�����\����o]��{x�����D<I�񷏣�����|yә���Xv#��;�0�{P�o"ߏl�9�G�SR%[{ʘ�`2�m�e�A Фp�H�S+��TG����d��m���Q�&/L��<0N�#2S&�uDIx�����x��1I���0E���ӆ�!Ҳ�X�^U�'Ì���ӰFd����SYd��F�j���5n��w#x�t�Y��4���CÐ0�����g�i����C|D�U5�u� �˛���UJ㚔��#)s$tص��Y��Ѡ�7�ә��8T�r&�^M$;k]dN1ɜM�$2�x����Q��@Z�9�8�8��h"E�D�ܶG�X���ٍ�$�?PwX�%�����o�E(��kJ�8���i�Ҡ���'�4!�fA ��z}7x+-ŧ1@J��
%������)$��hm�O��C���l�<{� ���T��+�DU��F��z5�zA�����Ѥ����v6�I�Ovk�\h�::�Jqm`�~#z��";X�$06���-p��r��p��ԮtM?ijV�y���~Is0k�P�����J�Y���;W;�EU1W@�%E�*�g���j8�%�31��M �	z@�nxDt6y��v�u#=��2�RP�1Ҁ�8ɡ��[?�]���<�����إDo�0WW�g9l�To��
R�J�~C�^	h�"�GU�3qB۞=�x�n.ݚ`)�{Zt�I�����X��kv
��y|�U�(v�W��VP�?��.���%�%�}v��<��/㝶�u r��yr��M���>]}�^W�Ň���t�g,��ۄ���q�q�x�z�U>l��CHLm{_��}���.`ק���A��J�̖�#"�u�|]M��s.������,�9��{��"���+�#��/���m�R����4-�[ɭ�GQ� k|�;�pg����y�v���^��*z+2�ۈ>�G�"��X�חLH�ɖ3{�u��)�=�m��)�"�+��x������W���#]`�m*��%���?��i�ţ��u�I��Q�B���cjo�劔��vk��)Ң�n̵o6�=ci�����6�j����c��^�p��~����P���O!1�ݛ�3�5c������˛*�T}��8�B��}[����Jt�1?L�E�F�'���4�^������r >�����6�Y�WQM׫�Gz�7��g5G��t������|����V�ד�Mc�y��O��G��/��D*� �I�+��l�������?6��Ukww�D[�&,XC�s�LA`R�u�\E$Ӊ�ac�vT���BG$�A��l�8����%�L��"�ήML�P�
�k�5m��Fz��z�6����a_ ��D�v�C�F�	V�+&��md��Sq��"�PN-�~{Odm�>a
t�`_3���4S��.o}���+5��$s`�CGm��&[N<�D��3WM]���7�B����^���ꕰ�n���CıO�yj#���X���|0���I�E@xO"��#��ψ�[�����ujmXP��Y��o%H.�1��F�3p�K��ЛR������k��^��B ��}F�}���Y��w�~Ʃb�U�<�y������>�HY/�Z��Z��\
��|L�#���VbL��G:�h�r��p0���?w�iJ�� �B�_~�V��R���-��J�%�;������@,�H��aa�~+�	�kI �m5&��ߧ,�=�m��0������� �1�At 9�E�M� �"f�����DC���1�7H���	����vP� M�ѥ-}�� �:B�k��TG�d�*��M�h�Ә;/x���K!j�6q��ԭBlw��g߆����յ9����!h� %)^^(!�Up���i3���"���|'X�\Y�C�.NuM�~�1�^0n�� �,DH�Eg�����B�������ۈ��8s"W�_X���+gq5׭!�=d��o�;�AI��������<Z���hټg`9�`�OT1Y����A!��x��ȟ!1�@���$����yd)�B
g6�ҧl����a���g&�:�{ͪ�Q[�z��~G��B�G�{�'xͭCf�����$ �	���g�mz��Hg�(s�n%
�,��d<�m�l� �U�]�U�B�lΥ+�`UWC��\pM���K#����γֲe��3w�P4Oֱe�]e�G��ڜw	����Rz��G0J�.�x=���X3��.@rT���6�x�z�}〉)~�~BEP�f��V�GiIp�<����}c��\����R��+63k����h�ݯ�NC͘l�g�n@5�}P��l.}��'��TGM��w��jf�)\�>ő�M��v��&���.�v� 0�%æ���U��{�~*��:�ܠ���=�u&�
�,��i��ּ\��-�I�)��E����V����c.��he�O����+������`ӈ8��p%�{`d��il�I�K��p�Q�"C��d>��*?�4�J"��͖G��/��2g�EA��ē�`�%`P��+f�:S	�э襛}�+t�gNt�R=i��/�K�d�k�c_�D�0:%Y?��@�o@���lN]��(���2 ^g<�(��bf%�D��e8���ח�����BUݻ�R�8,6'�
_I�DH���B��hM��	%"���}���A!�J�u�a�(�[Qb���*�EjxT@y�XU�9��~��c_���ʚΥ����i����D�� ��zJ�z�����J�\�������~�t��&h��@&�����azv
�Y��Ϯ� �` ;�z�tٯ�i��,!�-�}�N�ŲQ��3)��K��"�y�6�Q�fc����X>�Ɣ�km¶�ﷲ	8 B��� ��m��M��A��)�C�L��gP��	�j�ű�R�SئG$~�#�=>��Ϝ��j|���L伈��D�Ɩg�S��t��yg���@^�&eH&g�H�+6Y��d\Emwy�l#d�`�B�k�D(s���	*/GĀ�N6 j�5��<���q�<D�0N۰K#�DN������
@������^��\]1��F���< ��26U����O���a�KU�7/�p�{i�OUx�L3l$�JA'H5GP�+Y�A��z�9�^�M%z�K�0j�'�(��MH��v�paK
���ʝ`�|�^� ���~�D�P�e���Z	޻X��Y޹�i�Xa`��Ds�m�X�B����Y�슪�f9����O�c�p+Z�9̨���eP-�:��S��V�t��>�FF�c�|��qg�k(�5x�@���PF��8O����s�o���y-�p�G>���f�R�A�!�~��b��$��V���{�����Cu��X� 6nY�������ַ�h&�����RH�L(Gܓ�VT����Y���)�+�e��	K_Y{Uq��1'K�3j+���E�ˁr>:�ҏ��������au0,�g��e ��{��?�g��ꭰژ�қy4dD7��e���H�{��:;߈�ݦ�8 ϿUNX ��c,�I(�����}��r�2Ԧ��F{w���Rb�=�%	�G�:m;Y��uE5V��ڛIқ+�������W'�*�z�Q$m%w�\��d38k4b7�۩�������ԉ[�ɘ��|x�v�o�G�~Eqw�J�+��o��t�p	�Б�;���l�����9�C�2c���D.�	�
- c���� Gq��
�v�&����K!3�P�*-=�z�Q����F��ى����8��H;�|����%UM�х
U��J��x���"�1ʗtq�����"b����)�h"��j��Vo�&�F�f�q�k�k%� ��<��W�{��q�gӲ֕͸���y"e����c���Gʄ�]��PjYG3�v�Дj[S�o�z�ߪ6x%É�*�"�|�yHX��ߒ��v{��T	�;d���nD��`�=/���Q�6S�:�ka�U*�E�#���?s[ER����-����Z�W��0%�X��l_�=�O�r�VF��^!�P5�A ٌ����ȉG.�6��:��j�8:}�V��s�F7@$u�Q���C_��Л�&WҀ;,C��;1�Ћ������IG�w!I��*�MX��ɞ�9޶�~5�C��,�&�y�`hW���Pnnє���O]&a��#%f���U��Q!���#4�Noj����Ḹ�׾�SQ@��I"�RS�Y��閕�)�;>�It�̂�Q����ɻ�N�4A��6��	�4��qt0�2�M+lS����y԰<���}�t;ҾV#�V��I�e���Y�t��y�|7�\;[gW���s�7���y|���&vYӵgTb��L��V_Vb�&n21���(�M�'"T�1�*�	�����ZC��e��J��:�ZŔ�3�OHT>	~�2������ww �� ��� ��������Ȅ�� b�_��ˣ�	�O����dUH6#��l -0��ff�0iH�w��0	���o���o��I�@�w��w��E�r�۝,��T֕���7|�`�J6k`� ���K:��������WL��-|T��ϙ�	�ߎ5�O���G2,��=��\��oz�S�4��`�W��xT��k�?�[�k�J>b�F�N��%�NQ��[	�z.I^b�s��.[[%=�\&r��M��6t�1��;�Ѿ�xv-�v�Y#%�h<�t�^���s�����skT5�C�=�����^���G��^(&=#g�����H�{��%pl$FuG�t��G��%h5���>�<:���hc�H.�kS9��&�}6�/����
��\��M?�ֶ�Z1�9��J��BT{PG�e��Tn��f\:����[ʁĹ�w�N��)H�9�ZWMx�3LmaL��Ouk�#��Pk�<�ϔ]' S���ͽ�+��/�ɝjЕ��R�e��{;*Ư9��+��"z�\{R�c���S��zf�!�X�Wp��^(�������c���dl�8 �Z��o37�g^�/&QoV�Eǝ�����ǔ�SԊ��y�kԕ��Z���<�(�e��{,���r�}��h���n�h�L�:5=��of���TÖUCsI��Y��
������mܱ������������(��}0�FS1��
����&��~޹�;	'���gh���N^�_�J�b%&E?���:��DVGa�i!�|�x�ȡ6��Q��ݣ��i�qs�� ؒ�C@� ��m��A�;�����ӕ��.�H��Jz>Q.]��戴6��ÁX�B ����Yfiƹ#î]�+�`��SL;���
�{暍bFT��������,-�P�И�V7���3�xA����fJ<��z�|��'���cQ Հ&M5��Kq��on%Ω�T�������>�`)~���*����}�⬁�W��"��/K�����
��
q�l���G�x]����ۀ���[�A�_7�GnЫLF��m�� K�䢲��x˰<����1bk�u��^���%�`��+f!+�� j� ,R�_�KA+�����O�2��z�ⴢq���w�G{@���*|��W���ˏ� �9uhk��$q� ��j�c|!���O��}�M�h�4@�{��ơ�����`�G\#[��IP�9tn�.�A�G�߻� ��l�,�z�U���Y���0cU�5�F=�e��U�h,֟^u�%,狁�kx^1>�!�݈�n���QC���KF�h��òY�5�E"�6����������.��8Q����,�5w}��ک@i3���$�*���9uq��J��$��W�[2�;�TЖ���K
�Q��������b�������$���w��C'��+,�lG�k�����\�(��*ZH'���(�|� iJ��0��e��W@`p�R�0�Ξ襍n������B�7`��;M����b�>�N�,VVY=���d��Y#,� [�;��?+��?��p�����+��%��4�DMc?�VSb��)�H�~X}�n�:F�qְi�� ����mа:d*�X�+"ϟ�-7�����}��0���'���;7>�����;�2��|��m��|�:\m�)�{"')�+q�t���V��H�52q�nPKo��Bl��r_�J[�l'y�mQiY�4���Ⅹ�of_�w*<!*�feZ���|�y�)Ẽ�i��fJJ���gƨ��5 ��Rv��