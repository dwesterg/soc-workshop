��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�@lEG��T?��B�^�*�w= (��s��ٰ�gC!���d��L��	 �!�����,����̂�(�=��@^���}{O���	*S_J��%,V��M(G�uպn��Sy�6Y�	`E7�/��1�܇(���S�(]DA�D���1�Q��Ӌ�pDQTS�%<�g����#��Y;p���鮲������WM���B��~u�6^�M@iV�����Z�ѳ��]��JVlźx\��N����������MB��h�w��(�F���WI�eq�!�kqYd��V��B�?晢��T���eT*!���)"�"�`�&^���;ڑ>�v�� �Ǝ�N�bOD�8�}Q_�c8MrJ.��������am�p|OFL��u �g�ᗉ�o]W�z<���!W^�HA��u�H-�ђ��T��%����{���k����Q����$��?��O&bʣ>�Сx��C��"B_����_M'���c�=��+�a%��a��~��ʍ�	 &�(DPN>(�4u����Zx|�q_"�i�� ��V�_u�f�>�P����:$�"��/����q.h���խ�}�m���Uu _[�=x�OH�����Vn��ګ�ͼ|R"`q[K�R��6��O���������:��Fvh�#c_��Ɂ�a-a�����/��cZ!�}�)���m�x�
�Om�	��Z�y}Ĩ��S�� r��6�_}?u�Vg��ٻ��3�s�ʋ�3�Vzy�WuNm�C���D?��`X]9#}?f[��y_c/��5���7CA��`�N�:��_���f;�paF�/��,�wҒQ��[@CH��E	}�&�@�-�+��BE�;�jՊ��ˮ.+b��I�;������	�V� �D�g�}K':L!T#�-���Ň�^v!~p>���� ���n�,�DܘpT�z������/�4Ѩc�a�4�EPȄ ���g�Q��2��]À?j�n���Dm��pk���J��_x%eҶ�w��b ���c�qSP���8��l��λ�p������Rj�J�I#I2��AB�#�$[��w��۶1��S�f�]��G�-Z2���!br�8��iGm��}��4@���R�&�^p����E�|JՐ�y��(lQv�?호���HN�!	7(C9��39����U2B�Cx�c�E�w�����O(�P�r��B_�gcV�# ����9���^��!��$���NTg'/R[-V|����v@c��J��L4L��,Y����=RjND=���|u$q�8Gdad�D�N<�g�y���%���sn^(���R�!��s��`<��]�7�������F��� ���Pf���E�p֥���x��b>_��=����qSۛ�tP��:��W16K
�ǯ�,%��$�@�yw �!�����b!�gS&(_�Ǹ F�o�}�I8:!����f����h�km���sPy-�>	�5 I��g�u�N64C-	�]��W��xn$H���?T�� p��!et�!�>��t�`[��D�-�im!^g讖�"<�\����T�I6X������������"�#ڊ	�)�e~l��2
D����:E?6��ga��
<������&��^	 � %�(��Z8s��5�q'z��;rs����	���'�B��MA�?\�ړ8(�%7���3������L�������@��xl��quu��H�KU�XHt^x%m����VRɫac�Ԭ�q|�bU�sl*;�~R0Kn0_f�<�w�]Y�B���U/I5U�R"��[�|�n��o�(��K�b/�f��s�C������.[n��##W�A@
6�&C��_@�{�횕�}�kp���[�B�՜_-$e��E@'��5��&�Xp���n�c���BE�]Z�#���(�~��1ռ�Y��y��w#}�ZL;KP�~=�+|��svj_��p���{j��1�n�b8Q��Q��b�zPe������e�Jg!��{���=a�فa�X3�\�[�;�D��{��37v�/eR�b�-U��L?uPGj&�58�{	s��7����7��>�� �B	O�XNR�H��I
�R���H{��A�hXJ�<:���
�E�-Bs;�	�+v�b ��Fe�4�f�S�}��K�ȜQd�5�j_��3.G�O>����m�������1�*��.�)�����R���@�a�S���*h`7����2��H��r�K�J��R ��购,HΤ�^ʛn%E\3���e�9�%Y�@^-��LT$�{��%��9|U�����w?�.�"l^�{N���f���f�F�*��b���,��Ne_�[��p(�Y��xʀ��o�sm���l"�W�33�/.�p<:K(�(����dϹ{��t��@޸ޙ;z���͓<��i*��$grQ� c��c�͠Dk���蠟bCUUSf~�.��2�ߪ�7��p��_���CW�r�H�R�ש��~��|1�^�t�t\��}z(��	��Ākˊ��}�~�u}ȍ���	�A��R�'�G�n��ѾġzҷV#�kH���i��RW�SwƝ� �>�i""$���HFb��Қ�Hq�|2��>L�s���pK\Y��s��hFW����/ �G��)ë�&>��!ق�[`I�|��)�2G5��s�v9��]�gK�þ8���J�z�.;�FM5[�!�!꺈�y���6�ɫ�O��؀2u`��
}	���wI�~�r�M��j��V�.}lx,I݄��$���#��xɊOJa�j�gЊU7G�1/+nSL�w�������}v��8����mw��~m,{-�Dn�5"a�'���O�S>���e4j�h�&��Wj%K�j=�Ij�U�R"�P�$��vϜ"���:N/���Y��O���l�-w�[����t�t	j�h�3���X��&�.�M�Q
sE�kØ�g�W�B���.��3V{x�K�u����e����N_���<`�U"�t1��I���]P�ɸW{�}��s��!K�� ����/a1�#�qpb�W�O����p����O��+?QY9�g�_��/J��}=۳p4��&X|]s��y�@�_�)�o�P�&\}�y�Wc�Š��Ӆ-[���Q�B��٘rR�S� Ⱥ}�..�/ZP͠�1䕇o���+GԒ�J6h`wV�Q?pyUƘF��v�Ġ�F����hyBPgĘ��_X��qf>������d���n9�[~��g`T�뀹���f��gV��,Q��O5.:T
A�Ȱ��X�')?	c�6|2ǲjiv�+��<C��g$&�(P]����(r(ϮKĜr��,�oƴ&�s�$�	��eA���R�O�5�_�A�ݘ�~�[�� �ٮ���>��#
�+���;�\[��e��!���]��;���8�xQ�ݝ8�MϚG;3|��A?��L�ji���|`�r[�����᡹ �����Q�]=e��QB�v�`�
�r ���<������?��d�QG���9�
�Uf�\�;��I�Χ��6:�-���[��たv
DR�(+R0�+�����%���ƶpgÔ��(��C�4ޕ�I�1�$��U�V�=8 AO���:�7�v_��9����-g#�*F���-�����9[V%c�lod������IV���wx�K%��;i��/�l�����;�4���dJ?�ӛ���,�#�������x��%y�6�F��=&\RH�P�̚'����ň!�]M�zl���Y���z��i��d��e�&��_b���~��s]bVOz�N�F��Ӕo�Ė��x/7%��U݀=�t{;Ұ�Y����Q[mN��8�=�����ʆ=-�W����{��	�7��|y�ן�_գ�Q�r��&�׬��46�O�7)�A}�ie˭O�<�E�,5�^'�kiY�m"脌������̿�س�O(����ݝ��	6��}���-�E�ǖL���ea^0o��PL���	���)�`�[��V&�p�\?�?E�d3;7a��$�W�-�P�C6:R�+(k!|~�r�+�/a�;����]�0��(�uxy�mg��NБ>x�'�����)�ҷ�j��/q<���Y��H ������^�pŁ�TTW�JM�%�~7q'b$T[��3�����<+oG��f�|?�T$�8ǉVǹ���L�z�H#��G�?_wR YL5o�gw釭*.�7�AبEEt���w1e>B��]�9���($#�ya?�}%kl)�ۄ�}��z�5c�u{:�#������?Ӓ=��h���,ґn@@G��߬�)�C	)���T��:$S���v�>F�V���!`jDT��UC������)�_�j�FfG �`��Ê	�b�R=$7���H��g�n��%�ð��=��>�y"t��n=�d#�,|�W ��]�kgm"5�	�������壧���;�M����x�d��<Wf��
o著ܱ��:(� uZp���^4*�0ǯ�}�wp��/�D���xP𜛭F	�x�/G+Տ�C��~^i�E_Y"��
��4�i�����xuq(Ω��o�*-�9���1����{wb�Q�E_o�Y5ڸ@r�D��s��-�:���ȭu�^-��櫪��>Ͷ�P_�:j+TOf6WB�|�9q��fqI?��л_����g�u�}�j>�!�@4�ں@�7z�Ivx���ƃS�}�]�sy�Jg����c�&��S��E-���	�``o��ƣ�?>9��%v�����F!|�R¡����ٲ�U�i��[ǐv�@���#r��ft��H�\�&��|����t'Q{@�VG|s��*�IDOp���d�5����3�7�Gz�"b���y�Ǉ��5`��a��.7_8����1���stL�I���߭,_�������A>#6�"qc�!���+r��qs_�F�k����Gk7qv��hј��y$���nK��נ�e�K����}׻��b�`��zI{��n�y�����Ϝ;)��m��f��\oi�F��^}�?���Ef VN-UIс(�+�?B��]�'�(7��@�͒lu3�yɥ�#�v_�(�ׇx@=~r>��K�c�_�;�T,4��쨹�x�7@��r0w��8�^!���z�`��w�q�S�[O[��!��������%n�7E�F�)�ʣ���8+ծ�x�GOܮ/����]��?���:��pv�'3	��_�v�A�o�-b��	�o�vL��j#:)
`t�����S�D_#qр��7I*�)k�K��@���X�$���`Ĝ����δ����;�{лMC*fPm�$��L�2L)�B�r!�z2%���K�.�s�_���!��͂�&��(�"�L�tHtַ�.Aԓȯ%/�nY�,�{�c���C������mN�EJq���Wڮ25����@_����'>�L��H��������jxM��Ik?���Vm�����xRYcD)d��S�7ҵ�V��T�J¸�e��c�lw�7 ��D|�$[^��%��S����ޏ�3�x��_�lx ��6��t�g��tBQ)}��f��U�n�~�����%�H�*�'�푡W�5��u��0��X0c[J�B�nd��G����%�������FPS�u���eJ�С�f=QB�;�oX�Ⱦ��p�T-��Ԝ�H/ȷ4
rx���{�p���m�o��ߵ]���<���Ȃ!�-nl�����W���p���x����d�Ri�}�N�n�\�!��G���ݤ|o��p�R"KR~]�'��{	��@��uy�b��zJ3tar��_�D���6'�.�ڎ�l�HT�˙^t0p=
�a�����fb�0��x7�Ο�L7��`����={�O�{8��%f˗`�/�Y������R���lP��lq�!-��,��˜x�d��m�(�P�$���K��W���g7�<���3x�R�KT��&�|���tP�a��*�ۿ>��JL��$@��o��<��}��ğw�	��Nm�� =źD/p�#I�,i������e����o@ǠJ��>oN�E���P�A�\�P�ΐ�f�\O��4��z���s^�=�ְY*ŴZ���P"�����f��b {4�� f�]����}�4���ђmc��c��ۦ��|bר�-u � ��I���Y�?u �W>���H�^	��x�@���*����hH���pTeT�,*��Z��ɏ�9JC��f����r����=`�*T��aP�<�"JߎZ����?���.MԫcFk�[,�AH"���ׅv]jޓ��/���3�����r���tނ�-�瘽��&7E��̀�:T ��.�nm��7�4��m����)<FUc��ǨD���JS!�Ɵ��x�(��#ah?ܜ���ᔼy�GA��_����"a��%n��;�%n����F�Mt@�	(ۉ�yML��0S&����Q���t�(�00Zu�E�iXE��,t��YD�8�W=�����O･9�􍄴@���x��N\7/�+ ���s�J3����e:��T�\SƢ�=�r5�g�L�$�!�Š�bI����gJ͙Ұ�h�
[C���ᩔvȉ�	���1�@1=7��jg�����Su��R|cO��`���~ot�qFޠ���/��{A}��5��&e��#��S$a�L��Z��B���zW�\\ �eRw8V$�M`����	������U�������/�B����l�CK{�N�C>o�}��h�{���2�i$�9�p�P�TQ#�a�3��)>�ڍ%��g�]B2���:��J�`������e�����
c~���MV�5�������]li_��IJTA�W}`�O+T�PݘՠŇ-�ߌ��3m�gPIT�]�)n��Ӵ٨oq@��4�����w�b�r.R�O�F�;$^�^;.02�pY~3���+#\1e�]x����S	lI�������<[k�{(4�
a	���M#�H�~H�7��V���B�KN�5ņ���R5\���w)?P\��27��Efqa=�x�f]=���ٌØ�G�}�s&%�Վ	���w�p�]Т�g�?�e퓏#<2���/�M~�t�K"��(�u�޼�7�=%*��^���"���I�X9��(1$���� ^x	�J�~a��[��S�܅Ʈ���	Z!`���%��.HK.��P*�1'9�	��'�rC�L^��!uu����sI�н���p!ǰ�c�{��c.�����['��b��ಟ�r��Wx�d��k'��o�uC�8�M� ���X�-�ѹ�W>�ju��C����oێ��V����Zߖ1Q�����1M%�y�]I�Ǐ?wגwƇ���g�%��xC
_�b�!�B��.�\c�v�r(���Tv����O=�X���BJ�ˢ�)#��l����������g��⾰�cꜩ�Ŋ�vN���;ϓ�X}��&J��UCיw1Q3��^�u2H�Yx��ᩚ���S��'�F@6C��{Yxk՘{��E2�|ve�(�;�ҫ?i�.�H������4�$��)�D�/B�����������7}�2���OZ���-0�L�jJ��)���GO����]bh=
�r��@_��vw����ِ����Л5/�7L<;�j���DtC����>�"]sX#g�+~Hp�!gϕ�~Z��i/d�1�}C��k���ګSr�R	�+,��.�g~~))���['�"�� <�e���)2��K��?��~˂J��N��`hLlL�Bw��[u6AC>n����D:���;��?�百1��&�V���6���'}3�����
s�ޖ�
��0��3/�][�)��>1jd�b,�)����jN�@`Fۄ����n�ul�m%���q�ӫ��P�{�����A�J+X����}��܋e6͇�c�];T��W�ns��2틝5U���8�D���4uz���"|-����ln
�0܏jK����B㝓!y�$�g��$�?��K\��</2/Ø�ڕ�4�p����/o)8�R��_�M�ot
�}̣q�k���y*��"�0�wu�U h��3E�{*�2��\{� �䑰��<�]A��=�?��Z�#�|���єO���L��`���3�kl%2��P�߹�=�A�Å%l�h�5���ZR:����|�-;F��X�b�F6�ג'0��i�e�������P\f�b�e1�����+&{��_;������c߉�4���)�Ug�]W������w�$,x��,���Z��˗K���Z��/��Q���5]�`���Z�L�5@'�[;�Mn�1��)�+CHL�E��CJ��94��,/���<E���1����'�#R.d�!�5PK��)�� �.Wƪi e�Kރ#�G�,(fm�sI�>�ֆ?��s,@e(g��J�`%��ϲ�ՔbKl4�`�]ER�bG�^Ƹf������]�ZS��6����V����Xm��wZd~��7�$�DK#����eLqKh���4@�MP�Z�k�r#�����H��G����Lp\�lY��탶�ӵxw%������t�7���BĂl�0ٮ��Q�F�2���P��?�ɔ��p�o!?OX��Vu U���ߢ U���ql��)b��rg���=8�Eg3U������M7��Z�Rx`���ffB'�M2�SD���'�� ��m��9�W< _���0�J@l�Bl˹���&*=���W#X��H_��̶瑈+��$ۼ�8��OZ$�0���0_�F��G1��t���/bĸȷlrN]��?��װ����o�Y/��Z�;&��1_<ͤ#HN�8�eդ�e�}���E%.������
 �Vnc;�_�7\;C��Oq���6m��<�S��l'A>�T�o��h��B0W�b��.x$��,��Ɍ�Ļ�YCיr����ݩ2l��Nm�h�r5i����TnkJ��Qe,�ɏ���-���\�At5<�NՁTLy�z�a?#ɰC;3c��f�$P���Ey�Ȭ_��P!C�9ܱb'�%ab`:�ǌ�������]��jj�J8'G;�#ښ�U��ǭ��b�,���,jaxH��:yM�#E~"NAU�V�g�Nu����E�<���1�V�׮��M���ӾA�H�ᶽd;BD��i� �-̉/��Gʿ7��9�^4��I���E���Rn龓+2O�DO�*T�K�*D�Ve�}��/t�
ӊZ<��xr2L;͒^^\�����o����/!�������CF\M��M9�%�Ŗ�d�i�A��y���x',��4'~�|KѶt֤�T9Ei���8/��VF�����;oa�&��Kdss��	� e�>v��mX�Z`��/����"1��1��[�;M���?J��(Q{����Z�����\tj�\Ȳsa�:�E�z�	��y�$ŕY��t�K)ٍ�����`�\[9� ��p7�C�d��YM���ZA�zp�����>I�1]ͣ��o�*��*�bR��B&�ewFE��wfV�����D3��әǉ1�&.䃁�\���}�:�S��b�������G����u�n�U �f�#��P�op���_�!�˶e5YO$�੢����yV[-�8i#^��+4I�Tr�&k��/�߃�o)ɭZ}o�a���%��8��o�
_�j���ၲ57~�^]�"j�V%����`{�J����Hf!�/H�|r�&so��u�xH�xg��e�{���P\�,.x�P����d�)<��HP1��\p*�]��W�0k�x��whL�n�����Ff�:60�>�e���dr/ZH�nKw+��j��`����w6�����i��P�c�����:�z��*�|�'9�|��f��\�V���
bх0�k�S�&|ߗd����
��:,��=D�������r@�{��J��$�y����˄�	���s�\���W��d�{�}��T�ˈR>�.F
����T���ֈ���Q��Sȕ� >��9}M���d�2�qu.���O�
�a_�N*i �S^��[��82%����Kv7|1��q�ȊΌ!g� �[By
�u�	q��x�����CL�@��k��FB���.u�U���� g�Z����A�Ic,Q˹�*3��'����?�󏌛�p���#gyH�p�l�b6^�`]�x�[�z��q���*5l��<��FG���<��Ӫo������c �a	�L��$8~��ȝ�v* ��P�wu1u�=6�?��|���P�Y�91O��ƿ��y���v�"}����\>ò����V�bϔ��C��LO�cmDyq�6BQ!d�l�(v��7>�Q����ǚ%�[1�>�
��d.���'�bB=E�*9	]B�E-������l�@l�����C2���4ĸM�8%@��k��öxu	/g�N��8�'-
��s�x�
�2��Q���!&�穕)��ӉͲ;��o�qB�?
K��(�"�����o��A魯,���:v�+;<�8�?�V�tܿ:�P�p��%+����n�����ZH���.r�T��d�Z?s�I��o��l�5�ϣ����������A���i���EՔ��Eq���g �!5�|��̖=6�ҿ���'/Z�`��N���Y�Z1�o��iZQ��Q�k���O{.�
���̀X��}.Y���%&Z�z�c��"x�87���W�
6L>L��'�fpo�[�S�f�$�ώ�Z?�+�؍x[�X�26�6cPp2��f����F����%D��r���HgL�\2�O�<b�ԝ4�Wf�bpN+�p�JU�8�F�w����=����.�*P�3.�%�q��k�CHW�I���c��w�	��⨼��3d�y�M���I�_]����$���(�i��-_n�2����h;|�� I�	��w%$���|��e-{��8BjEEA6+!�R��/V���������/ȅQ��kKg��L�wv��2�y\#�n��^GRn[|;N_L�D�(�_h��
��2�f�. q[7����-�UU��M&�����Q4ж]F���;u4lx�P��iL���"�0B�����z�5��}�;J���l�8�z�������$u����$����>F7ss���6��A��ɪ��d���R���F:_��S�fG�d=u��18���R�`n`�H
����>���:�U݄���ф �n�T���M��7�Ұx�ֹ��)�����r�LR"j�h.�Pε���G4C��N�V����L�#i�7e�}��bv��9�ۚ�S0�!�}�3"]�!���b�]���6x_����BqL4�4~�7I^��3�����:��.5����x��k���<����6P�J+@̂����C�v������/*u|�F�\��3it�d�/�D�����S����V��_l��Yߤ����dc����Eg�Zc�s��_΄E���d'(8�p]k��"�����n�x���n���R]�,�Q%u����B�B�8����Rw��h�)S�ì�ߊ�+ʋ(p��i:��g��;�-Cg&@��$H����ô���)'4�:V��O��	r��@�w�_���DA� ��B�f��p4�T��L�׽����5X\$E_�@���k2b�?�,A)�v;��g��'\(�S��N�ho��G ��=����x�=JT�Tv�Y����9Əjk��c�Ǧ��&&�p��c!��j!ɴ�Q�޼C-�
J���ҝNI�&���% 1�����߷TH8����;�q�NA�&�bڄfDE�]p�G��-�����.cB����`Q�&@��H��!; �U�X����y���x�qUl��v�LF+#`�3�k.W�Z��D'���m���F��i�eB*�b*j�3��i�w�:�S3~�bu@��j5I����V�1�"��+$N���&H��②�4�~G2X�@�>_��Dq7`*F�v�����0k$<�c�}Sw������ڮ�����o�%��W$��<���I@F�H��Ky�|̓��c��&�*)��V�#ғ����Jlm��Mnx�	�����m��y�1%*��\�|�g<��J܎l7J,�]�ܨ�z��C�I�����	�N���Q^�-�'UB��U��Ib��]�y���.�3����)B��Z��|�S�2��l�n���{�
���ҵ�BBυ����a���#�R�I3��V��~�>�/>)��^��	�J���B���'9��B�!ڸ�yԂ,�(�$I��#�:(���5��4vd-rW�J%��xof�����M�Q�L��U���Hq��Σ�v-j^��;�|0� -sw��}���f���`�o;���^j�H`T=X��u�X�,ʹTC���
�\HMqL��:�?��G�X[��@�g�W�64���֪F��GiΧی�iKс��	��9��<B����Jj����M�����Tn�,�2�D��)TR1'	+�6��ũ�*��V_0�
LL!+f�mv�f�K��j7l��7�E��\^ ����x���n��Hq�9o��"�f��t� U�	YxTjyj_L�a��En��3��p�b"ė�{$��0,�F&"�A#��.=��%-�`-� n�օ�0%�䅍�y-�!�{�Sh��H�^BZ�op/[�@������W9�y@@�`)���[ÆW�4�i9� &E����s�}}qo�?UMC#-�%�F(	�}iD0~pt4�\\��������zG�݃��g�n`(\�?u��
�\W�2��������QnB�r��(���ɯ\�3aa+�$6Oˇ�7��3�~�%�%G�>�D�\y�j���q�
*h���d�|L4YֽK���3�.g��,���o/�����Ĭ�)�+��g���!!�wbM���1(�����t�	J�2o���V Z�{���R�i09��B#�����0�l�o�5��m���{���CR�W���ھ1��!�+⍇�3���
T^���p?���oڻυ�6�N�Z�#9����x�Yq9�.�[��QB� �F�<�0r�M���c��dO3�k~R/PZZ0>��;�#��{+Gn�޷������3��!�&y�����C���c/7  �Rٍ:E��?��f�����G�G����_�5<E#4�Q����LO��8�^վY-ͬ.��^�!�*��e�~�*2\I��_D��=��}�S��qnB�Dh��QMdE���x�R���qU�+pu9<=D�h��;f�S����7���v��{�J�9��Nd����p��t���+�9^$腻M� a��S�p�v������N�[��uK�n{�鉟+�9-˸�\幏�W��p1|�x�`"����5��|5��E���"@MX	:E��9$�3�Dy��E�6�Fa%�~{
�K����TͩM{�2�y+�
���73�
��%_�D�S����9B�C}�8}ד1bx�����6�NVC��(�,{9rM��sq���|������&cG�A[�j^rn���<��ϼ����L'��霩��d���D}Y����kkT�"R�ycݟ��cC���8�}����ҥ���c
p��'��3�Ё�����ǧ���h���W;��0��7�]j�IAD;K�`���g>>, \����հؑB/}R���&'���T�N}��7S  R�
OX�p�A��M��L�~�ξ��e�钜	���L0��rԥ��h=g<hW7���8)̇�Ȥ�_猛�J#
�j/�Y���]�R���$�����K]������o\T��ܯ�3xz�p�Q�bօm��W7�x,�^��Ϛ\i�<F�q���'�ZwV����r��z�k%N1���񼥛�u* �iPcT��pn�e�1� 5��x�WךW-j"�C�����a7��8͖̬��t�H+~���� e��៳��/_P�/�����^S4� ��$��&��~�B�7��O/�O�Y�# .cw�m.^խo���X�-ɔ�%�اϊx�Y���:��wu��&�I�I6Tr8ەۨ��៘����T?
�X��I�Q�Ii�Z`?��HŔ��Eњ��P�R�����C�!���Y�>uT�?>�i����jj
��)؄(���1��d�D�f�����a���F�V�8�N^,>Š�n3��`Α�g$�J{��"R��e�Ӷd��⚬��b牏kQ���;[��1�z�Z�ކ,:��t��l���җ6�,&� B��
��oH�q'[V�`���i5�qg�/?ε�g���2W�c��h��[�*�ȌS��/E����?����h�> H1���=y�Q7�O~��:tf�n�\��L9�O:��.L*"x��[^U�ḧ�����=�q�m����"9pο<h�(���II��o��]��fw��9�O1��e���O<�<_]����Z;ʩ�zyT�T��Y^r⼏���T"@S�iX���Z�9;o����M�}�FY��0��!���s�CN%�߇����4O��c�|@�*�*����9�P7\��s�,_e^�B��#���	I����wYo@�%��<ө�&2Qg\���΃?6��|�9������ޑ\-#y����=��"A�X��Y�l[m-#��p76.cF��+.�I���.���Bм��㔦]*��.[�Ɔ����vc!��,�񰋖���������
����>UU�,�J� Z�6��!�2�[�$��VC~�O�V���4K�1xڀ̽��t�"߅0�bv���sdJ&u 7�����|~<�@?�'j�scC����b)���Sb�-`2Ծ����춺��s��:�~�f�(< rL�#(�JS����D��J�0.�����h���[�����\����ѧ�XB�-yt�F7�!����#d�y�[jg���X���s:u�n�/���o����s6%���D-��#ןSב��3����OQ۶�/�:gɺ'K�0x���S�G��-��Yz9�gAƻN��tx����]%sG�iZ�3�i��sM7�8�;�N�����[p)0����;���e��X���RV�҈��-�t�ϧ:=��J�`ME�~����}���'�g���!nI0=Y�$tU�a+��S�s�6�����ߍ��[�S�'�7q	�q���_"��J�ZMf3�]�:���EY���ͤ���m��k9d��x�?�Z�%B�mGr�T�f�K C�LD-:2����ݔD��D��L{�"�6X���?(�f�V{<���&�M����0.]�g�S&�Cz?,�}M��'�w�%�0
t󎬏�����c]A�-��1@9����G�y�b)�����M��y�a0���u���(U'ױ�i��F9lH$�4"�;��@�R���шoR�d@���p�6Č�����"���ghnVi\���Z��y�O<L�j
~>��hyдJ��A:K=�_Ѯ��`>�9Ya��s;���;�Qj��G4�]�r��4�R���d�T�އc��9�Q)�9��4����~�Y��Gړ�>mVN����W��-V �l�w:Ɇ��¯f�S�Mcݱ� xr�u�j�Lf��p�2��|��ˬ�߂�D=����U���R�`���p�G<�ʱ>�Z�=ً#��6|�@��[]�u��Pq�ɫ%����z���S�����[�燍�6�h�)�R�y��H&�Hp��Y�
�kJ����!��B�F����o�K'M��*`wʹߤJv�ƒ�
�B�2?�'ƀ�g�5�H�0Ϝ��c�B��Z�F�Zt�՝]��p�oF	��b��4�g�v��;xb����c O��2�q���� ��|����LK��=�g�z@.�1�묑�0�<+���^:���P��\>UI����r����֌ۓmsb������G(�G��IӭǄ7��d�Uu5�'�K�X��"F�z�C�;?g�X�fz���B �x�u1��锏�Nס��)=�=�N�ս�^O��Q�y^�[�{���z�����$�7��g�Fx�!�zsGC����Q?�F�3{�6��3���_g:���=}W���}6��>O/���>��ޒ��M?��&����ԣe�?9�W���z&T���b�RV�-�+��k��Dj���~P�šG�a��*f?�����|�iQ��jF��x-����l\9҄�;g�#a���9�}��P��\H?(fh�}�u�'�,i`4���]?Е�0�}�=u��ĢM�e(�1�=�,�[vh/�ޭ�K._�qȀ��@�
��D
��GG��R׏�����vS�G@�3�.�1����Ϣ����vS�"Mm�{�{�< ǿdm��a̗��3fҚ����i�
�<'�8�Y'UF^�
7d�^�B��^Q�}
\����L�g�5j�F�(�����i�'��%�3��|43#�:Ԋ��m����bL%֨�et�pFx�	�@�6�3�A�sO����&8��#F�������;6ݚͪ_��zUoR-O�F�SƂ��~��W6^	����'E�`��t�`��āYoR���ǉ::r�C}�_Ga+����Vj������&0PS�K)�W$���7�P��ӫ�����ð��˓3x��X	p��.-�Er`ߤ��L���n������#��y2I���Ô:�F�vN����&`	�u\s���!jR�!�1t�E�k�=��C�MЧ�ƍ�4:	O��/FU�; B�6���]���#���G��bw��X���w����z:h���w9�����wL�:@e��jt���p�,�`����|�m��z
��T�4H��oi����FѪk2���7/f��d�L��7m����ð�9����}��fҩi|�R�(�iS�.QH��:;D�a���:����w�Ύ�ۓ�����o�d����1t������$n �0��AP#�֎��h�\(-�qd�I�(���/�%�o�R���5Q�p��!����)�"qo��v�Tح��b.7��~#ZN߉��5��G�x��02����訨kF"�Y NZ�$�:G'����`D�`�j���+�Vs��G���^�߾kFw�IW5ga���x[�l�/��OW{ԛ�7뼈��I3�9�Ԃ�i���J길��U�Q�'9�%׶;�j( ��;�F�LsQh�jD*%	e2"�<��R��ʺ\�I,C�!���*���Y>���4�c��m��2e��*�\�\��J>�)�w=�����4��fz��:U����Rd������4�IH���k�!)�FyS����ICP݉n�L=�c�qG�=��Vm������ژ��5_�����&�:�O,�}��̙�r�T�l��[�s`VE�h���2)#D},�f���lۃ����v��߇�,��Xz�I5M�"*|Sj�'��������ԫ�2���%��E"�K��gi,��p�HhW�������}�)I��%T��g.	G�@Lmɪ����+E�G���(�Xd)R#�Q�ø ؓMts5 g$��̦���i? ��,+,p��id�+�� Ԧ}9�!�w�Κ�F.��"�iw�0u��W&h� �%�c����¸�ۧ�O|S��CN�(�r��KI���(��!l�W#�	�9�3��sdW�N��%�H:���ݓ㣲sؘW�R�Pv&g����"�C�;-R���囊,���zA�P��QgϹ��ҧcĲzan�%�����_9F�?@z6\�6��e~��Ķ9����<L"g�<D�5p�1m��\���^�_Q�մ�}���5;N�J�KV|�QÒa������ZUG7(���5h��ȱ9���hP0( �u��Y(rKn=�/����v+P)�6�$H����j(_��4�����III�$Xh��M�Ƶ��gKԎR������̤6�ůĽ8D������/"�D4C2���D�l�w�~樂���")�N:e�-���猠�]y��ϚTh��%)�?ln�y�딁�P�I������p��m�bP���,ʏG�ʰ�z*��0�)
����$O�%L����ܩlxDO�f�/ذ�	קB�-�;#�zM%¸<>{e|��e�f�����OPƥ��A���2ò*�z0Ől:�d�U�"�-x&߸pvn���yPu*��F	��qXA�̃�:èW�H���Q�si��^\���5���@�:%�GAri �'dJ���V� �+��م�gq�ם�8�;��CX�FO�ƕ���i�����g�3�et��+�g�ò�f-Κ��Q���x0+t�b�&�'�u�v��ȬA����Ź8�i�2]���"j��V�ZC~�l��[Y1�q�#?h�dAJ�?+@Ǟë��,���X}>4S��2��.��G����X#��SIf�/���Ku�	�^k :J��� �(J�'-�w?��v�R�\L3c7 �&Q����`|��ş��:q!��ąb�#���@Wֹ;��Wd�1��Tb����\��\����vjD���G[ȑ����U����O�2u�GG�.o��a�L_	F>�xzn��	�[3�k��.��y.�ڧ��Bʾ�w-- ��-�:O�x��3��hQ��B��exZV��!E�3��8gg1�i�(uL�J�7%�X�Hd-��0��XFٯr�%�P
,�d���);21��Q�[�>��"����LgNm�k]��ʀ���G�uk�>�Q�N�2De#�E���lO����Ȑ��M|>�rfYV�G5w��#�w����H��v]|�1��>�DAb�ڇ�(6�6>q�	W�&{��RMN���B��!j⎍�궬/xx٦o���ٯ�/u���/�R���6��yw�}y�*J�En?k���%�̔ﵣ):������$�{��ٹ˘�b��;<�!vy���,d�ή%�Q ������Pg|��ԕ�`!����}���ҭ�1C:ia�?(-���g&����3'w^\=���"��ǂ�xn�El�>���^/5����yd44�k�OBys�d	�g�7~�)B�GF�hJN��M� D��Kp�BJ�{�q4����|���?���2)���A��\�O9���O�s+�_��4�V6�Gi�M�]��e�m�7�I���8��~�R0�S����#s\kG�.�_X�Bk��ڟ���}�I���y�����|�k���|�;J�>��'i���֘�Mj�RN'C�1�v�Ճ�ٜ�)N�{ՒHC�42=�������bL����zwI�"b�dq����i�E-��`²;Q�����fTN!��Y�4G���d���]g�,N���f���y�2q_��d���`���~+�}��)�D\7�c�t������ �,�k�	�N�_%K}�q���R?�N���Z$a}��u�0�K�e��v��Q*�y:�����d��6�=��_���q3"�_���]����5����ki8����ߜ�7�d�h����\��2��V]r8LSݑ(�Gd~�u^����e����-�4SIJ������`-U�3T�b�� �84�������<�ǉ�8"�"&oͅ[�JH�I7zF�	�|s�\�`�$p���}��<(3�J���1�A�bg6����a��-}��+H�{�e�k��~���M��N��G�\���<ߣHu	2�a�p��a���ǥW���YZ<Q| ����m_K;�CGrW`� Ue�ց�JA5k��%E}ϐ�bp�v���}����#�%[��zJ�X��n[��="�5
�}5�IqZF�z�7N�mm��fpi����- �aGYt/�7$�"�����tZ	�
�D2���O=�[0��\����x��V�9qcP�	���=ȣb�l�S�ׇ�m�k�V�IO�pFb6^�s��9ͻ]��5��]a�rt��"�P+��w��!r#�U����q����D��g+u�.?�oUK���)��R�-Fa�j5�I�K�=U!�3ey�?g����J�b��NP�G!- �U��w�݁%�r2ݝ�e(\.�(ĭkFSo���?u'��QM���5-!��/aEȅI�H'�4G�xJ������٘�q9X�����Vt�#]�����(�x��[^[>skv��'+�>u���B����d_t���Q�;S���ɐ�n�\ƈ��j<�eS.!6�/ѡ4�A�	�5ߋ����68�D3��:P����	c#np'�OA}�����܎�
pj>2<6
FׇP&�z�L�0���p/m�9�cg9GZ�t��!�E+�� ������f�U��'���.ܾk�R�G�R_���Ȓ��޾���w���Es�~Usm�EؚL䠤=(�sf���k�7>,�K��C��<�M͘�^������i����X��1�����֭/��nl���D-IK����.V~v+�rMNW2�*ㅂU��{N��%���	8_z��/�8�c�.%D:k�H,�u����@҇׋�	�a|�� q�e��:3�4���_"�B꿬��`h���4����('�^X�bV�G���Mg�u%u�E����"�%8GG-ds�״�����a$`^B��j�k�q;iNAvA]	��Zuo��
�F���l���}�}���/z��R;�N�w,���1A"�3��-`�S�(���9�hXi�4h��a�i�ͨc�\�[�����u�m���hU�B)"��c׶��J >6d�K�r<����s����wϒ�,\�&:e'V H������A��^�6�����
���L19��{ 8z?"����>��(1� �5���w����`�1����55�����d��q|�s��3U��Ybf<vXS�1�>Sʡ��v�+��	s �7L#|Jc���<C,m�����1:��q|���۝T�~� ���^$���&�遷��p����B~�!�#mu[�J�tjj0�<]���,���Fylq<��3��O�#Go*z��/ =ß	�$j^�;2�c-�\	��Ŋ��{Vc#��-3�n�,���Q�F��qx�z��be��9`��Q|�ӣm#�0���x��Q�ޣi#�]s�6�2Z��Z�rG��4�W-z�Dϐ9�����Ã��ݮ�E�1��{oB����ԛ\�����dܻ��$;8�]� ��gW���If��]p���3�_s�H�ł�۔���k���ܦ��Dv��H`���%k85��*�������=M���yf��y������U��N�_�S��B��!΂�@���wv).��F(P���ί(���"�ȩrO�82O�>¢���'u��pxd���=R�OZ�gج��9�B�s��}8w&Xޜ��[H�,�3��e���)�#ix}a��K��"{��b;[��}�+m�}��I;�v�x'���RC-.���w�S���g��`��Ȓ���{yJb��hv�Fa�uZ/��=��_�����-��G�k��T�1��G&D�WE���l �	�к,�H5�ŀ����l�� T�z�9���B컧��&�{��kRO��-U-Ύ���d	�u@DT��fbY�Lj=B�.�e�kꉤq��$�9�����8.�Ƣ��]���5B�slU�V�e+��>,�Շ|>ǍN�,&'��,�&��,T��wG�F5�^:v���/P�����f��v����2rG��D9C�1z�#��	�7��w�T'3�L��4��ZH�\�����_���#�c��CPn6R��{~S"���<<,�e�9���և?г�v��-G;����j�c� �;�a.��/K�x��DY�@�zP�Nwv��T���Sّ���O��婽4a�]���L�N+�A�L�|�
:��bJ��2��B��"��P���7~�w��^`0wV-oz�}jK�KȀ��#�ӓ5!� ���p�u$ڿ#R���T��<HPz9Ey����3X*F{���t��)����n����#(������$��PYW�b^�Y�/]m)�F��?p�A���M70���$y,�����f�DŁ�M��5�%%B�L��ʊ��@cלگ�q�ҁ�J����Z6��?��c�Zehn�Z�(f�逩z/[��Nѱ�h)v;c!��^�� s��KF������`��hV��y�04�I�W.{�dΔr��B ��u�J�o�
�r���Ě��3�n�'L�t����a��zϱ���j9��p��!��Rpc�2N�QЁ��k�{#6 t�n�������p�j��-r�X���a�րı�ZT��5nMge��4,2�����O\.�9ȏ�HfLߤ�4ۘZv!~�N �ɩ!ֿT��E��#�3��]�o3�cy��1�]���u��	.<VI�ٵ�����7}�K�������_��\��w�?B�{�%�OI�$��|tޠ�L�}�9�O��A��9=^�0(�=�')����z�7p���s=�����S��r~��xh������Y�@����5�=垁ܑ��b�r7��9m�W$��]�Vǂ��R{�ʜi��2ф@ȋZ8}aY:n�|���<�뉪��2?�E��3�0�/��r�D����i(��զ�Q�4>�Y-:�uY�*�,X�gS�IeXZƜ�P�����=�ШX"؃�����W����Lc���4���ڭ���rr�����Y�����G$�G���^W6/�_��3"(d4��1�$v�*s�.�	σ��T��M�(cd㴪S_�1oµǇJ��R���������!��d�&�p.О,E���|
���2���0��}%��]�������V2���Ͷ7(�(����0��!�&}Y�I�#�ce$/�u���X�u���:(1��ZF΃���,`0E]l������q���g����P[ �,6�]{�Su`z�~�=LYq���D?U0��7��ފ�ѭ��^�S��
cKM�#>t��R���%�F��	�l���S�G<�S�G������m��妍���Xwk3�ɀ�l����H�8ޓͩ��gK�!�̛^�:<^�,/tC��r�yo+��a��w���p��3�-��ө4��/t�R���&�aUpS�*�j�΂�P&A�tK�%�ՆYzckn�:�i���!������o&�ʓ��{D���4�������c*� �@�-Kׅ}!m���Dz���1Ҥ7f=m>a��,;1=3{L{e�� �^?g�S����G��x>���!��dD��̏kVT�"d#������{^n����y6d����c�0