��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0q6 ��ܥ�̬/�-��!djΌb0vѭ�%�b͝&�^�u@�]���&���C��N-l�� ����E����T�]����Z�;�uN2Ґ����/�w7������8E	�Ҡ�w�|�����V��5`�M�|}INU�b셟�(�F�j(OŇ�j��7^^�%o�b�����fBQ:"A�o�l�/�2n9�2)�;�zg;` s����̧>e���d2(9�H��\�S̒�V�XfT5�����@ m�"�����sۈ� q�'+��P���ڴ�<R|[�5V@&:�L��'z̉�6l�f�ƒ���'������ܔ'V�؞~n�<x���>������r�ư�O�zR�:Y~Q���չD%y�(F�����(�����;�@��5����(�v>��5���x�5Xڇ��r����̋��W���[cy����
ǚ�˫��a+�1[��8�R��[����"qx�����_?·��r�R�ݡb䓯3�6�k��D��ۃ~q�:	�"pX�^�w�Ɓ|��A$���ר�q�B��/Ɍ���X��t���M��3��+\4(;6Yդ�nXb󕜋�T>���oj�;R�Ox�ޫ��7�L��_�M`������?�ƚs���6s_���Whv�I�^H��Ee�Fu_0 ��ENPv��F��8h���o��Z�0�R��J��,�v���Zbgm{���\:~�|��Tc(X�h�~5�R�G������B$ͷح揪{[KC�R���g��d��Nu���+3��]�-��g��G����e��|�<���Èd#Kn`�K"�cֺ̿?�,�f�:)I�<;�5�q6��
�l�~��=*�gzJV���ye$?�`o�e)�l�.���;�]'�:o�v��0Y���DN�
`�a���F�d�9��QH
�]͓�m2'&�^}��v㈜��ә��pRW.�#!�Ow���A�x�Уg>NӏƖ�I���e�D׽أ!��S�8�����
�5,qm;�S�1�V�j�L�+82<0^�;�*۴���o��)��`*�	�䴖c�;��v��d:)�z�P9���H��fy�A[.n�|c�;#��F��/T��<�b_ �{n���i�O�D�'���&���?�x�����7�ɇ�'���n��E�4|m�]�	gD��t�4��wk��(T�ǬB��0��!jIZiH"O�z�헢Ha���~@��f��Ex�' ��S���~6���j2�2��熰�Vj�3�l�q!F'��C�`k��p>�ڎ\��'dԚ挎�F�+��XW,�_j��K0��	8���&L]�P�3�$�ލ���j�*J����tH��<���ƶ����mj�/��`���D1����F`�[�؝5��������xw2^�De7hwk�O@ے���=�5yvr��_���^q:��M59T+a�L0sM)�A�'�ⳝ������"��?��i�a�.a��C n������+���N��0��Ք_<� ���贯μ��|�f�l���A�J��k��I��O��:մ���,���r�h?"��8/��2�pZ�3�ğ�11-�o{Xł��ЯJ�i�Ķ$����_xK�'�I&*|N�e�Ҽ���'��1�Jޣ~P���.���х�����1n����+I�vrW���H=�Ψk�IBqR��KQ�#�;kw�܊��\Y�8:L�@�F!�8V���ы��<�7�*t�do�*݀�������<⻢4���T�;mr���  �I�Cj��S��m9 _qφ5ʊ\�8� �h�nxo��2�h���܃`m�P\�{������BW��J�rT��ec9��+�d�m�9i>t��ͫ=�4qMn86�f�7�	Hߨ�6��%��!è���U0�C���y��-]g+��Pqc| k��q&(sA,��ԋꅖ�,����� ��<����9�w'�X�5Z�\g��C�m�zJMw��"���d��r2߯m{Be���-s1eR�5zA(�$�h��=*��9$a0ą>�������s��>��%�5	�)���"@�����8�;;�����@��0z���
�C}o?����_fk�PC4&߫scش�q�UX���$�L�#�b�0�f���\l�Sϙ�:���4Kc��yi\�[`��8(����:vM� 	G�Z�����-u^��eg�78~�j��`w�cy�҆Jw3�����Y�[N����"�M��穵<�P!Iˢ�b9��2,BS0H��N��5,�}]n�xlBg�5�vxl���ؐ.�]F�
�Ѓ(xx]�Ŷ�J��qʜݜ=��V�^�PُR;XV�C"(�$zw�-	�<9łQ�1NC�R��,�P>�-��)K,x:L��^�$�K�j�L�Oa3�����6�9"n�R��֬���SJ$ѥ��;s��d`]���O���\�@ z������[��k�z����+�
��˟[6B@XA4�Z_導��dN�,)��jE��qic��P�ڽ�rN%YLsIU�E�C��o�Z8%�D�01�����!@����Y�+�|},�qyS�<F,9Xz�-��6r��@A�!��K�Q�߳��Ĭ�OA2s������"�} ��jꔛz�z�~cj���kYCF�D�~�b�x�H��j�آ$�YW����W�&(l.��4OC��{�AJSA�Op�IE�����g�``��1�_��U����w��+e{a����a�x_������O�	��֋]8E�8�����ـ�)Z7YW ���Z�w�"�Ҧ�_���>�`Wv��:��53w�tu��*Zķ;}/TUlWb�DY�������VA���~�����M��۲�Ƣ�
�`��Eu�A���#�S,^�(q�bdyM�d�C�%XT'���[0��"D��5����9�_�|�Np��_�P�L祓�d��x�@9��_��ͪ�izb6*R��*]��H�VW��|�=�Ir1�1X�{��2�yu�+�	k����Ղs]�	��Gb��t��ޣ��t��<�f
9���_���v�S�30ے�'�n:�@xZ��$%m�Tb�{��gG��d�T��x�ּ`����Y�[�YG�ç&&��<�����|�@��2���� x�E��:O���ȓD�x�������e���C��{�����Q��ھ*7!�P&-HÚH��ö�M�a׮3"nS�J
�l�",Ӌ���*b�m��L�L/ո�5͈:�y��[���3��il
W�Ne�GEqK�c�X&i�����yQ�DE-\��s�s��`+���g��cDѓ]_0*K_3HW�q:ڐ�G��Q4�D��y xna*�fuǲ���&�B�kIt4�h4�US`m�,��1����32�7&��nr��HE(#�\x/��'Ͼ�R5yo|���pg�W���O\脻�
��0�8���Mg�)��_����~A�^~\kl���9o`���x�.p�#����, f��;�5UM*��P%������^Ikj �����ߋ=��2:��l���֗;��H����(j��A�KSRa4���*Y*ys�_.s�)�Qi���I\��ծp���,�^Uqz:�����W����h�v-Y�/��BkQ"���������F��W��O���g��f/֮+c@$E�I�.�X�NY]�P������n�?l��C���9���v)eM�/�9���>�#:��GJ�"큡���[�/���9 jEF��yA��)JM��D�����x�,Ž����`��Y���T�����1De�[dp}Yɰ����I�ˀ��s��&�ىB�!��ӏ¯*
�G���G�w@��^3�*��K(���~}�Z�N+���"A�D����� �Ny�"]Ǌ���"����z~�)%���a��4h�օb@v����BP2���	��M
�b��?�6D>�W�Z �9`#eҠ���w���Z�����M�KE!���W ������ɞ���p��O[�!�X�o�C5۲ɈU�����{>:��g�^�i�z�M��{l�a����m����2��r�cXPe�WF ��N�M����V��qo���A���nX�ά�0\z�1��l��m����z5��"dN�>0�RH�����e� �v� ��'"�9y�BXZl�eЉػ�v$J^� ��I�`o��<v�b�^-�w��k��Ex�e��t�;D��C�}��qVh�1�+����i3�mb�7}PC�<`�Rn&���<ڲ�\m���[^��~���U4m���v]�DO�zU�����ih��Y��_+a�߳&����v��PR+�:)�>&� �1ED�����ߒy;�cG��6Y�T鯟�!�u��n2�Ja!��3o�|\t�qӟ�\L�Ko-�gg�aOl���f��*�{�*Yӷ.�����6ڧ2�9/�	&��������o�
��C ,qt��zěcS�(�x\n=�4��f �e��%jGx|Dx�.�3������n�HĪ,
}���}ϱ�⽰�����2�2�����e��o���	,k������hF<�=[-�g�� oy`��5����q��Y��g��2� ��rT�T�/_@_�9NqA���h���������L5�(�N�
��N��yEs��Z�r*�A��P�2��er�'�B�����w+���m�4?�,ƚk�ib����<9/�k6�Xa���DC�(�"��t�<B�u��haW�B�C���F��Z�H`�����6Yt�Ʈb���������[�
A�����g\;Ǳ�O*�i�,�����	��e"u
�������V�5�,�9u=��z����<Q���,�1	%�4	�`��$H��V���Q�)P�C���oCڰ$�z�t}����g��ǽ/ח�%R�c�X-"�'x>{7��%���j,8A���Np�<�x1�q�u��z�LX+V�o��e=zz�Yl�o�K5(���W�����%��/ �W;3<����-�d̎��EeX����~H{�/M�{�Ok�
��ɲp��yi���%�4t@�f�L�jN�3/��!a�#/�ϛk�� ].��(�es  �'6hZdx�[�_n�(�F��C��Ȁ"���){��a�2,�U��`C,F�{�k��T0���|⏗���й�����"N)ڷ&�����GS<����Ĉ���w�%)�0���?,�4q��c�x��dʛ���jp���6��Y=R0���l�o0��q�}cʷ����eFl�Q�Ŭ2HQ�,m\�"���r��h6Zz�O���`Rͯ���~�@���L�i�Bg��M�j��}��*����Ƶ]����x*�"����� �7{��ƭr:�=:�6��v���
��u��<�L����/�%���}��\��8���#�Pc��!��������J��tv����@�Mレ���&h�eq=0�`�q\e���3�E���e��6?�|�ݨ���$�n�L�{�L��OC�kKȟG��#�n�s��Ӝo���7}g+M^L�f��mcZ�-��b��؉��Y�����6�Q��O�?([�D�K|�@'�$��G�xD��`��4��;0�GW��1S����������Jׄ�ҍ��Qb��W=��~͗�ܼ�>J(&��le�/���hN���D?.�[�a����,�&�.�NY���jq
�5p<T���Z���3&t�5�AYx�LfXu�#j!� M�i'�%GȜ����/���U�7h�4��u�{zݙ������R�	B<�m�L��{Z��p�߿�$�.V{�NAWq����nHM�[��#�\!'�L�CV��N��J[d����u$C~q�Ct�F���_�7�y�h����X�Q����;�I��� ���m&�(wJv6�xѝ����G,�O%�N�%̿n������F�j�X��XO��I|�,��Jci��щ�	PȞ�f�2FD�n��,W2��L�Mf��kP|��EC#w�
G1��S$\�+k�`$@8�������u�����ӻ��W��xߘ�x�i�I��fM����ԔYa������Ia>`<�-0 I>��iH�RR'�����kEh�,����@�n��$V�!���q���|��>�l�[vm�>���/�u":<��	��k?`+��΋aj���&!c΃Q
*�!ʞ/<����$��P~���KL�L%����H҇�'+"d>��>7�^4�٘���d� :��L��˜1�(�?c��<E8��B�}xZu��71���n �v��{	IJYΠ�Q���)V�y:�Ce~