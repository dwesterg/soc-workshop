��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv MCই,�i��������^�xuC���^�	��g���|0�P��짆���N*i?�&���h��x2r�ZS3����L�뵬"�I��x/���uB��XB��\l�s�	�k�ڂN�d׵�"�'��4	��X�� �x�<�	�����ߙm]�bM5#[0����K�	.�d�;��*&z��gz�:�i��!tFr%����?$�,_ ��Ƙ����(��cV�W�>���A�"iպ��!?=��M)[�;�C#��oF"�5~&���2��R�,��a|Q�뺍;6��~��uWjbh:%Lt3�E},��y�ض�Of���9�u��j���Ѷ�{�hԝxĢmK�Y���Yά�#`��q8��=� �S�޽&���|׶o���sp�v�=��Kh�%~�����7y��S�e�h�2�'x읽1γl5��e�����M���[�YB�8�ɿrFa� M�2m흹k(�6��~Q��t��O^t^U����D��oYkLh�Њ�E��'�ۄ�G��{�~��&t��a��ĉ�(��b���kF?9)�z�Ǎ���N���%a������I��D�n�V����>�om��D���2���n[�i�݊��Zz���]*=Y�0�	
��Y=�ˉ��4���7iw��*t!=��#�{�;(Z�Af@A�+�N�r���s����K���r��Ύy���C�y���Vf��UNg�!�{Z\�t��:�Y����ä�'a�ܿ��G�o�i���y,���ƕ�d�Й&b:�+A&���2)�:9|�������QP��0l�>_�;�iۮ(�i3Z�~eW�G*��b2���z��/��X�X`}��e��¢��LN���G�e<Y�3��A���:IG���柤i���a�<TY7 ��1����d�h�+8��2��"�J�`!�aFeS)D�4NT��S�*�(m!娄���$��'m��A�_D�`�����z��K�X�	B"U�ƺ��en�L���Sw�ϷQV6�b��v3�[�DI�jݙ���\VM��	G�/�55q�&Iě!�p|w�LWw��2�E'6%��ѕ)ts���?(��ÄAЫ��&3�ǆ�*�~��&�]�����s��T�Hyϫ?7~����LU`f���Ŭ��f����v��E�>!bj�<t���c��ep��l�T�LTa0�o刚�c�J3�:R���WTgN���^/�(�^ ��V��4��3i(D��\�NA�ߓ'�p�_�A*��J|��_���;�]3ԉ�@��Ҋ�sq�,Ѓ��DjH�l�y�ܤ~��&P��j������1}j���ZY�{��*��s|�n��&���!��2�,�~5=k@����Ee��v;?�&�����@5���~U��v6�[e��m����'O$[��l?�鷁s�~��!#I��">)�|�@q��rug��'����	�n>�.k޸������A��jmM���Wh�t���+���)��AP�	��a���E�q����p�m>�?eh�L�)���L|�,惛_3�'}���#S�Zg@�nuϴ�j��P{�Qώ���$�=�o8���#��^�Xn���{�:�0AD������S����e��K<��gك#��Xrg�^�S{�܅��H{E�]H��6�\L�v����,J�b~VN-*S�z�1�('͢��(sӸ�����s/���Ė.�&��Wc���'�/4�M�B�H��!�� �V�K�9�H��6$���~���,9e-���Ո 4�~�Qۭ���F (�?C*�	߇]�5z��+D�F���_҉@즜J��n9<JU\��>w���=9/�K����C:�t>#g$�#�W����9Z_x��=�kE��kM2�W���u�N�b7���/��X΍��Y�$��,�GV�)}*�9��LV�R��}��Fd0��7�x���~�������+��{G@���?�����`P�C��mw	al�7��7�nE�~w�v�Z*����u�u#F:D�������ʭcJVk&�@��dX4��i_(����s�8]�f_��Z��z�;r8��C�dImD��=��׶Lh�2����Ĝ�Թ��@������H�נ��XC��x~�,����SI��/Ȗx��O����e� /�R*0)�N��Vz��U��v����8����Y�����zJ'��f��#�H"��/�4��a�n�>�������d�#�=dO�76���`&*��2�O��i��M��7�֥�N{B������+W��6�'s[���6]-Ñ�����!X/�*�K�!����a.7�0J�n�^2?�<0��| c2�{{xɹ_��'@� #7c�nT����f��p������p~8o���'!�hr 
a���!oE9a���'p�|T���KW��s$���βWv�F��a-O5�L�����(@�>�8��(N�y���� �
� ��<�/������I�x�@�M+q����}����������ΛR%���^L��$J3�z-�ߵ����UυJ���?�	�#މ�Y�$���?�S�ǖ�Yh	8��k%��YUӆcW\�-�H��ӁM^r��ê�{4���*)��vy��i玔WM	��"ߒDG����h`2R��Z�Ѹ������fpGГH�Eo1�p-���7�[�@��hJ·=k:K������g�
�h$!�xt\��r�4��*P�Vy���jBYxR#eX�"���g�%'����ț5<�|싂
֨�]?VF2|4�L�l5Y�	5�6F�e�~辻��<��>ԓ/|���{/�v�t��A2�#��+u�Q��N耜R�m`�A'Pl�|����f�+ ���;.��`�ga���V�M���UI,5xT%�;A��um�����I�6���ץA08�T�/.�<E��9�����%�� B�~���T����\�f�>{k(�UPN*��Y/U�RL��X<M�z�B��CD.�LǏ�
8{^8ǀ��>���!/�w, ��k�
�*G�	����Sx�ކ�W0?bH��fm�B��X�'�ѩ�Ө]���J�����j%?0�_b���N̢�+�6CC����g�{��9<�`�+W{,��$2ApY�3�#����K�0,�N��8d��1�-'�]	�kDJiU��T�L���=:�:$ȥ�����gg@u�__�W�/���Щ�I��Rii`y��&k��j���fafo^Gi�;X=Q��z��nrT�p�O�ݩ�{.a�H�����FY#�|��Sd��(���;��ֶG���x��ɟ��j��6o�+��W@�!���o��"Y��Zk�Α�̴�~��X5�P�Ӭ�u�����
0�Z.����Y�kaR7>�=q�А\h�Yk���D�w���4 ��r
&]֏Gq$�Zh�n�!�'Bt���U���D��D!�
0�`l�T�)yכ��w��W���7��?��GO�)��5���1Ҝ�8���T0�z���:b��iE*9�����G��gI�rnj4�y�	|�^��9��x���G��T��\�����o����Q?8:x'oX�D�K�8c����R�9�CE�e�	�3�ZJ��%ж�  l�#������?�1嫩���Z7��"�R�!���┖.��&�M�$���@sު� ����_�>*��R��gK��8u6](���5AW�e��6��l
`�0uUe���#e�u(4��#���0f�n�6p2n�c�ˠ�\��<�Bo0���Q�Uz�k���u�Z�����,��=B~,��j A� m�E��d�@;�� �f�o��h�2��%���Mg��qP�,��w�w�5���z�z��Y/"��6+���Lnco #�ٷޫ�*&�Jho>�I�=_&�G�A�t��
�	�34�WS�*W~�����z�W�x��mKn�'�~v��5�A�)"w��s���y�'Ξ䡼���B���R�|t8@y�͈��_��ڛ�nBO�c�Z���׺�-�=k�n�o¶xLr��m�P��z�e����<�����p"�"�r��`��S�����Y t�x�A�G4��+Ŏ���/Xk�y�e=����_������d�Up�"�Nܹ��B�<�7~\� M�8����*&��Y�8c����#v6������ͻ��:�e�z�1¿�x���r5�P���)�p5���T����*�ċ_A�x����#D��W��$�IN�?��Vh����B�f�����l<��m�E��|[)Q�th��V&�L"�W��3��ɱ:�}�h|L��v�i�rd����"�`��\wZܗz�Z��Q�1�nt�����GE�V/�ʺ>���sS_pD�����c/%l0��&Ǚ� ����,��5Zl��mm��7\LXV|Q��~�V�	'��:2�?+8G����N����އ4VPTj	�}��-}6s{T����E��F>U����p���JM�
���8^~���[LP���W�zoe3ʕ'p���x�z=�r�E2C��%VC9�dZ�ţa��۳�lG�	#� �MC�T��+���=.��X�*I���Lp��4�W)^��J��d,�L����\$�h�ֺB��=Cҏ������o�8��#L
UNG&2Զ7?�*ҽ�T`�4����C����P=��s6����ŋM4�P�E���;e�?��Hb��|>�]E4(��'��'��v~��V���EY�o'$�����}��Q*콮p��g����Uv|кV.���`��$�P�ƴ����>�l2=�7�s�&R��+Ð)��ݴvEE��A �c�{����
��+v����g��i�i���osC7G�7�vTd�`Z 7���� ]M.��`������1P�͆b ��͢8eZH�e(,r����z���	)ħױ���\ݼ��_�J��a�P����fǃ���+��Ϊ���Ob���t"�{�����2���9�a;GI������z���[�Yb���nl�_���Jo�1��%u�mY��#W��#/�s�,\ǋ=�f���"*�W���Ό-�&6��cX8��v�"�k���`۰���-�Z8;�g��hhW���Z�Ш۳�G9hoP�U�:�Kg|�f�fi���p��59D���tI�� Tχ5`��޶,��ߋ�2h僮T�$d��b�h" 뀚j�A]b��Wױ��|o�#�~��$Z�����UPkp�]�ve�J[�Nו���_��m�
�+c���*i���K��B����~D�����J�А������y�'V�����;U��'m2kߺ�P�CL>w-'�T��Z�F�ҁ��k�r�v�Q����e��sj����RL�}��ĺB�L��tG]��2�p��N���H4\��P�ʨ�c������'b�ef9q����-eu����^T^�9��JM�F�*h�:���'��";>d��嵗wyPx��c�Ω�3[ʺ��c˧uhx"d�F�h�a���<�蚫�� w$^�A]!�M*W�F�;|Ӻ��Z�'�Isx��ľ89��4 C��C���<��r۔��1�������$�k��( +#�<�o����X�� ���DQ��������#q��TxN�c3���ȍ%�J��<dvxf���SKwD߸4�UڅC�.?���-c::P����y`�M
Q�k�@=c[q�1ČVK�1�q%4���}r�D�T�jG�?]L�r���%�c8�M�V,�g3z�~o�^�@�{K��7*K�gl�-F.�&�G%P-Z���Y&��j_9����ƣDZ�k�e@��̛L[c9+*��@��A�����]�k��f.�ѡ�:�d]����k�
�4C���jqu��*������ͺ�h�ߔ�0�ǈJ��3�ڷ��K6�J~�I$S6����됙�1H�m�z�q�1����O�u܈�O2�T:��Bڥ5Lz��˥���d�w�{��*��k���d�Ҝ�@G�<.��A��]�B;���&o�-¢��˴��}L�!1=�1Nޝtvyj��c�]��:)���v�i�b ��b�އ��-�7��aGyz��z�Er�r��򲻰v���]E�ꕦ��$��:2���EO�e��t,Y�:���r�D�C�
3��ʋ��o��9��Yr�KZ�]x+�����K�d�v��`-��%��eE��r�QIS�������X�+�LԾ����Z`� �G�n�+C��`����Y�k�B Us�K�(:�
g�#�<�V�	J� &g>l5q�bY\�_fڐ*&�d�Qn�Q�e�W�:n����x� ���}P�a�;Ւ��l"P(d�N
PR���>j��(�����4�6y\�j��qKn�ɽf!�)�in��i?L�����ȩ<�F��\;�.�h���d��f���@(U���P����S��cO��:����|�Eּҷ�l�C��;h:�k���W��R��P38��%��;��3�A��m9n�+S�Ľ8�&dG���;BCF�4
��f03k;ȩ«�� Q�x){�u
-�,�!`�J�Q�g�����Ӆ�M�=�&�ˑ�=���f�	>ŷ�)��n��+
bc�/�=�st��qC�$�%���yy��y(z�龦I#^�K�a��~������~^���>��-I�LU����F)��VN�sQP�'��eP244&xOրP�j ��΋_ekjT^Cux�X��S�pى��ݯ��n!D��5i�"���xz������C��@8��5�Z�X7�AW�b�=�|�gU!��?���Ħ�����yή�9HR�����!]i��EԌ��;������ϸ����GE�O ���˄�bm�$YZ?B�R4!��R�H{Y�$��������h�K������C�XksH?�'�L�)d���b�f���E����j�[�8Z�����#� ������mI*P����;�=5���_�-�AC"V��[&v�&y�4���!�;�����m���>��*fꗫ��V��N ;lM�����������N�-1�s�x5zx�L�Lm[���Y�ƹ�5n�>+��Ж,.�mD/�e����f��}��m(0����t�O;���h�?�$�y��&%W$�jH��'�d��Ѡ:D��=ѓ}�.W�DQ�e��:�w��f�\�%�{苪��'|%����×�<q%��yw`��`8�+�c�K�n��~���A֌R�iZSʈ,���e�#
��kmr���v���)����Qi�F�e��鷘���1�f�bݕdMj>��Ga��6�]u�p��8�F_0�׆g1�>��-��9l�U��
Tc{��q ���"K�?��9�u�m�{�&7٩:�v�O�x�hH������������̘�^�Vވ����u���6�I�Q��O�ЬȒ��p�j���se�Zb����a�E����K�˗�D�ؗ!�6S+��Pe(�VP�MN���C�|���V��#�)��(6�w�4B���S���ը�����W�>3�h��.F*C�5ȅ#j&#X��,#m��ɲC#
��=�d]%���E(�o���EW�
�)�>�3������Ĕy�yM����V*^݅W@�{*���,��	6�!B�(���E�l9�4�x�ݰ��D� ^�Z����8j���7"�~���)���'�]1IB#�_Wv�}xm���m�~�!f���z!���x�D��� �8��>�P��d,��=���u��&���*A����H���˻����r.���j�EQ	����XO���[�J��-�g���a�x �f��9��i���pr�94GP>�9�����\�_g��Z��Kh��X�����7�%��{_Ւ��Ɬ,����՟Y]K�9e��H��+����u���G+|�n�`�.�@J�}�
%���<�.���]��B���׺*;�+"|oW�$�	����(���ё���-���E�����C@��!���'��%:]���q�j��Q5�i��^Pi�����&(t�>Uj�ٞ�T�%?�W���E��.�+���
+���o���j*��.�\��U�b!������Y˩!�f
'8��q�<�v��x�e��\G�Vq��*)�u��d�>5��$&
���t0�^��Ψ�G��;|���|�����r#b�o�Y�R0G˱0��B�c1�vA++(�'I�G��(H����
�_�	��i�p��B��̌x?��D��(z���c��-hZ�!GE"m�w=gD�`�0^���T���:
�sAJ�% {nM�>b�˛X�N�c�l��f$K��hd�$M�?�ۿ�.��5ף�ESzЧ��oKh:��Ln@�����z=�*K��x�������q,���B�߶G2��G��hLH�P�����$���I��]
�Ldt�}��X<�kV����?"�<�m��<�~��F��5G��^H��p�Tr��ɪ���WK�˂,�
����[�)�,�0y��K�����f!5@�K�F	�YɈ��f��'t��&Z���2��(T�#wZ�F�&B�8A��?�n����������5�L��O_��옖<�vY"���1���F���P%�N�0R�A�w�'s»�g��΁Х֟�y_@1[�o�0��C��Tz/at��ߊ�����
2����吏ХlJDe)��W���$�d��&�����=���z� ���T���wq�C`��P� ٯ��n�u�<W��&�����_y��P�|�א#W`s�V���}k�m�*^�	z����*��m�\d��=h���.�[�t��/�T�1͝b����l#����F��z�I�F�<I&[IMߎY.Od���|T?r�N �eoY!�h��r��R%UҐ����V^��T����R;�6�8�4��9��g
��~ͧ�\ރ��5<c�qH�5�B;�pv�I�,Sh/_ϵ08��(X(*0O�׊�Y}���4��Y홬��ap�H�^|{��E
�@�t�*��,�T7(�$Q#X��Q�/�T�-9��$A�o���� �vc}
(yFuAy;P�n����(j�X%�N���R��7����<�@�l7�1� ��#�ܙ[����Cyn�AҀ�]o�z��UP% �����أ���N??����"�^V�xrP�uGh�n�eV�BrK����>|ĉ����7��O���%@|������7}G�0�J�fV9|Rt�=:ntC�ȣ��@�3w0���-�>�#���ȇ|���Xi�	&�劂���$�ߩ=���K�.�J4:8.#�Uژ��8��=�Ψ5��� T�Q1qH�,��^P�Jj!Q�3�O�a�7��R��O!��#/�^�����V�}���f�F�Q&�h9��0�g`\<'�d��Сus�HzM���M�f�i���&8�/�$@�	��8[?�5��B�z�Ҳw��^�4%dD�����i�������J -�"���1���%3d�ޏ��w5�J	���qGxW���~�ϥ�ׅ�lY���J�<�� -d-����e�����e������a{_�^#�:�E�	�9)"��b)�&�py�f&�f�3׀�w!���(�����Ą�{�4TS�,�KP�'�z$������o��ʡ����8q�mo����ݝJ���2��͋s�]���Y�ƺ��)�`us$�a�0HM(��%�)"��Z׬�X�Mi�V�́"o��e��f�l
S��4�ۜr�V�Ks�;����7�%����P�M��7Ǔ�!lхp��8�������H�{���i;�jr�ީO�	�Jb�X�1��,��Mт������Hs�AT����G�a~B�:�P�ua�#�F+�K��e�h��T��xf�M;C��j'��ؖ��x�vp�B��������n��؂f`�"�s%Ֆ�y9C���_�}�xX��eV �ޚ����P�Nd�t�AA�2�:�Ԙ�!Y�f�V4��GҊ�=5��J���r��[84�9���c�cSƾ�I�{|�$��3��m5J��X�C���:��sW٢���æ���ފǒ�6�~�=��u�q(>'��$a9Ȋȹ����[��>��Il�E&w�W~֐1.7R~���k,8�S��WJ��[O)�ǫ̅X�nC��ȝ���ߤ���i�H�yy����/4�ЬNS����a�]�S64d��L�x �6�pg���()e�5��[��-lǢsO]�
�*�E���2$� ���X�D��P�6�<�.��R���o#١�$I���ߤ��L���VEk�`�Tq����FC����Kp��ǵ��d'�+��9�v�@+LZ�ټ�,8�Gv��`��Ҷ�Q&�X�8M����V�/6���{W�ͺ��-���aK!!���Rݹ�m��E�2��}���M�Q7s���,���e���cɭI.����Za�/ܬ�Bh'˨��U%�)�c0�H7� 
�W��n�~IҭXY��%Ш�*��Q@ޯ�`q����r��a��G\kT_h_�m_�_d@	DT�2��W��L0֢K����-�f��Q�,=@��ca�Ps��U輔�a�ό����w�8)S�E��������h���CN�^0�\Q�',�� u������G)���Ws��s 撑S�R��a����x���`��hZ�O��нa<f���x����+�<_�ČH1����kA� ��K�E43W�!Um�Q���ςI�qc�2��7��4V�(4T�c_N^�u��ɈaD┼o��^Bٯ$�0S���x�S�q$������P�`wcx`�T�+xn,x���JŌ��H�
{��B<���0��\�8͐�I��.�P�h- ��B/6� ���~s��T�ܻ�ޟP�~���4��X�b4�&�mH?gC!`��h����9���Э6p��1��_b��	qP�Z�4{5��%���N�u-Q�5�帿S8������}N��.�Ns�
���h�|�%b��v<B���
�q���+gm�Dw;
U6�r�3��:n�JD�QH�(oْ� )c��#a����edJ�*a����r%��ŪL�ǧ�TM*���D?�_�}^ou��լ� ߟ���J"t��UEYv\ݸ�^6NmLt�����K����xI7wc��3�e����w�ws\�7��J�UG:�t\<.�%y��ou[I�h�R���r�ѱ^�ǯ����J��#d�"�����?����N�]A�[|t�᫸[����z���p!�Hzθ_Ȝq��E?#t5�b����Ss!��.��YY'0k����"&Z�\b���h~��J�k����'����%_��p3G=£X7�`{�(�ōBTI]Yf�Ud���D?W�ز�ո�9'�ʯ���3���)�Ot^�g���ǋfv���MbȦu�� �}�	�LU
w��H�wQ�gZk�&��0��9&�mXP@����FUH�XR &s���Ms>VBw�׺~E�:�5#�N,�v�����>����|���N�}�.�"����?˲��	��[�Zkc3;��˵>���T�bX�;e/�f�=:��u�U�G����i�.}�H�m��e8���(5^���JNSͧ�<I��n������Q�1��tj����
 ��̒jؤCS%`�&d3���t��C�KV�����'��Ug�#I&�7qi6~"T����Ѭ��i��[�W�
g9i���O�|x�2�\��/+\�	v�K����jFE�����L1����뺠&(J�s�M	�QL��A0�����\;E�I��nl>�y9o	9��j����/ ���c`r�s��>R����t��ؽ)��R��o���Ԍ��k���亂��r���H[��S�NG�T0������/�^�/���K��Є}�Ojέ�e��8���|�׳�����>K��
>q�9Eo��{n4��&^	� E��(�F��Q�s�_��YB����x���jz��Ĝ�K�q��<����}	�~w ��O�����y�O��$B�Σ.F�t��K�GT���(IQ�W��W�y~vށ[#]V�P��"��rt����)���r�!�<	���������� ��7o�� ��*L���a��0���7�]�N�����ځf��'�?p�jf�T���%��r�K~p����k4�N§ �(c���RW,��N_F�b�E�>joPb�uV��1w,����u3��œ"Vt� Y�k���bU��@c��K��y�:�F�����5fT���i���R�wAlsF�*M>.+����k�P^��$��R�� �J�%�&o�'Z=�|t����T�ڐ���V�J��z�f��K
k����>;�A��+Ń���OS���Gpv"|E�y=lu4@�%:���`�*��0��� .�sI�J���8��?�e�#w@���ܗ����pN+!�Ǭ��|%�:S�ϋm���$;��5�ɘ����J���<�#���/Q��[�Հ�{����<��'	2�qd^�u�ȹ*������g�����'����^]<��+����(�����A%kS\dc�>�f�o���^�n���g	�BR�꺈�C�(��\j���A=��,���.؊��6Q�K��p�D�^x�\��k@�)��J���V7�4(ΏA�.���^)f�y��<�����,'3e�����G��{f���[�O���?���\�xyF\�������� �g�W�	B����nw�Eذ������.ի�5o�X�~��Be�t�s�7�@͖f�`n�����;�����vB��A٫���Ԡ�.v�Q��j[�"�%�m�������U�ɍ�x>�8��,�k��O��6���s���H�`7�ٖ�4�7���ٕ3occ���w���$��<��P?��#nx'�0wmMV����$+��������k�7L�O����4�c$��{�8��`~́���P	�zT����b�T�j�b��rc���آϠ�ta6b���sn5���1\�k30[�I�(D�L�ۦ�Ca�}A
M�/�}�g�C��C�jMF�ʜ &�K�ڱ�Q��մ�����>�t����-<a�ٿCnH���)�_�طh�M�ϛ���`��Y�H��`s�ˠ!o�������n
5�n��F��|"���;�7�n0a��>u�i>
�2����0���V+���"k�^�����&@#m8���⺤�C>}ߺ�H	������5e��ֵ9�)���;*r�8I�L���W#����?*Ig�M�����K� HB�Ӵ� `�^�)��W��+�M�_:���{K�L�o���	�S�}�%�O���L=�\!m�B����^@Oԫ5�h��)�V�o��4%|÷v�<R8��/�\��H?H�$~�.�˿��ǵQ�?��VѨ[A|9�׭��f��+>��*q��4�ע�F�;��`���EM���4���K[�p�,�	���b�CM?2�����l!�K�aX�p�٣�`-A��\]��f"��f���3hEi�o�$�e ,��?��;J�Q}|�qa.��N�����M�;*�c�YLc
��7�"l�q���U�&�?2]0f�'��c0���lg"�� ����8����\�l���3 r%�Y��mQ]YkSں�sG�Gg���O�S~q|��ӛ�"����Oa��҅��c-��KZ�un1�A�A&PFθ��Z�_���ٌWo��=L�f��u��{�8��J)+���J�࡛����8�E�RK���&T5�+@>hbםT�Xr@��d�=]pt��&Y�
�7\r�>�F|�l-�'wC����y�*���S,%z�79���!�A���}z�ň�����~.�P��6�*'���+�"��<ջ��PM�=qF_V�EICy��43��\���ɟ���G��"K,�u��}������B�ފE ��zW�	}���=Qr��1�7������T1&2�U�ݎ���r=c�Y�*�Z��]cZ�[ϒ.���b��-K�#5mw��Φ�g�Oŏ�(b	3�^p�F]+^� <6c;�ϊ��C��I�P�'|����6��lR���&�g
��p>�1��>�������a��4���YM�v9�\��:�x��5� �U�J��!�����)���Go�k�)�'��2�}�B���j��ըB<p��¹��n�4jyMk7�W�nI� a2�8Ȥ��D�ӵ�s�,�}������Jۑ�<��A(\_e�����?=y��Š�^� }�P+�����N�R��f|!V5���\�w.Z:|�`\v�Q��i�@�C��6��?rxH�(�����|-�9��Cv����SQWT��{�{˓��VD;���E�~�&U��	��BTG<6��Aϫ�tN��+-�L���ԙWq�9	�_���!]��f?�H�����v�PC
���>�W0x��BL��,N�8����������1�}?|��'����,q�����:�zJ�<�a����w��x�J���(�,k���:�S��<�-�Z���9�ƴں�f�
�t7�˭�0s�.�x8�a�7ʵ�}G������a}�H����i K`J��=]��"�:�q��E3��q�`.�ޠ�W��'�OҤ�ه�$�0$U��K�mt�,�5��"U�4�ϱ���p��PeGp�*9���S�3	���U��I��h�-�we�]?R��E~����hMD�>y�
ó��y��'ka{���,�{n���(���Ww�����4�"�k�*Hݚ�.C�Eo��[\��w���J�1y�B)�C'�I3j��[WW�`�k��!� 2L����5P�K�h�U1s��Ð��8�7|	&������-�;(d�*3���N�7���a�e-�=��*�zpW��#�?T�Gj��9�z�ȧ:6t�E�weW']�c�~V��2י�Q�i�T�v��k�J�ɳ�np��8̯Z�C�y�?��Y"�q�4ҭ�A�v�)m75��^�	-l�Th�i�ڶ�(:�łB,3�F5GW������*.˃�&n��I�I��E�J�\�>q�|5���(L�g�	D��M����؊cdb�(��W,o���}��g���S}b[���\'�� n)�}}U�S��{w-@�ol� ��BW
0HHO]}�^�v3�kҙ�����u���y6�6#��YM��,V�7G���Y��%{��E��,(����}9�j4"vNh��A�{�S���8P"�����`��d�t��\����CD�ѡX��μ�@�x�m�_wn���Y�rW*�����Z���|?�`Pq�̬̈�a%kA��y�ө��;y�N���2��k�[�iٞ�#�T�B��7Ik�&We(�:g3M��ΙfT�ӟ�+�m^��X+����J?0G�gM��0�0^h�)�i���h֦u�-�*����U�(x����i(��΃��ż_��dL�H��ǕW3�u?���Ŋ3` f����R8��W*�=��4��XT�>�*���6`ϖ.ƹ������ �#��;�Ȼ�T"o����@"��&���I�G�X�1�D�N�+dg�)�{�YuDm�.���3��m�T"�\����7�`Z���R����hٟ��*�o�ѳ���s���9��r��z�XC��x���}����2�Ѽ���3w��>�<����Į�m�|6��\&a�p�U�K��gz��tt���<p��~��a�T�7ze�VGk�P���w�G:��NDǷtP�6ig��\�-����S���nδ/��0���
/��"�'���U�������t�ĽN�q�^�n֑���s����v�I��,Eg��z훺�7���Vg,*�ܽW;dä���6�
K����꫊L�^%������*ct�y)E�}�Ԗ}�����������{eEI�Z'!�[��1�=+S�%�v(�X�b���(�4�q������A�j>�])#�k륇�&�mJj����\:0%P2_BC�����?�Z��7or2�%	s�c���l��j���y�������8��/0��<�5�����}���������rddYh
hoϽ��Y[�Q�!M�>�l�c��E��I3*HhM�c6� �K���&���V�L^��}�|�}�Z�	�f�G]O�=x��GGܐV�a�ky��$k+�o��`�-�߁T%"
?yI��|�~��:���u�k`�|=�P��P��TQ�2љ���v]m���h[��v[��A0����8 3Z<��8���-������洇�;���f�fa&�4J��LHO
��<�Rо���U�f/�U�4b�#���'�r�_4]����6��i��uGo�'���h�^�.A�}��`�0��d���e �kAyP��;����	�8!�Ѣ�	 �s���R�n�P�����c�.��L�Q�� H��f*��l�X�Bh\��$��×�i�c�x��w���[Ζ��P��	���0}��L2 ,�uF�G�w3��)@T�������%�����"f��u��i���Hĥv�q{vXt�_m���t�:FHf�U;BX�R��K�~���?A��$�`������=�����������k_�����hLT�$x��t��/��{��ԃ+�X�e�����U���cs'�*0�C
EA�z��q��PW ��f��ئQ$�棑�J����$�$!&N)�4>v��bP��ۺ�s���4�����=�~70�Uղ�'�G��a�D�#������s|���(���^�����o|�]�
9��!�٢�"���T��Y� ���؆�L��T0>��ܿgrQJ���(�#TP����W6�@��c�|ť��p��\V�;ɪ8$���V��/�����7��Qֻ�kR({���:��f�U�F)E����P���ArX�[��.$�j�y�^����\�`�����FG/6wq�0��H7!A�@�'؝8�6 �(�nѢ��~˒��ۮ�TE��!����������E�V�u֡��� ���Q���BT>q)�Ç�K��j
B�s�3W��A�͕
tV��s����j�l˴����9*Q"�,M
��O�`�XUBߥ�M�8��Z�yH�l"�#���~3P�����ۣlsa�R����qmZ�},${F�� L��Ո�7j�����r�`BӮ;�m�d���؋�G�(�B��]>�Є���asQ�.��)��VX�`�ּ�y�j�h,�p͔Y���q6�3VW0��4
����h����� {�`.T���}��t��\����԰��� �@�o�y9�����������3}�ỉBㇽ�Q�(L�����(	�2Ysow���M�~)�����й�Q���y�
$ePe&=y�e��y�+I"sȒ�X���5<`�b�JV�xVH�fg;$n,�K���'M, �?�O�U��d�m5:�;>�?�tqA��.��o��ٱta� ��$pWF\]d�	�©=>[�aɣ�7F��_J���PŨs�Br�N��:�nA0r��q�&.r��Qi�Q��kғ+W%��\�HK`E4�.�a�^b�l���1��\82uV��q��*7�%��~�-���CWќt橷k��I�����&|� �*�j��9�k���D�O�Q����JO4�ϖ�/MQJ�7�j�3c�R�L�'��^����v�U���q޶�������T���^��h�h>YrN�
�#���}/cHt�x�
i|Ӌ��a&/����me�ty��Or�T���}֔ i�������U���vΒ�5y�a0������H߬<!(>�Hӗ����ne>��&�M&KZ�hZ��c!��a���m�7l����4�	G�Te���03?�C�-�����ӚV���}99}U��1!LVA��j���*O?X�T&KAԡ���Uof�T#�Cۮ?�o��$�Z�^
Ǚ�w'w[| �l"h��؟��쌂�5s��k�E~���c�<�c�����&bj�ߍx���IV�(��pm�s6~&�q�z��Eڵ^9o֡j��\�ҍ�)�R��Dr^�,F�&�Ր�xR�R��	�+�PX�T/0���}m�����
)�Y��]MY9�kd�}��)�PMچ,�pI���ns�0H���m1i�O9��d������X ֝�R5��I4�E�r�{��;�dҶ��^����P ��o�}Y�e�%��g�M-��.kR�],�6��T[7a� �!R�޽=���f5���k$}\� ?����h`�3�r�\uh��ҧ���h	�w��y�݁���-���7ݑ8neg;����gcC�y~X�X�̖T�B�<���HM��piK.N�*݉���ם������b�-`c;����Ζ��JDP���\��Ywx�kO�]��y.@�����:�>���� S7iijw��+��}�߶6�G�Z*S�6�$��l�$�`���r���������� Xa���'��>�.G�m��\Ud.��~�H��*Vc�0�a�g��+`���c��_��m�Eo3C����7/;'.��Y���e������u<Y&OU��L9 =�}?�)wA��r�R8|������A\`�Ȧ;�ԁ��{ܙM`Q��X�i� v�|`[�O*�maY��Z��1�ڠ�ž�03A�)ŖDoh��Q�eM�i���X-�]����]K�W>-�I=�2:���);�H�/_�lv�_��F{pnZ�.z�(=nq��I���B��e��hR�W��_ ca-t?��)��p8�Tfx��R�7B�����H�8
��՚Âs.VS�[�ӿL(�{�59촘�d��a��#zЦP-��Oњ��\�t�
޷��b���_����f\?��	S4_f�xX��N��E�ҩ>j͵ˎ��*X���-�pt��L�S{dwƾ`�N���D*�;���WP@]�B��a&���Q~�d�v��M����ޅ�R��(ː��2����c��X�s) j�@�K��)Bab"#y�K��I� V�,���z4��ԩq�Q-��86R~�S�]Ԍ�ݧ��C�!���%'(}�t-1���)��l�؋��o�P�	#�Q�~��ڼ0�e\�.K�	qך<��6@�d^z�	7e1H��bJv�fF�$�?׳��qOK$�	w�h �Se"��|O�D%��������Pe^ʥH�C�Y�����z�U�{��;0O�d�t�i��06�T9)uxLkߏ���%cU|�|�H�q0J^C�Z>&��D��42?d��PR��C;��e�S�j��T�)I�!����R�^B4-�yC<b&���^t�7����e�L�R���Bs����a�#�`��9�2#tG��-��a��-�'�����R��GU'I�w�x�Ռ�n��7��$������rɞ�-�PFJ����m9�nh�fNNSͲ�>;,q*�`�O:F$�����.|A�z"�Y5�	)
���.a۾�D�Xx 0-�l�ʌ�}ޯ�[d�{�N�鯇@;�� �P� ��}���Z�k�p�)T�m�\W������-!�. �s?b�R���t��ŧ�Y�xeB�wڒ?`?ͭ}�L�#���8g�}D-�Z-
�Ӿ�'��R����iڟ[���t�����TSIUϺ3{�s�:�,�ͼ���c�K�W��b��o�����;�(�>�@�&5�	 >�X�9)ell�U����9�^=8?��Y�A4ǭ9���AH��_��G<�4��)��K=*.�c_7POx�h��g
~�� ��:�h��8�aa3AGJ0�G��Ev� %~��H���S�
d���,��r��ޣ�),��,1Ǚ��+DY�;���I��+��^�#�x�m���,��	5Ӽ����Q�e�vb��M����L�GG���@�ºPߎE��|^9�\-�C��P�$\y��6���@UI.7$�Ա���)Hc�UZ��T,J�t�����%�]�\-w)&%���u{��d����� BnDoEM"2��Y��ʑs�� ��x�I{ι/��>�����B2%x�
{BO��5=�Yۻ��<� �KO�-e��:1rb����i�Ŧ�"�O���w��k�z����.f�M����K}/2��#�~�/ �+���b;c���x�V������
�p$$K���܍;{�8|�I)9Ȧ8�>J/e��!^�m�)C>7|�ˣ*��XI���lf \\��Ia�J�c~��I�-'BqBPsp��Z�dpN��9q�����NAp��>��V>�G09�t:�T��T��[��Z���ɫ��~�f�T��t��\�4���1M8JA	��{�&}AQq�,���\՘�� 6�����/�kC�c��㽻M��y����[Ӡ^��˳�|=M��ⱋ8gZ3�p��������P+3���J@-�,���7Ks-�t����U��c�戧ض�cF��B��E��iԯ�j�<�gS��~!�{��%4�zں&��D�{�z\z;�n��)r��K5�m�G�U%��TH�~��$~�i�f�̙{8�!��]�,#�n�pR�P��)x�8`G���gz��e Q���e;Ϧp�;�"r��e��^%J�o=
�UhȖ4�xfi�n�-��E���ԬOy6�,�����py6�h�1��H=m���\�E61���T��/��2M|Vʉ�ε�y�\�9yfJAG	K6W���W�j�s*-�n%�+���&k %��}2��0�����"�ܮ�-���q��6�A-��$���"��+P�^a�09Ɛ��O�-d�v)3���
]�R��"�`�����F�X�ߌ����Pp F��U}^R� )����k��)��4K�ɼa���TNZP�	��<'�l�"����e��DX_(���[0�?8��gp�MH���b9QY�Fe�Y��w�Z��~[Țݛ��r�W?cAm\��GMR>~�4���w?`�ީ��5�鉧6sqU<�J3!����T��\*|N��h<o��)�L�Z�����r�����X���R�wJ�; =]�.�
9	�2:���d5�ye9΂����C�59&a�$��@ax­����<K����v�����Λ!R�`>�����G�h�?X "��c�	HJ������x#��M#O��쑵����̓_*��Dka-�_kL�-�����aќ��Ȇ�����]zDc�D�Nxh9+�a�y;��Z2�	�� ��<O;��u�Z�,�wn�pZ�Eq��r��Zs#�z3�R�l_��?�N�i�Ew�arP� ެ�;��F�O"�gU��h|엾+��껟'�#N��7	6�yB
���y�'�M���� 寄|�0i^�h���aVG��c�=���X8;F�����wD�T�����=E1�u�*}�R�<O�p!��È�~��V�@,�����8vO���a���Bp6�Z�=�|�7?�c?u��Tl�I�#����θ�z�l���xߤnH�yß+
��QϣK����y���llHgD*u{pz�]\{.�&	�2P2{�+��BW������ǫ���EP@g�X�n�u�W
8�����,��>�J�ά;�%п���M*�h�5� {�	��/��Ѥ��f�
0��oS�k�^����T��[��
�A9�r�~�b�֒�(��i�O7{=��hxXS-���Qɨ��0,x
`a؜���f����X���Ê�lI0-����|�b��s�bj]�(�E%%��A��tz���v��|(ch���b���$�^��*�`�.`yA�Ԑ놕&�\����V��Tt�Qc�`��.�W2E0v��W�H0TH���� ��D��G�FEdy��y�c���K�@Sl���)l8����;Ȣ�ܴ4�\�2�q���Y��7G��lʩ��&� I�ZݐE�,�e������R�O�b�[�Y\�%c�U�۠1���"�<�W���g�^����t�ϰ�;y\��C��*�K���j�v�RT�,�]x����f��V�]Z�����1�0��qcF~���
�@������A�/?�g�����J3�D�*Є�$�m!������A�=���X!"�Sy#�{�s\l���F�j�${a��4�׈��t���XY8e�	���0�JZ�àE��t�$~ut�Z挄���	�܋]u�6/迮U�����¤�,���WA�ϹI���vD�	�%��P�͡�`.�n��0���4O���;K�M'**Ƕ�׺n��mK	�u'�k��/���X�Š�_���l�����gЯl|�=M`�