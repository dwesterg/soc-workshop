��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U��:hZ'� ���k��WO6�����x@
�K'���,��������4�V�����ws%4pD4�DC��[:(�ف�0m%؝��z�}*�˦��|�[���h��%[=�M:`�!]	2-�v���o��r�Z��B��l\[�������[�1�/�Jo��������u�wk�H\��,�\C؝m&�3�P��Jd��|MA�������8��z3���=�Hd��&�6J�9�úH�T��j�������@Ș��.@E�{Eҝz�� ט�5Z5�d��i���8b=J��y���YW.PSN�MSΉ��I�փ9-��Čv�4,���@�t�vŰ[����Ϩ���r<���᥶TQ��u�0��n$B�����Fɢ��G���E4]A�hx�hC����Lw7� hŰ�%my�7�Ik5��S���h2Q~~�y���Y��T��2��+;r���R]�G�W��1-ne~�X���R��$��ڞ����C�fGQ�e՞d�m�~�kW�e�� �\���~��PԳ̉��;�U�0k�*O�����Ţ^U�e�uRi�!yDΠ�BK�r�`wX���"je?���bl@'$x��+��-�'5�#LA5j���T0���U�A_])��@�&��zH�I���qD�ǔ�	V�(�׌�gs �����{�R��Ϊ\r$��\��Z0��6;g���-��E|�A�yv#"ָ=[��3r��c�� �z]3�;���d��ų�Z��>�� �\�&]}z����ΰ͙-�>���qv���Ӏ���~���v�?@�6.���Ĵƽ��J�A�ʊ�p:�P�"��%ԩx'��ҷ��"a-�����93�z���,�נ^m��t��T��'��g�FY&����-Q�%�����B�fMM�r��A�J:Q32����6uĒKt{~��������Yu������Y�\��^+��늼��P�O��e}#�1�XA�q�"K�f���c���յ�i߫^=b�����D-�~N�����4O�H��ؼ�W�Y�Yy����R���X�N�QF�_Y����	-�,'t�u>�v�3�8[���t�8�>����+Q~���Y[�p����-<i�	�ༀ��gR"ז�S#}��U�1�i�j���$��%f�!���7ߢ������35ug�\-7�k3�Q^��g(�m��5N���y����
z��=V�@��OK��e{��\hQQJ�,5�Վ�$c;U���E�h����WϤfgR�D?�Cp!�vm�_l���]�"�zMn̿e�[�eI�%I1i�1��}{!�	!~j�P���ѱټU�&^�B��T�:��T}s.��w�����k�@G�I��9�[Y�=/���D��7u����@P.����۱��	u\q��*,]�fT��mb�rٵ�έ�g�7��Y��,��P��<b���=�W?}b&g7"��tg������� ��,τk�	<O��d̢��=8L5ބ�>��
�f����>��v�ۡO�5/\*����A�����07Qy|���v�=��E��gO��ۉ(ڦ�L/ރ4Ob��&�Y0뭈��0��!���:C"�X��Phw>���������G��_.���]&��������j�I�����Uat�uk���)�w��$z��35.ݤ�bW1��D&���Ҷ)ٕ���sWz�b[Ћ�^��I�؁Mz�x��'��F�:���}����X%��{���V�2�A;���8�e��%��^0D���^������	�<a)BP@��E=go��v��b�%1x��h��w�^V<�\JIq�I?Tq|�;u��^	#���.�2Q,m��!:5�o�[f�f��bf��(�t�J`$|.��2̀�U���ض`�+�x��{�*��_��x�CεT/uQr�M"7�b
T��.
ю�bYJ�	���Tj��;� ���h��Ғ��/�p��~��n��ڄ���h) t�����8�ʇ�\?�r��'�H�%�����ssZ_�.��`<:��������Q��v��A퍬��,������-}��*m�j���P�TRs�"Yc�����rX�_f��v~�T�ZTj�Pb4��#Ht���&/� �S������]�l��i��]/��V�N�R�-%�s>Hx�������^qxz�55��"2m@��;���o
�&�Y(Ӯ��Y1xTZ�%Pe���<������K�_�}3d����m��?���Goۮ!w�i$�%1>�Z�P� D���w�/`�ܓ��K����ϋ=��U����㋬�v��
Ȏ��c��x��ޫFl��:�#ˁk|�tf�2��#^	瓕��L@��ܱ��#�\V� ��8*s%�&(@���yyN ����}W3ç]/Kg���d���K� �,,�`od�,�{	Z��]
D��"d8|���u}H��EQn�I�K�&A�Q7%���U!q�/��@2�B��^��Vtf���|L�KJ��R��,�K���Jp��Y	[��D��T=um�R�i9���@]���?�!�
�o�]�Nэ��	u�:��&P"q������t}�;���D��|Ɓs�d.hy�A΃cV&��N�''�A�:==���!Q���R�#���M�rRסԕ������o��<!��DOS���m��
���(i
֟�V���ć����3{��U!/���SR��['P�ਅe��}�;�w<f�ǟ�W1��5�0����3
��	�����1��C�ِ���:�iV.p������ߣ^���%��g�P^n!A[f���P���̜���եx�����Z��>I0��r6���N�ы_��w%��^�m6-Y�K��D�W�����W�;���r����s��*��SGn�H�$�Ȋ0Ǽ{�[��<�Wv.4�uD,��0���V.sD:���q5�w�����.i{:!	4�ʙO�]G(��*-�i+w�b�_��]�o�]��Ki���a�64���Z�;Z�r�v�g�aX�o6����QGr���2ۧg�a�6����0bΘ�.���>�	��π�Qj�C�j
��>I����#����!�]���@�BiY��=
Jۜ��j��A��k�5-E�{;/#�d8��z�hYi;���gr�2�1����/�W�7Ql��P�{nn�F���G��O%yP=X ���W��i8G�A_�F�|o��0���!����v����E%���Q�R�<��5qCw	�5�4�ٍ�K�Z)� ���.��q��<j�(�B%w�����ɪf��Es<+��K�Vݼ`m�,��F�I٫��6�v�w�#�[a�;B�O����4��J��8��r��ϟ��~�LS���f��A{����s����r�F�bɭ�9RV�s�sIt����UA$Qw��Z�P���#8�}���m��ϼ�D�h���4�]��P�yo����Ѷսw��,1VJ�6BC*����,zN���P���HJ�������<�}�K&���F�����$�X��~�-���<8[�ևb1�5;��.<�{\}��پ�Վ�o��Θ#2���Ȳ-��rV� Cwń��m{N~b��+��vީ�JjZB<f����2�S����)�N�W�\�c��&�$�ԝ$�[�A��"�"u�C.=.#���+jze^�,BXG&���
)-=׹6ݦ�Py��#S]g�K4d�O|���̂h�����M6w3���r����h¡�Wg*j��ީ"��B����|�T��?��¿$ӱ{���K�.�
�l}/�2�92�p����,��,ܡ��F^
`����湮�l��WSr%^�ྦྷᚓ(Gv�,�����TR �x�vOY��ߣ�Ȯ�e�+�)�#�s��� �ـھbb���U��#Vt�����X�tpjeÈ�[�{�zc5�;E4ZR��;�[�aJx�������3gp}�D�2#��V'�`h���Jlƚf�\�/�$@�\)�v#ƻ������<��f�����ĳX�˃���6�������&y*(��M����KbZ`����H�.e;j����צ�� �v89*.RuE�A���	^vA�O�5�%�s�s�����M�J6�R�m�}�F�߅,ipg<�=WГ�TwG�����Ļ���q�:v+Ѓ*��1� �"J�<��w�IS~������_i�:���b2�L�'��a:�@�C�b�J�E�,�6�6�3pO�!�n,���G"�~�HҰ�u��w�ύ���'1����q�'e4K-{�Ejdjx���xU�qu�%;Ҕ�����HU����/��#��x�e߶ƔT���x9@3B�Xeo*�y��٫o�ˌ�53}��P!~����ns{���`��L�S!D��������B�=s﷎N�0�xʩ,Ѝ�x'��R��T��w��"���7<@���K��5;_X
V�:����g�X�A���͑��Q���(�%#2�7��2��B��u�9�όw�!�J����
� �o�W;4(�i���%�/	򪗚9j����;���ܽ�����¿��?�8�%��5�/?U0��aAmYb�<�������aۻ�}��m�uU�FS��B��}ʛ���C�i�:�<�(����7f�;�7�<��5^�\D/t��0�0��Wi��}���.�G�sR�&,:#�/������	w�~KE��z�ۉ&-x��� \��$� �c��I����
)�\�jG*�)WM��EJ�	tF�OF�uw��ܤTH�3����{����W$��%��P{�k(�b���iL'�k��~�6T!�KB�"%���R��/?��>�$a��q2��P�(�S^�2b��7��j��KRb�eK�i�o*������<���
�9������Y�Qq������ZB@@�8����L���Э��8��m�ߥ��Ϊ�z�3���oJ�\Y�70����l=�y_�D^vvK��L�@�a���p4�H��ShE5
E�ȉ��~i-�����_�K�+H�M7�9�^���0Q41{�C޴u �O"G
���{(����$��(��qE��8@ʓ0����vyd���6S��W�����7�+�xV�XgRϚ_#����d�aR��=)�JY��:�VYfo����D*���&�����L���Zy�����Ԍ�s���9����W�$X�X�[|��#�76���?I��s�!�S
jg�m����7u`�G�H���n����A{̣��zF�~���
�/ϩ<����]%	�G�OC���j��F�7���]h4Bk��g�r)�� �6�D���^+��2�$0G����j����\\
@$�+_ۖt����(�(Ϥv�K^CJ�SFUȵM(�vBT�O{e�X��ʰ'��*�����E��:��������mʹ��*���h��Sx��Q����C3p����5���=����{R	���:�f%�����N��hU�~��N�-�ذ�w�G�Ȼ�8�֞MUQȺ��-��Ԏ�J%F�<h֓<�����m�=������S(��^�����>�݉����+L��s@�A4Ν�_+�}*���.��>�Hz�VqZC���C�n��7���j �����6,�J�'
��#Y�i7�O@ ǻ�ۛ_�Ƌ\��Ԑ�B!���M¬/N��
�
����sL�џ�СK��2��� 2�*DWE!r� �F�'#ߟ(,$����1oMyM����5���g�Z�����Ś�:#�+aO�eV�ÐG$ѡP�dS_c������Sh�N6 8������Ӡ;��T�)W.qAr�cQ�Oj']���!�vY���g��柳x��i��ј�Er�Z#l��/�w���a<p[�]-5��I�滁��0�c&��!�����T�����Z���S8vN׌g�J�9|����B\/�Y�w��k�_�L����H2��B��0���,�HLe�� ��)V��y�y} ?Ⲯo����&����#��Sd�S������WA��ml3�W�\P���d�>��}.��}vCm�[�m�G�W�f����[���n���Q��CY�HL��U�~�o`�E���-�� #����2"2����J�qh�������Oؔ4�b Y�������z����p9�.ET��Zd����!��ז���64�*A�j�t�[�Ü�������2�]�Y�B2�q��'/�n������O�Wcy8��\9��U�i~�B$;Or4�")��u?��9�n�A^� t^O�|-��c�j8��:[T����~�%��d��'	�(R�q��&
2���Dpƈ�_y��ˢ�%Q�G������3�D�VA�g��1���ez�VJ�p��[�$�	f���E�ue���f�~�`��a��zQ��R�š۵}"m�_�8��l��I�5��K��ؽtWW���JҬ���SI�����Y�)	H���Fq�?�Og�DU�䒯��{'ĲO_+��BQ�PW*
N�kW��Ǖm��v�&'��ޟZIjfɝP@�74�P��Qׄ��	�[�H� VK���ꅌ�
�&mGаª�<܊���.�'�V�w7�Q �7bmD�I��1�)��U!Bs��w�j,\L��9�#�?�"ʙұ�li}���!aO�ǝ,]�%@Q	ˠ4���iP/�ڝ����;i�>k!)�N�=B�YP����=o���P>��{�����E�ȿ7��:�j�\�Ȭ�j�ޜO1��X�R�Q��T��g�~"ͮ�Ѿ(�z��4�����9��N:��lR����(��YoO�������M`�aQ�C��F�)�K��a%��~���i)*��A�n�ߵP�Yk���.�[t�򹖏�|�wJu���p���2P
6O�Rd5������T�x=w7�L�j�r�an_�>���ՏC*�%��>I����c�y��Ϛ�/ �V���&>�����{\\�ܺ=����F)/ۘ*v��MU�����I1d����֙��� V 	�'��B�Y�sԝ����Ƣq���Z���*��M:8Yr�l{E�k��BY/������@x�NB���(��1#,e�j���pm���j�N�T4���E��"�6v �s�@� !�j�BI�'��ɪ:4TĮ�Ax���4c ��[����^�՚57&}��x�+W��o��٧�:ț�X�'@YZ��#��W_[�m����`�����u��q2�>n����� Ca{"VJ�]�̋�3����p�oJ��5"�mV"�1�l\ui�Y��P���F����ɿ�@v�=Sp��f�f��n��j=�c��I5�;5�K��((#7�	�?���
ל��
�ų�>-���L�0
;��b��V�=�K�գ�R��v�i�9x;���3߫��+��=v�Ia�\��kK���X�Ǟ�NU:����`�=�+q/�� @tˤ��;ZxR�(QsK֡Fh�Of����Pk�o�5�h�O��Pt��h��<�g,�q<^��X���d9���
��e�i\��G��mh��� ��9H� �o��jio3x���<���&4�h0�W��,k.�ְI$)�j�����Fk6�I�8�Qi�8~l^_KsF���^������x��"��\;�[�^]��Z���F����GJ�`gʓ�-�R0aƣ���-^ QQ��Qx��<J �X�`G�
!��??���͋"$6�0}���Ȼ!B�͛��`�y�ҙrXn��q�VrE�0�����B����xo9����bYzo+��eN�����F�����l �E%;@7��Z�����[��ݫ�/�Z����Ț��^�Z)R�L�%U�W�5�~-1C���2�����e�4Z�!!E��xR�t#&x���{ X����
ws�P�FA�9M�&��ٲ��2��d��Z���I�ײz�29���v�f��Y��[k��a�6��C�����p����z��7^[N�O{ô@�n�=���Ģ�a���7\_u!�n� %?��"<a�2�-����j|,���s�+n�i����HF���=:��fIf�\|�}6w��zz̩'u.��+5W~a̙����W�7��1v�W���'��`�HI���Eђ�����$��X�W����RH����0���,�O�(9ׁ0rf_�I��C�,��W�m>����J�F9�~u�Ѱ޸F�u\l"j���j��[�[|��H*��x-�\S(�����=V +t_��A�M5��%9�/{wf�V�l ���[΋{���%���o܉������@�#�J��n�=�Fދ����`��]�5���7]Y0Д!f���QMH�K�p%���QZ�D�/C��
�B=��x�5�?��E��
��6��xO���G��9�,�c�׋h�ǘ�h�m����m�[Ԃ�r�iY�k����9�e���@y/T� >=(�ބC��Z�؏^���Q�k��y*kf��;Zڶ�Ӷ��I�k�ILa��@���gR��C��$�cs�����=�n��I@%��g	���z���|���EMh^�����σ���ڑV�^���N��V���G�XrV�o��9�^�mN�I� Q�2��=�j��D;>���y�9�Xgh�f�ԇCwPW��-w�&��2E�X��{��h:��5��l�3�����o3�T[�ߣ2"	~��J��L�Ŋ��+������u����s��0�{��>���F������Ĉ�C_��WQe��Ms[�ܜ,�?�� ^j��'�r�ڳD7�X͈�vpYEIܡ$k����U����_�i���W`Z��~�p�P�!��o�Z���]���J ~�i���������ũdg�ν�#5ˬ#�����s�"��M�4�%�$��+z��������q��ѭ�s��.�=(��B��L� |i�p�ͯ09MjwF�60�g�7y��p�k3iE��&s�B=��O$��Ͷ���#��37?�$A?�)'ى݈zŴ�,�.Vz>��ө��=엕�RB��{���/|#$��.pl�vo�2�OC]�`�e�Vy5�ծ^xҋ} �$ ����&g!�+�a��������d��`�*.�y�,Yz����� ���B��@�rI�ˁL���D���E�J���6�3�������й�^���h=p�ʕM�=.�+�k�Š�ZQ�!3�N����Y��k��/�ƱM���6z��*�ޙ�z�cwJ�)b�ڧ%���ʿw���ś��i$`����NdCD�;+O��;��~�
3���z&����F�Aͷ�"K��~��	s/#<���d�W�q�":��y)N�c�הkBǛKq��v�`����{��#Su�a���ɧL��� G�[P&ѷ�έ���n?�����BUr$b0�]/�"Ǔ�(V&����
f�^m���#|c�	Ԛ�� �DZ|�w�0�廞�>�캋����X�.�g ?zͻ�
)�*�4I���C�����+،�y�Yu��q"��@66Ж���Su��|��!��1�`WaȀ�h,D=q����N	���D�Ѥ��!���� �\<�%��
��S�K����|nM���j�`��Tr�"�y��1|���cG��VnG��6��P��K�����D�͢k�<�_ƪ�!pB�a:LVt���!}�y؋�-Y&�M^�)	V'@3�����\�l�����U�5']����ߩ*����g.�
��I��[7GԺV��O�Txd���X��������Myo�NiJ<NJ��	�w&���|l�w1Z/�K�_�]����=����c>�yz���@}�6vQ� �J!�Qt�'��L�l�7�n�`��d��C��9���j^I2�Kp��bsv���R���F6��]��.����]�c�]��چ�L�Ss�-Pb��%,+��י��>{Z2��P��ϋ�
f�_6]���fc;e���
-*�U|�y)�
���d;��cL���Eˑ	W��K��uٳ������Cq�/�sSW=�oU���:�CO�sʛx�'\�M������
x�ʑ���D��W޺!�e�aȌ�-����)�e�o6��b�Pe�	߯R���1�K�8K�I��t��<�s����H�����F>����ج�wI�Z�u���qJ>@p\�Q�`�R�K���L��h{+��ght{8e�A�ޗTxF8�d�ڀ5m�:�U��G�G��H����*�be��c���PY�ҭح#[��x�f�v�b���F~3��Ȭ-�c����cUU�)!�h���M�N��;8���;���N vL��c!_Wb!��TS	+�GxǙ���뭺,Q��u����L5p�*�/oh����hB��1��}���4�0T�{��8!Ǝ�#��� X�̊X�%�1f#;&���hp����Azo����)�]�{���\c�In��­A�eyu#@Aa�%��ަ���m�K����������Xq3�O�
rk:���*G#>b�>�f؀k:�DTe��B�P��!?�}�	M�^�կ#;e]�'g#m�_H��F��5T���0�v�z`�柋o�s�TPiA��ɯ׵�:hٷ(�(�ld�<6��R�L����Y�"i>c1hC�,�\�{�#@�$HO+:Wt�$���i&��|J�8�*�^��[��U�`Z <���݅�_���K���wTFؘ,��8�7s ���N����3	�!io�[؆�`���Y��)H�-��+΢=ǈ��-Q�L9�S�[���=��Aa�E��c}��~d�J`j���l)r��/1��.YWqU-�/��2�;u�jC�YK�G��K���14��!�}URو|*��Ci��lf4�"xcsnz-��ITG�����wpPKm��ζ0׵?39b�,(�= ���[Je����F�ŗ���fV%A$�)�t�"��pf�U��OV�?5"�����ׅ�	K5�h��Y���Æ�h)������\<:�2��2W�ӷʰg����J�RL
���n�^٬��`�^?���+Ĺ��`Kn��{���Z��WBRy}�b-��Z�L�l��	�2�`�c���13BƮ#ᶥ-����M=��jx#vي�׹2(c�+�����l�$:@w[ۡ:E��hkq?�
�ڬ�*}(O�k�H��ei)C���0��T}v�YE2�26�畱z�j�^v�J��ٮ�)�����_�QqV}s�>�	W�k�ڪ��D5U�	�O�"���T��*59P�뎒� 9�b%�Ճ�8��kKO�	]s��OF%������D(9������'�-�"��(�s*Do�']W][n]^���y��1��}rG�����Ku�tD�ު$�b+�E%���"�I�
P�uUBq�zSk:�_�4�W��0ΨYXyC�nr1�q!�ph�S>��v��_�:�Z4BBa����^q�R{)~ٜ���'J{�5L�W��#�E^*$�-�����uhG��73Y`�U��_�$	.�� ����]ْ�N[x�ov���w���G�ݞߜ�rʃ'�Iȝ�U��߈�Z��cnr��	i���N���PL����0��e>C���|BJ��]�~�W�d�U���Z����i�ƳV!hZg�U���0�yq�_>g�b���q�"�r��s2�bG@&��J�S��?��	��YS6��M.M; ����O��������X.pG"�~#R�b��P�g,-�
5V��5IME���f;�͵	�/�H�F`7�+Fs�)�(��b����'�]��T�+"�X��T���ueI�m�b�$��s����L��e������~���$����p���#Q��F7�]U��PӘ��d#��b���哓�Pa��D��y�̏�u�-y��0�'9�˕W��
&��'T𬰛i�у��D-��P�ğ5\�1x~���!k<f�����aA�,O׃B�����X0k6�qL!.7�w(�����nP
�l��D�-���Ʃ��[{�3�+IS�$�KA��`g+����o�5��(����S�X�1�H�)Qj�bI�e��:8эW�ul��Z8b�_��A�Bm#L��MO.}wlq�	�'�v����й5_R����w��?��j�]?H��Qrʖ�(�����V0�������1�A��*���^�Mn���I`��#g�k�94P������+A�m��HQ�:���.��Q�*�E����P�1P��2�?�$��>��������W��5��M�������������� ��҂"-�;S�ʋ�Q�ڤ�w����U/��EB4G�Wɓ�Z�c����2��pk���<0�O�d��H���0�2�Q��{ダz�\$�ՕDD�*��]������֮�P�J�A+=?��e"ϣC��De뾛���y��v�UQ�K�5QUͅ�D����F�1�OZ���^�V�U�:ɠЇ���Gr���>[t|�u���������F[�מ��/ �wk��
�B@x��I�EjD�7��.)R�+��);��6R�+5+'��H��GK`��#�JY�2k��-�p�V��]��m�6�t[bX�W���B
�y|�f@�^�8�Z!�^֬�͸w��*�K��dz���'�"w�e��a�i ��8Z�Q��̝g.}����\���a`5�5=�����Z�|=�rԉ��4���
#��T��td�R�2r3��(��lY�!��P)xv<�^���U�c6�[��͸8��)�K%!����z��jw�q�QB^I&�TWpn�Z�T,@�x(O�c������Ʋ�5�����؄��n7�Պ=~J�ٽ�Ԗ�*�ll��:C�N�78�f��X��G����}w{A�+��C��;�A�5�������<��R�'��߀XJ_�)�GP-�ƀܐ`�^�z�y��q�5��G�L7��pTڀ��!R�ho�t~ب���֋`Z�0[��7�ɍ�wMi�!L�x��^�9g��w!�������ו�EdCE���v�n2Ԡ��}��gN�K����z�H��J7��t7�{�4�]�T�Hh-i��q��V}��9i~��HuC$ǹj<{�N#5��cxRE[P�Qڜ^�]q��3n����Q�{�4���+$R
xIlm=*P
�+��,2�,�V�}]7�4��=�>/�̢zH8�P�`q��h,yJ�m}n�m�J���u�z&�ʕ�1��d�+�<r��	�t���"7���# ��!��9O}��/��lP��_�%5]jAq/���f�@�!EkOAL�l�S�g�aQ��V˰a��9Dc��	Z=��?)K�[(z���Gs��0Q��c�,g5E�-�Q7Z�z�rKLѫ!�L%��&\2ʍ�4�-x��?|������x#�*n=��iД���qL�W�����%�\��o��
��f�l���?��Z�k�n3��v"&�`>l�/�g����]]��2(#%<c�\��!E����]?7`�91�
=r�W�h���S..�`Q&_�*�Ȋ�"���|39������l���Nn��������ř;�Eh!���u=�W7�ĭw cm]8���<���+����x��)�{�$��x�'�N���r��w7~���!-��A��6c��O�q#y�Y�$�}�Cqo�	������7�σڶ�|�T�2b��ik�萙�M��o[�پ{���$4���7�1˛�WT�CW`PN5�Q�Q�K'hi�)�b_�f�������d(38�)�b�t1W�%~(b�>L��4U�/��n��ͭ�,��d��e,�ҥJEt�w���*����� �d�v�x���5�a�C�yĞd:z�N\��cX��X�	�<UՉ�=��/��D]da�(�󊿇�_�����f/�eC���;���x�O�g�W�$�AG6�l��+m6yL<ȏ�{��-P��N��3:�� Ɩ,�Cx�V·��G�&��n;�Qd1��Tl���ʁ$�si���.���j�-��_CZ]'��Y����Zp���=ga'�A�u��\��y\���ꛏ���o����ͥ��>�*��On�X�q�A��1J^���7�.f�*ؒ)�$��s�eH�'|f�gQ��X��Q�b4����k� �������=ؐ]V�Z�{D�a