��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�íT��0!�2�� ^F����mWTP�~�rn�N�]a̋�}�Gm�#�%9ч�W��p�hSgD?�W=�՚�VG��14�J�D!�C*����ȩ���	b�T�r�W0ٖ\��xa��ȣq.�J�0Tp]�)}��LW�y�d's����,>"��_QJ��g����'���P(� �Z��e$a�HN�3��>&`�B��4�,���	�	'����|�(3#2mf��a~R.�u��HO�yrʃwM{qo#0�v� TBV''��K֥�Og\��;Fy��lހC��H���,"���2ѮX�c='�K�&iɋ?���)�N�}��F�b��d TEO�p��F��.�((�bN��1s`�$��#�d�^��U�ڒ�i	��pَ&�mcKrc�b?j�h��_��(B+8��-�sx�H<�tn���g���eW����21u�<����w���y��4MY�4�+]':���O�]^�T�]�1��6\��L�

I�6����rտ���v�(�Wušhhc
������9�`�B����iс�. ��©b/d��?A�U���� �yӂʡg]-L�57�6m��U�n��i��rCD��͠m��I�����F5���&��z'��t����!�S��*��*+���@v��o���0��yǌzڥ�e��ӱ✤w$�� wwm�1�f��pd{�w���w�$wU�T��� `��gj
�B��J�
K6�y�۴�����	��#�L�_8	h�'�@�|-�$T~�d(+��4�ʧeD����aA��r/@�q�wC�z)��u�)_-Ha����������M�ݑ]/oo�t���%ǭ{�S�}��p���T(�G�7ޓ��DJ�T��{�V�o�T��i�v�� �L����ʹ̷����(Y8BU�U�5�"�C�R����� �@\�DH,�o-f�ص�>�<�q�a��GI+Ѹy���x6攆P�N�6[��m Nc�(��yԭ=�63Lo�$�����SD&3 �
_K$���_�om�ڮ�R����G �J?��@h��냻�"��G�/�2%�K����0eX0��q���+����k%*�=�V��A�-5/��T(�� X����_vc�\�����/t��z=���wG�n�Z'��YZ�W����L����kI	$���h���KJ��Α�/R0��}�����o�C��칌:��I��K��3�7[�������7��ey��Կ�V�*Q꽖�����b����5Q��(2C6����211������mX7d��mzZ�"�0���X�"|�uج�ֵzI[B��q�����l�D�P�ah[�ӧ�J ���$����5:�`��K&ws^gB�פ�����9g0���a�vF��jbcY��ڀ�$%��XÈ6��{C1� �/���Kgj��W���Tj=�BזFl�׊r��AYM)p�Ac��l��%�r�ŚJ'��.dTO�lh��/R�yk# a��(��sFV^#�h ��� [ze��:d�h��ULg,~�鎏��
�9X�[�?Ȳ?NȺ%��� ��q;�Z	Aymf�w��k�e�L�>';σX��XP��4{C�[��
3u��>�+1�I��mi;�G
�\����|}:Z���"�AuI��?���ɕ��{�E����?D����˺;����`_��@�������T;���@̆�����;��U%~��l?�I{U����Ԋ��(�����U��Z�h2����0�rK�:�Y���G�Y-�Ӫ�^v��V�^�u�xoG�³�e_��D�vF��_F?:,�W�K���0�2g���d&�1Q"/���_).�<Ť�����a��N��]#`��|�1�)����#{�f|��F^~��b�8bl$}���6��}�Ia�D��-���<�ԛ�D�e�2��gS-��F�#r��L�[:��ô��Lߕ`J�"�s�,s��"�e�t{�˲����F�>x	�L5]D�/���T�M_�8J��/6-8��'���9�dX�S
L�|5{��1�W���9��-��
�����r���C��7�f���:B 	3U��Re�k��3������0�0�i�,丟25���G�.�������U@R��Q+hs�
}\IK��������+]t$c/�﷍o��lD�UV6�''[�Z~��� �Ѥ9�]Mb���;l�՜lV7�+��ޓ�HV�N��NQ���M59�<���V�0 ؎�����״x��ij�ϡBy�/��a$��;�#�^�ۜ�'�v��sSr�§)N�	a�h�1�@�W4����7E�i�z8�2�E�W:�e�Q�P����[���\��8.�On�&���9ÌZ���w��lհHƬ|;^�_�n�Y�W[�Pّ^�Z������Ch[�[ 4\nG�R%�i0q�2��ض�$�2�ɧ>lX8���?{�yd���щ�6Lڂ?&^�j���+R 0	"\fP-`Txi��w�9n���
&$$�ѵ)�5�~���Y�1>	���Vya#�53h�Ձ-`��>#:mPwN2)y�ߵ9��Xq���?1{�Vƿ�hEGQ8'�2�z��a��u�=/sT����E���ʺ}�N�j��D��퓓��!�*̘d���O��fh��O�¬�%��5?^vo���j���̬b�1��ԛjx ѯ�Ƅ��n� }�K-0B{u�PA6:K��]sU��P���*�A9G�I��Y���(��=9����/��� ���T�mJ7k;f8E�OկR�,i�Qw�������0�'�{#��w�a���h+ǂ�>`Aؔ��
�-]F2`b�����K���c r��zN 8��Xc�j��NV�$WX_� ��<�E�V�-��%�H⻰��}�+�o��������Y���Ai|H���@p�Q���3X���B1^��I�>[{!$OC/�[�y��p{(��3b�'�L��)�>S���[�&�]��ãT�a��k��H��g��ϐ{-4�a�C}ی]�`}j�*ff�o�0��L�����Ə^�����z�����]��k�7kA��t/���R]�U)��Ͷ #�`������4R{v�3/��fa�?8;S���2j_	�<�ކt~�T�^��l���ơ�MӠf�>O��Pڥɧ����͛�D�\�O∐��l�o��/�0���&�o���2�N��%�f#���g$ �m��[��d�$���a��\�����;��B��,
Ї)� f�.{�N�J��^ש[VEE֎A�(2��(��;z,WE?>�=�����=)4$f<U�8����`�s`Y�'��� Gv澠q�CWb���u �l�E+S��l�ja�u�M��͇U��Z���2 ՝�'ItAL�0|LB�Tث�1�<!��U�����JJ���)�P��/��)��K�ֳ�O���z����4S/'��j�j�.3qϦ+۵��D����{�I���d�l���?��d�Zv� �blv�3ۯ�i�m�E%ga^���3��ֹ<�Y��T�(c�
2��qm���]�u8�d�,�J ΊD!��(�v�I-�<:f5xZ6�+P�H�=q �+?d�ٖ'�2�� ��k�v�eaukq;�5\Sب>x����[g���(49/->m*r�SĶ�i!'!Gq<5�2Z�|mJ�3Pܰ����%Jn,1l��7��R3�T�En��s�l7�m��lly#ih�)�R�H�}BHD ��L;=�kB����<*23Ūǣ(,�~b��[B��J��`��l��o�Zx"�����B��[��`�@�stj�W���Xkp��tQ?PPv� =t���ψu	!{�D�P�"RZ�*c�KX;�&����Ŏ���<r��}�i�>q�5i��(u���O��BU&��̎�i�1ot�ʹ��k���]�����>h:$׎�bx(	Cm��u�sX�X�e= ��ԣK:�,=��#F\�|���I1�&'�`���'?����gsڞ���T��E��Eh�o������.��&nE9b���S��� 3��������u����`�8- ��	tl�_1�|�����C1����0��>:ǭ�)�ܽ�
�s�����G���������?(QO�E�̧�!�s��3ט��۪��BM��?;�A}mq��l�Kh�I���"�`l�#'#�3��p���+��#���x��3�N-G�!�6�ř��W68�/gQ�9{�`��F~줞�F���j����~�:I�lro�T�O�߳u�!��N��D����������<of��a*��>�o@�G��L~|�����qE�!�Gҡ`W���3�"!�� �7�����v;��'ȯY�4��T���>1����#����~v܉gM�V�>I}F���n���*��4�CO9P�k���0�����~Mb��4JR�$�`������ސ���%���i\����M�ǭ[#6m[5�eG:赅}�͕W�oF��@���H¡'1YLm%�#�	����˷��]�9���m*������DQQ���h��Xt*���	�d.����n�E�0D����Y�Z.��i�a���˯v��<�L0��Df4�(T7�dW����(-���2��HŐZ#���λ��hdɢ(<<O8�ز>S�(|�:�Q(�`#�J�X/=baH8	#�<+k/4���1I�)總���p����fջ)�n�<���\q�BZ5��4�4`(dA`����W�Q�]�C�����7sΤAH�a�t��u5��?�-p4Fc�����C3�^��A
�'��'��B�_2B/�<�{aerM�}|�N����{ y1�t�<��V%s��Oq�7ɽ��@� b��P���� }�����BE8U^yJ~�/hf�ZopM0b�cd!E�
iO�.X��o������Z�i���h�s�s���k���YC݄�v�W�U�7�&��F�ϻ���vl��Z�]����M"�N��%s�BQ}�)!�������s-�|�LGa�ؕ��.�\n.D=��\�N��o\���OctG����me$g-��ξ\���M=r�%Z;_���ƨj�p� �8��%I��8!x8U| c]B5�c�==�hES���u��E�3Du�Nqd�`�U<����Ҍ��@��`XǨO��a��>{u�ƠP���8�o�Cr	$���rb���6�ah�ND��m��lgxA��t�%m]�m�J�!8}��\�]�Σl+סj��zAt��vg�%$��)3@��z�-����C�4E.k��Y��Ŷ#|���Y�U=����8A
�
��㩣%֟�rˡ/v�t"c0����U�kb�旴��~t�/�"��d(8�dV��7�ĳ]@~M${��@*p,:�C�y``����@9Eh��1��oo�M ��	�(���X���Lm|�#�2�8mѴJ-J�������#�	����CӞ��g��U�,#bΦy嚈��;�\�!�RsTp�7��4���
�EK;.��q|5�>��?t ��f�r8�{ˆ����##c�ͯL�*gǟuUpr�_ Xg���ݠ�	��Cv�X��IR���H�#q�\�4�v:o�c!��1��Y�P�8Ѐʽ�L�܃��3�Ї�
E�P-�&fBYAo8W��]a�u�ܡ�n�����>1�W���X�5BH$��G��4Ʒ �) � D����.r´�۞�˱�'���`@�-�*,�|pk$�N����B�z`ь�;��^~��` �� 4.VYd�*E�׆\�Z犩Ж����W,���2U�f��g�Z
��F�汈8R�^���˩�.��BGq�����Ƿ[bK:�H�f���[^����Ć�:�)���#B`�Q�{U���=V��D?�D����#�|k�3C��B�m�`�0(��4J�ߤ�[��$<bC~���۷� ��ˁ̟%k�#��h]_�f&�ki�|�;�t7��5t�=Q�x�_DBk&�e�ҒZw@X���c[!�plWqD'����zN�eZ��x�Z���g�	���Si��.�u�	_FN���� EJ1���(���t��[&���{l(~��Y�iH�/i8�O�ջz����!ȃ�d��2���'{Z\=Yoݞ�g��G�#�����?ӥQ*���<�M&�@���n�XF'"*OӅ��fs��oD�"����?O�*K�������P�tO��prI�S��o���:Յ]Ƶ��0�t��H��<�)í;ԡ���u{�AϬ�/x���E�b����^'�E�0 q��:�N�C����a>���*�G5���I���]��>�S�3�!��W����ͪ-��nƢ!�B�i�o�wL��Z�n��vV�t�Iw�U��g��rR5��,�(-����O��Čr<e4���A�a�+Ta���V7ڄoc�V	/�8�lV�\�Qel)��%�L:~�Ϲ�qe��(��Β�/zvb����q^ߥ��}�ڔ3D��-�ф�i@YH��	�o�:��g+x0�|lu�G��I`��ȉ�] ��Ҝ%%cd�S@����1v�)��벸��IGY�pS�}�F�#�>�f<F7��~���Q�i�w����^�Щ�����oE�L��pȠ<K<ͱܢ��<5i�H-󤙹�ٔ���O���-Y+�F�)���dxR.w�n���\���N�s�)X>; ����hr$�^��k,{n'�݌Ynd��^���r_�T1˛�Ϊ
2�?A?ja��Z`�2����8�r!D���Ym�/���uBe����j	Ƽ�a�עNяR c�I�*l��s�E��t�������hӻ���W�$��䔌���:{�ֱF�@���lXi�Hl��z���ڝS�3?�_��