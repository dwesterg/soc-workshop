��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t�Ģ�H?����H�Nʳ�d�[ii�Tr���XH�����%��&�d)ɻr�x!�]#d)���H���"�x��8"S�+h/�8��:Вz��������-���@�<�
���m-pi��טʏ����|�q8�Z8G�ӡ� ��߂�L9�����O6D��u��ꍛ�=x*�ٱ��qiJİe ��D�X�T���[�D�����Tkpٱ��dH�&��FA%BF�|�5��p!����K���S�� /��6�`ܫ�����3 P�B�((����v(���`�	���IlOC��f�[��:͓ᜭQ��CУ_��+U�5kܞq��֨�e��Š�|��x�
}�^�"x:e �EI�Yq����=\�̂���T�z��Nz�����QD�쳠�� KM�m8��Wc6X����2���kбB��Ʌ�������ș
=�
�y�[�`̣��f��	���<��u7���ӕk1е�,� 4S�Q��h�e2M�$_X!��ۢ_�`�|��d�H�C��Ή]�D#%��ri�����4��.��,Yl�S׊��
�s�6 Tq��p6�l���u���B�z 0�(�}���l���% �%����2�1񸙅;���!\�fM��{���ܒg@�ߦ�"qvHL���,�v�P�y��v��R��	^[K�ӣn5qT}�!uO��}��h/G�T@�̜�F�w�H-y�<�
�o��{����u���1�1'w��_8d��_�pE��J���Sf)x(>�tݝ=�i����F�<����8�7T3��][>�O'7��$\5iQ#���yR��D?�'���jio�?��a�U�y��H�������ٌ�d˵|�+gL���2kJ�z�V�_ �"?<O]ļ(�Ы+2����+�ah_�k�F�3JMF��*n���u�R��|C* 0�
��(���#�k�.� ᨒ�����p3
����m;#T������by���S!m�p��-_2��@���G �@AlT�&�g���@��(h�l��u㯚��5x{2�Br��( �gFb�A���_�3�#��h g����\4��s`������R.+��T����P�W�GN��o��9-2�/�YE���E���L��%��<�~����ð&����6�h�՗����T j`��65Q�T"����Ml�蚴�k���,�;->���s��bj2���XH��$R�
w�E�ɦ4K6����U_��a<>��]�dF\�yFE��[�t˚Ht��6���x(Q�V�P�-�e�>��%��=Kx`)�d?4ij��yw�4�>G?V�dׄ�mb.�
T�~�RA"-�`AS�f���O����d�ͳ��Y��ܻÊ��1�sY�M}�h� ��t����Y�ye��6��cF��	/�06(�ę(������l�ԑq�.?�5����<�$R���Z$�/�*��+�:�̪TV��2G�vU|H�V(�O����=�[�{��e=6��؁�×����Æpt�@0<'%����ٽ��c�X��U$�P&g��?�⽛p�jQ���k���� ��猌�B�O����b*J"�y��s*�s�@8�^��"4E�'w�rW0��@v���jcX�*��"d�D6�]!<:0>Q�������64ŵ�w�=؟7�
�n��Tx�ZcU\�S���kP{|�l6ƀ���0,	�7tF��2*��b}�0��+�-�b#[�9Ϻ&83����e��=�9q�-��O�	5"�o#����ID*������\S��ɍ<B߮ܔ*��<=�gg`�jg���{�}��N��g�����jb����e�����Y�IT��j�����/��O����M�5p���c7�75�hA"�5�ޟ׀%=X���N. @�>�Qcf�D���A��©�<���/�D��rI�3�5�����0Y_Gq#�H�JSӕ����jc6�i;�~��=�Hf��_��*K�i �K�
�yL���-��K|&v��ph'�=�fI@a��7Ҷg�����h��p�`���u/%	*DO���qb���'�Ȓt��T|�� �P/��������o���M���{��qoy$_� '?��"�tqF�Yr�	<7;N�e#��d���$L`zw��E�[���GZ!״���~(YC�Y��x�g<�v�Y�f.� �����/8�¥��K�(U��}KDF�$�s��������Qq�kB�����5'�}��j�[�+��z�ӟ��xCs>��Ɉ� &.� ���S�j.��$� �1ϓ�+tkI�T������q�.�)KZ'JY2���9�_�2�g� f����﫹o̼�<���+�/��ǹ䊋� 9Ѣ ��1��<�J�&w�Y���Ci�	\dk��%q_ՇA �`t;���z�:G8�p�Y[T&R!�z;b�;���|��1��gD�$;�؉A�;��*]������R8�����y��k��`sd��EMK�N�"��
�T�:� �E��d2�
�џ�hl�Շ�\|%�=��j΋".8��)ذ-Ҥ	�5ԢbU�s. C	!��k�R!��*��﷦�hM?�4�3�H���@���v��6(�˽냭�#�,�▃���z�=v�:D�}�L(_�;O��Q��YΪSY�4�)�{�4[�)
Rx�ݚM*�NA�2���~mO^ ��Y���y=ug���#RO��V�8g���o�;Q�d�0�t�bQi�R��?ʙ���+�6��%,"|W�t7ଌ��)qM���
 ]Oǽ��	v��$4j���������Jh�������0�#3R����	�y�N�>U���%zQʝc��n�6�������U 1:3�������BE�5�z%�="�´`'��}ъ�j󱨫9I��
	SiBd��kI�n��W�,Kxr9!�N�F<h��J�W�M:�d�'C�S�&�8�蚞>�{��hE��A+�A���[N:T�x?ʸ�o�r:ᰱp�4aƭ�Bi�^�}Y� ,_J搳r�ƹԱ��#i��%#���&�� �!&`���	&�d�md
"����0�2O��8��1%�^�����k��+@�aT�:tD ؤ�E�=00Y� ���08Pah7W��߄����fS��=/ (����ʾb�jr^+�|<��P3=g^w�y���~S�,JZr���܀CJvaa*"G�p�5A�z,���(��a�&����϶*��д��A�T�u�Hh��Az-*@-�i���Rj�ǧ����6�h�;�ǎ���:�A(����D�q8�L&w\������zX��h�37<��QJ=`L�ʹ2�}��$��1�b�%:[�4�nV��Ȓ�-�Qⷂ��M�h�&[��%���H��Oe/	0���H���%��j^��.��B�d���i����������F~�
�I^�� �Xw
�]NPv�|M�T�����Kޜ]%D���CZ 7���ot��ɎX~d�:���D69�z� ����|.����-��3+�#��	�'8"�w�V��n�+?�$I�E��Z��I�J�۝l�8�	h��ù�Z��@Ab��tW.&�=���c���>���%է�ĳ�뇆V;HO�?L�ٶ�׸����.�w��-a'�f���@+�D�����i�7*ʮ�����8��B
�X|g湄��(A�tp������h�i�aO4���D��M�����c�IS�N?�i�v,sf����%d�)�չ�R�bw��7�]���|�jŏ�e%���������ֵ**�(�Ȋ:��L�1���&�:��Fl�x�M{��j�ʴ5�#�+%�_�u"�OE8����/a✇�b�	�֜;�,�2�o��ם��z�[�;�a��38]K	uّra���$�y2���2�Gzx���(@�2m]0K˷�:���H(�q�>��%/e���s�#"���ק_�@�œE$�P�}~�� ��w�3FR<a��a-K.5	
��� ��
�6rem��H[�*Xx��tL�����Q>7��<�Eg#��3�������b �0�����r�����C��(�؀߆\w!�P�����+���`�✤��� ���;_��������sb�MbJ��E����*������^&{����:ʣ�8�m�|��:M��WFk��=Md���cB���ԩT���fn�p)	�Oec$V�����C&�%�#:�tn�T��l�O+�^`����|8�i���G�=~QP�HD�.O�4��x7���=o8;�R�|lo������8iS�����=}�Ӱ����f6��TDW�}A隑�3��A��`D�!�����֙�ƝIK���LtO`���B
ba��ꍖ���>'�»��l��,0�#,�4X}�g�h]����?E� ����k=�!�I������M�܆ ��/�U>KC�1�~s��P�5�d� ���#�V�S���$��0t���r,Seq�H=�*���R����:�g	śdĭl��)���<�]�a�d����^5���F����/��k\Ô/��yA�����=IKz���s�S���t�sZ1R�0�b!pe��g�w�{�rQ����ٙ���#ki1m(K�6���x������N����'%���I�I��h�:�rw: 7����X�@��k`�R���/}ǰܭ���.u)�,�?��������IQ.��	�y<�M� )ꮶ=/!������?̲�i{ଌ�� 9�v���	f���뇍�U�w󱥛8��+�#�-��G>�H��	�6{�2�iz�M�/��+�l�hj�9��#o���]��⥼VsD��g��)h%���a������OC���7���6���̍��)���/D)*{�9�b\�RӚ1����8!�|����c��p���*��s���&���ud�_N��\l��}�i���(s;��|��C�E�j�Bτ;����{(�@�~�6�0�{�RU?�mh!9��^y��6�ۅ
=��w�@ �k������w#��a������V_�H�7���VQ���Ge'�0��8���s��bc�m��z�8g޷���(7�A2�_�*tL3�T�2e4��[��`�}�D��G#����e���#��Ԡˑc�v��6����b���J9p(�P\͆�խ/G(8=@F��+lU{��0�=R+��E����T�m���j����L�֫�#t~�5�O-DY�u��-�o��j�5�U�PO����#'��G~?���7|��~4�,�3���l�ԕú�#���Q��c�Ly0k)���G�+�-Cn��o�8U�F������z��,�{g�{(�U_�P�Cg9�4[�9憅=,G�G��]>���Nr��/�iZs�&�j萖(�]��v�)�?F�9�P�"t�VCUB�����^���@�����r��vʯz��.6��c6�م�0�މM�}�F5���hBo
�_3j&����U��������m<�3��q�}"Z����0��}e '�������3XBp�N6	�#p�3�/�6Y�^��R:�l�Z
v�s�a)��sluVxA��6N%�?�.nլ5�c�q��H����s��O���C�؃^h���3����m%d��ț���c�<�Ej\3���s Y�xX �9N J}�	KP�v]m�*s���/T���C�mB��匢�IZ�mF���$�t}G���aX�_<>׿�1'����<� j%A�f.�����>�M�*���|�qی�>��������`��� �V�T�02+5f�T�s�s#�Rq�U�վ/��nf�$���7˕\Ƈ��<sٕQs����޺xom��VP7\ �7vEYe���7J�f�*��1R�2�z	���8����Pɀd�|O]�*��VFnP�v~Kr�!3T��i0|za���"G̞)¦��Zt�A����>�"�=�}so~<�@��^�!Y�R��[}%D����
%Ԉ���Hu�M������J$A/2/��1��3PT�t(:��� _y�iS�Lq�"�R;fQA�O��`
f+�M���Cŋ���N�<Ĭ���Ѯk�y`�y.w��>Ӊ�5�cC�"����k}#*4��V��}���Sh�/KZwV�#'�hu�;����/��=�K��.y�%r��`��n*`�5��*��Y Lw��&�|�V_��9�}@�@�E52�w��e�A�c+Dr��6Q�E^�SB�/E铨�Ͷk�e��.�v=1����f�<?6��R�_�&c�#0���hZ.P*d��e�w�8��q֓\�]e��3�s,Q�cbyc�5�u�̀�� _��c&C���4�lDV�Ւ�A +�҄uP� 0���J��xX�nW��.n�%��9e6!�����Wx#ԭ^���'�*�ܐ���F�%@���P��CR�q�ix4a�}G
��9��<q?w��ߵJ?�X^�C��)A�H6�N�Zԉ{oը��En"ɻkk����E1P#1�J)�M9����mI�hz��c"�,E���X�1٭���8����@}=`�M�a�G*<g��6�ڟ���������F�Yt!�W��A�����r��?w`u�%��OA�.���:�@#�pR\����r����\��:��{t�!r*�F��n�Yx��bm =�mU�{15vh���aq�� ~��,`s��C}o�����Wr�FF��k݇P ���Ac�j�I��5�y�7��X�\,ܵ���j}�������^QҞ�R��V5��g(~}�5�0xD2q��`b�����b]��ˊ���3	�;�;��q��X��7�q�A=Oq���ӛ�Գm��1��1Ç�jQqJ;ig{������L4���Vɹ{�;��ճBK`P;���"��ʴ_�?y[;%��8�e��p�S��_y����I�7i��o�5=����t.ր�5��F�w���_bK��=2�� �5;:��D�3��\qw���Fj��4 m�S�����ɗ*ǪO;>5�Ϟ�C�u�M���F�8���z� ��Z�Ƅ։4I��c��g
Z\�����/b!�
�M��Om��ӂ�l?���uL�!��C5=��E�zO�zvp�h�VP\AG��O��w��U�`�6�����g�ʣ1��w!1P�[�<?%�	]>��x^W�b���i��E?�h#����w�M�����\�,(�Ą[Lf儅'[ن4-�l�)S��������4��\��z#���Ź'HU���c�0�*o�'�� 7��-.�RIf�����]��e9BC#6��fX�:����r���  6���J�`CT�8��Rh`�0�kU�2���@�D\��*�X�h�Q��-P������%So��|}�;����I1�tD�٥�R�|!�_L��(ڦ+W^S��V�&��Im�(7�9q��]��a����8	�F��+��Ҟ��`��	��}>��E�.{X�Ê�:���>_����5uz8�e�u�*�fw@M:;�K��jiZW㇡�T܈ߺ���@�5 k(�me�!�W���JW�q2�2��.:�=�1��y�w��ݕ�����l�W|'~��pחY�`��u��l��U��G�Y�6��y*��+L�5�U�=ʶ�2���3�zu�i�$���X^۬P���1��nP�U� ( ʵz�(��n���!ҧ�ٱ�+��(�A�����K�F��i9�^x�����PW��F���}����uCDg��w4t��kW/
�ӷ�acAu��2�z�s;_Ҵ���d��^";=��~/26�����=H�X�%q�lO�^(�\��N��	ݡ|�CH�P��Bþi��F�K�m�X'δ߰�C*���TQh6��b��B9��PA,[[�`�"���^D��Sy�ȺaVվ�*�R6w���N���p�1w-�A��9��L�p��f&Џkb��.�쿔!��u@ROy��m�%Oh���������
��>�6zC�4�I.��DJ������$����e�QYJ-��9u��Jδ9i<���{!�)��:d(�i��[BNi9*%������$��([��Vb;W$��;�����+R97���3iF�0T?�*\�����=^��D���*���lZ�	���t]M½�����y;��O^�a�a������Xue��߫�H@EtV#�T����9# `�gG�:��@�t.��$#l����<l�Y�>�T�9����i�1��_�0n��m�߾(�2�b~�F2H���X��z��ĝ�*bvE���I�I�8r�d����{u
�y�(�a �^
 _Q>�����3��\)&��r�$Y��4�t��+L+]aZ����}G�0���}j}�w3!��c�x�FA"]��{R�ia��&E��WG�k*k��ZR�,4�H
"M����~�� ���cG�v�z�x	"�"�d�s�����L@^�ǙI�mJU�y�P����ϳc�0l�>	Q�#^K�b��˦Fv@� U[�w��=%��$[���y����!�� �u�B�ۀ7-�����E��v4T�h���i��[�:RD����h��\�w���YBsB�7	�#���)��	-��칵 ә�ܖ����IV��Vj�F���W�P�� N)�Z(� ��e�-��&�u�;rޏ1��J�M(�=:���1CPJ�.�o��l<S1�7�Yo�r���*�����4)�E�7�,^?G]��5!(�+�
������-C)�c���0;}P^b�İ��L��R��o�[��+��3���7���>����e>hf��|���E�\����X�԰�̝
_\Љ�'����vw��ls��$Xi9!��9���ЫszT�"n:;O����>Z�8TYK����ԣ	K'�$О1��MvZ'䞙�ߞ5 �sʓt�N~w <<��f6�G�5�����oo����Ӏ�(�h����8�3�yU�ś$��w\�^�[3�#Fз_��S�K��it�/�h�$G.:(]�j�ޏ, �ݦ�I`j�Yی���3N, vZ$�4��ɼ�Y$��U$\�y}bM>�<N���y�i�N��_�B���Q���.P��/�d���S	Eg�V�X� 3�5�����4�߅�m�`�P;3���kb�+f2��U���.��B}W�m�:7�=p-,B#y��$2�?B���3z�H^���M�@�����t��� 6%,A@<�x(Y+]�Yy�1F��^���;%=���u��H������3.��
��DH���B��	��!}Z�qq�*�����YUVF���(�::�>�)�H�?Z�V�]�%���W 8��I���/sofA�KH���'�ν�2��x���}�ڕ�s;� }��LgR��_�Q�R�I-�!-钅>�F��[1�-�4�L�* R�R�29�L@�.	����2
bU���D��H7x���ݫ���K񝐯?9ث�^��ɱ�.{.�;�D�o.�ȖII�6����Ӓ}F���/ԙ���eA2K�m����o|��87�	�i���% ����4{�е�K{�)!�)�-� ua�F�FZ�w�OӅ�tk�T3�˓4�V�m�|~<�$aėR����V�]y~xR��I�)掶C,�5��I_Vx��#��	�#]g�ci�;�9��:ĩ��Y�[�v��L��0V׀�tD�q����-�?k�=(�n�I�����4��a����$��5H�+�j����jABi���ŉ��ȿܪ�4R�m�L����� 1��p��|��ܲ�!z�MUP��}ab��n��-=��.;<�	e�؍d�Ml;D�$��1ֆ6�b�\�/�[�s��,�rϋr?�intjn����P!hy�}�9<��K�R��z��3�_�0l�T�{����^���APt���~����K8r�I&�50�H{�����a��Y<�m6CZ��Z�%�܇�.;yń&�$*f��R����+��p�\�|��Rq�8��Mf��5�Tf��.�}�Z�F��E��ͦ�GfEIq�K:i.Z�B��q�P�c����Z����r9jrFw)'�{(��������t��Mv(��»��^)�.�Y,�E�QT���n�z�1�3�#u�nC_��l-X����W�iH�or�\��<6��oNQ��CG�B�t�]����#|n-H�s��(\V�B�a}��\(�ҍ��7��m�r����Hdr�����);ǶV$�������Ȑb�z��h7L���{�~��h+Hw|�e|�XE���AL�oֺ���'4=���;OV��C��'�*�ĺ����<�y�\Bߚu�u��Vm
×>�������������d?͝�R�8%��g8(r����`����=.�MU���8d9�j�Z]���rl^�f�#���e:G/%�6�f���t�3��=���������Ɗ��7�W�^�G�>�[�Ѵ�Ŝi�J{���+���cb����$sCw*�':yG��������:�c��&�9¢oQ���ybpB���G$o���r�F�ϋH�S� ���� D^�Vшx^b����tf%��LC�E!z����BL��^�����Ɂf� /l���0�(�R�4�#�:fo�C>��}Ӽ��D�_3c?���EA���4��#
�n
~�ƭq^���/�XX\���}���5�p��[5V'�Vo�T@i/�^��+��	!��_��(����>��j�e}���N��t�.+r���\���}�u|�N�n!H-��x�ʻ�L�ж%qP�DJ[����>��e6�w6w��F�g�k����da��� �N����ˎ�QSQ�;m�O`��M)w�e���*��� �/KY4I���z�I%�y��ӱf��$_�d�aV����lqx�ٮ�i�m7b��b��\Hj&�܌4�S�$�X�qtN��FS�x�tr�[�[]����ɬ����eU��nЮ���	Z����/��p��쨇�����b���=M�U���uټ��� R�4S��A+!�(�6N�>�����פ��;��,�7��R�Fz�O�L�xrLbh��:�,�T� �K��֖"�HȐY_�9ВZ�8>�n���G�O���G����1 9�y:|Hޮ�!�����KN�t
�+^�(��Xa�{r��Y���`��q�[��71�g4��8^߲<��[A��[�q0_�=tҔL�]���}a�Q`��==�L��?_h^�=ʹ�{��|BoH�U��9�m8�f��-O���Rdy1�e�"a�C��~wW?�Ic��O�k3]?E��X1Y�Br)���w�?�>`m5�Ȑ$�)�ٶ�ߓ���;�.>(��2�x=:����ݒ�cs���h��;ـ����6h4���U�M�+0KV&�o�XzC!��GT�{i�H�,wp^�*U���Hlp���֐O�����>�!о6�R�Vܙ����q�F;Lꅧ��dm�t���� :Fo���3@��bv���D<O����E ��\�ͳ��[I�W(�h�
�j�]i� �24��3gƴ�Z夾��nۼ���0K�w���<:O�ڂ) '����N��foG�,F��E��� �bw���H��*�C2�.X��:%�#�N��LQC}�06����0p6�dAq;KB�ѡ��2��X/�0���Lt�0y{�UЪ��MXz��Bk�M�E���ISڪl4O���=è	p� �j��R��sR��1��i(��k�6��Lr�$�6JV���s\R�d�ϟ�عu{�C8G'
���eQY��^��be���to�s��U%��yS�qi���M���,�:�v�<����k�)>Ydm��3>!��}$��B�V9됡8k_u�#��ړm���"���;���9JKV��I���tH0�Se1�6q���j�ڼ������k�v�h�IG�_!m�@;+����  ��&��.�¢giy"��g\�q�uFV��.��/��%��]���<P�A�z���2 z�v�`�0v��g%~	�D�e#O�ɷ��|��ҋeЃ����)fò$mw{�0M�KI�b���x��-:����
4U��htɑ�X}���ے���~�N{(���������h�}7`h�g����������f`LY_+"���>����Z��Z�ՈX��8	@٭���k�̿���>\7�N�`��8���i�$�5��Y���P����F!�ʢ紻�,���/��p��#�Z���<�^�x�$�� ���@�`g��.������y����GPS/�	��C-�?0�w8T��:�p��%�z�o3�����6蜛��\h��H��?3�
�D��e��������\	5O�v��Cv/r�Oq���)�gf2�߫�J&pB���S,.s��i��c�o��U6N���\{���Լ/�p];�ns���&,��[����|�μ�)�z2'h�wN��[_YYx�'s��[ZR�K������qm�k_�O��f=�oO,8�����*Rh���t�j����M6݈�P�k�d_j
W�h?���\(�Y�U�p�n��[ 槢��A��u:P۳<	ʆt��$������#(�]�)��1��`��en%q��{��i"w��C�c��n�@�tU�`�j3捣�)'�Bq�GTK�=��h�# �.c�C�݀�#}<��S���+<�k�����ͣ'I��j����V�+���Ȇn7�C�-� j/F+�7�T��Q��d������2wґvz���0�D� ��4�����-m�h�������H�p�it�&�#�k����T�H+�G}H^��i�,�NtR!�'?��y�6�W!�G��)Ui�ʡ��I�M_ͳ�1���u,I�h&��rT��v��BB���K���_�z�x�Tˡ�
�}��W(Se�(���MV�(�J�8�Jh�f��Q�=��#�$�$��Mv�=��<���G�畷�)2A�O���A���C��]�[�bT�(|��-�>e����)gN	��;�!+4wf�ӗ�Ƞ��}�c��N�r������tc���+	����hs��o�L�	�z��������H~@����,+�!��S�m���q��̿c�Tc5�{%���:��X2wM�S���a���4�IIW�>�Ҭ����,n�R�4���$���ac�Z�*�p�}���r������x�3��c�y@�z8�3�~C|�#��0����W�gFd���Z���)/��Q2�3��.��\T9��H���͂X}����v9��!�SM�i.�b��u�L�'���Zٽ�3��Į�(~=��?�QJ2��B���酋d��9� C�e���N�Z�9T��� a�	Z��6C�nZ�Bfn����߇0BE�^ �?!�ѕ�瘝�G��=��^aP��[���>���U��r��Z����}����y;B��x���R�O�V}d�:Ha���k[R����I@K��Զ�A���6h=�T���}�f�)���?5pg~1����:/ac+���]��HX����qKuGc\��=�H�'���-o9�����0Rj�${��;}���	D.R�+JNǤ~*�����y�k7X��7�
� cjAb������w+�R��?�}(��ֆ�/F�D"o��0w��ѕ�&<�!��.�	�ͻ�G�o������M���T�%��7iK;���	��65�"h���r����wϫ�(r.�fQ��Fu�>�+|Cǻ�po�����qDt|�-�AJ=���񞭦�k�AHvt+��g�nq�U�#�����NaD@M0���e��~����Iڼ�1kk:�,���c�P�3����r�s������
*��f�µB���`�|�6j�.x�02$�c��<����R
��fɒU��jx@�J0;�R*`�/��9S�roF' �B1��c�3kݓ:��'2֏	�B2:~��R�@KݚɜJ�8���.pF���{qG.=�����P9š�SI�F�� #�V9��.�e[u���Ԧ_.��l���!5�ws��Q����v��������a+����
��y���ɴ�@������\��d����B7��9��~������w�!`��s�>_\���gq����XK�1���RbDh,G��U%�Y93����Y�.)Q5�-�B����1��U���smY���g;&�ML|�֧8r���^�;�wmes�=��`��O⠔@J�n|�$�7�������������e)�蚃WT����{��H�)��r���b8L'�92���H�n�4j.Pm�z:��`�xY���Mi���o]ԦO��p)ȏ��[1��������<a��1ڂ�-,��akl���������O�(�˨�Y����w������cY�!�"Q*?�ɪ8�O_�-?���	A�)_�:���{������g�q
�ewQ�Ӯ��0o�$���+<p�$�1����/�$g�:YN�.d�D�G�B��Ž4.�J�!�6���U�r�Y�����.�/"}����
���V�T�w�g��muH�,�nu�;sO�H��_Q/v4�_a��֒C�r�6� �a�9Cy�x�6���f��_|��Y5C�IJ�Yfef�-�o� �M�]a�k�O���[����J�sBW���u�$�D���v3+]�U)���u蠟��bOT����B4H���+��ɬ���Gn�t$%T~��8fy�^�9@��M�K����4>M��Se�78H�#9*H���|�Nx�����a�$���(��([i�nr�R��ż����2i�J�~�c�����L� ���n���y�$����{K�%��n����pw|��M�cF�V�-"��|9���5s΍�6�εߐ,f���?�x��NNR��#��vj�1d=�L�J��9x�zQ��vw���3��r�.k�t`ڍ����v?�V��ID	U2Ĵ�K��$�A��[c�6'	��K4_Hj��<Х>�Bd��׆O	��S�ѝK�}:.�ݓA��=��������~������ɲ[3sy׉���i�LR�ˣ�Q�����\�K��MP�dJ�:2S1{�T��U�)��6nq����oN�w�(�~�+'��Hr΃�d[�l��'��a��St����7_�:3x^fm��ɏ�R�\��M�j��J+y�6.����j��-׫�����\�/�~���(����z�D��9\���a�"�?����}u�z4�������߲���[��t�	�o�����mY���i� �X��̀�7���: ��.�6�� �dg�Q����QB�����,��(p*�HC������u��#�@0.Ȍ�r��M��a�@��z��$����������mbG�L�����p��e|e�M�Ơ���Nk-����lUa@�+��.*�3Sl��̀�?�>����,���Q�A�S��X�vYV��Qn��$"j{E��dY��\)%w���S���$��MD�՛���c�����lʟBs���H�g�ޫ����x���qJ	b���H[��;tf�mSH4mDN�������g�EOj	��n�'%ϱc�$�P�P+�)f����]��d�;��P��
	�LO�#��C)�L��+o�ɛ~�7�]�W� ����s�����p	v�մ���)��I��2Ed#(�@}q���!#Ȁ� &���)��;A8wZ� &���x�� ��)��K����|G�k�ȈUۍ'��&��O��Q"k�q���ۭ�S�>	=��	������/z�A�_iF����~j}�α��`�|���b딕J
���q2�
d#�����6I���8�ڊa�9ʀE=�U��7��1S4�Ҁ�1�^Ȕ�K*� tl�',�ò�^.#ot��!KY���lt��������X�<J)�����k�"�Aү��ڽ�\%IGRpY$8LW!p���$�m�/��Y�S��]L��x��:�F���H��W�n���ns��@B?z�R^s�_ޮ�*+}l��w�{J��2W];`'N��:�`�Dh�hi n�q��ݒY�]��Y��_du\�>�� �:C�?��{ f	�"�n��sr�^��	�l!�?��Ao���ix5�}�)�7n�K�� ��
�j�����c,L����9�z���/��1;��V�>����'j��Jz��ee|#o����6d������Z�+�>@&��La$����,c��V�ҹmX�vt�oap��裐��-�ۼ^�`�>��������4ey0!p��D]���T���@G��(�,�[�!�Ky�O&W�*��4��Sr���'��G�k���?V5�nI^Q(=��
�qvB�ܥ]o�=Tm;`k�>��E���r:��.(;��af�:�*�h:Gd�N��dl�M�f�bm]��^��d�"8��tKޤ�I��{圵�N�Ãȑ��?�@yo׺�,�������-��=��8sU���a��)e��T��`('F���̴��HT*�%h��楷 $6��C�DAݚ�|�U��Z�=X��֖�V̌�gHp+?��r}�@O_w(�orâg�:1�OyP�9h�$�=�qC����oؐt�l��$��9�YX�H�j	��0v���B�,'G���$LO�˧w�������v5�~�F��ϕ�u>��1�]��`\��]��R��� ؓ��o�&�N[���kPsN�}�Yt���\nٿ�f���㗢F-���ĭ��f�"#��o��n����?�Ad��?�BW�o�$R8o�g��̽����Ɖ;x���7�3��H~,X��V"�J�X�#Gkf,�g�l_��G:�ՠ~Xb��W�,���{*�ʑ�%����Q��fh��"�e�.���L�qgƴ�C�Z'K=Y����l��_�j·��U��z�:'��y2�_�=�QQ�e�S���vG 	/W��OF��F�_e�������/:�v@s+5���Tݘ\�����?�}�����e�+Kڵ���$���n\26�D�Aj,F��DKK l�s�P}���=�k���2pp;���kNlB�TU�ge5aɻ����F2>��AX��%ʢ��zo�=KWlM�!�HL�����兂�nF�Z�02H���d����M<X+r���:F+���g�����l��n�a3Thm�z��4�(z����s�J�0�YXs8ɢ zĉoȳĶ]3M����B��+=���)�ci`��_����<W�@/D }i�d�D�Lئ0)$�h�������X�g"�>�WN�pH�J�,��(�w����o �)�K=����Q�3�t0��`N�^���`����b�G�2��a'I�>�vArQP�Am���4�!��O��i$��{�D9��3ʃf�����f���b	`��˿�Z1�=�(/7�у��
H��� ����?W*��V�����by��˙{�ђD`��z���ā�]"��������c����=l�u	�EB������^� l/J�GV$k(�U��7
��:v�jF	A�
�(I\��
�I�l��r�`C2�BĨ�����y&�.�	��i����wǮ�;5������r��O���C���g��D`ؓ��_�e��N�Ɂ�%��ojf/����o_�Ӂ��0^K�� �]�?��A��Euy���m`��ē�7Ġؔk���h`��;�*k2P�_�r-� .k<cHkhD��zu��
���!FQ�fn1_���W�^��b�Lyh���~���.�w!�2��W���y���Cݚ�a��>�{T��K�7&���?���4��݆�,��]���u�~��j>D*�锱����_(�ҳ�}�qJ�Dep�?�o��������G;�c�w��'%�w42��ڸ�f˓�� �3	��`��3�`�^���A[ ��Rކ}-}�����v�L�%u��y�<�YT�lكXQ�������<m�FفLHYsZ�g�Y�+�.�r�wղ�t����a3���E��<JQU�����
�a�b��VmC���l�����-��ܡK���k��$Q�U��$(Jݐ0
����'&��Ib�a��Y�{m�N�����\�&�fK�7�����7�3�6�1��:6H���q�����I���7	0��̃K���kO��O��*J�/�6��\-�e9L�q�����ϵdFK�w�Q���5�V9�������O��K0���� Y⓫*����8~	���M?��;���Ίw��
N���f��G.��0����B?�$9l��B����؉/b�z+��]')�<�����I>2 �I�(��*�pq���{��ET�^'_?��5	X\�μ��ن�sB��7ms��O�����l�qX���Q��.�W��4��_�r-!F��\1��2�v{Q�n]3F�c�V��Mr�����Є��$�}�����~1�'�}9D���(i�?+٣t-�>����j���+�����թ͜��X�P�i �N�2�L1�N ��+Ba7����2���Q���0Д���k��.�<��cN{EXiw*�l�(�VWm��{+��aR,�a��t2Qk���X�y��4_��/54U���l6�ao�� gs�;S���m�
I��'K�{���V�o�.F����3���]u`�<��KV�(��]4f`�m��lo�h�j2 ׶�c�6].q�1!5��Í-�Q0�WV-���[�(�h$���-GS�@{�����LO��f����傌nj\���ϩ?A�v���fc�]Z7����4()�zjN(Gh0[�Zn��<�$��:sm�׵Sc�ʉ)���+�E�A18Hō�V@�(Q�%x���͜��F��M'H<��7ݭM��~�G{g��e�(���U��~��ؠȴ��R����v��6���G���m��Et��?�~��wٯ�P��+F)t���I5�Gd &�^���#����e�(���ˏ9p��Z�;�u�8 ��%h��r�yy.��������~8�k���*Y��
��;Ⱦ/DͿʌ�zGg<���L�� �]�r4P@!f_���&52Qd&���7Y�һcԺ���T�~�]��,t�CT	=A�I��Y����k�@�0�ܶwL]��A�Q���1�;���ľ�$r_%u�~anJi��� �Z"x��5�jl��#/�t���4���q��8�*Gs�Js�T�H���U�w�D>:�B͆s'U�f<�������?��ٵ.�)�!2��1g�H
X��9⊚�j�`Z?	y�G���Gֶ�;<|�k+a|����U���h�֯o��Wm�������H��u�򪫢�]��(���^�i��
�)>���o���^����Nz '	�Q�B�#O�i���r���t�Os�C�"dK��N vc���o�̴;ztp%,�V��l���0R;����Oj�I��J���W���-�o��=�?�fy�BZZ�qB "�R+le�bJ��$����n��ɔ?|�_��BT�uH��*�~ڛ�{� buAf��a�D��J�W���M[�Fv-G�Vc�a�8�x}6b�98���3��D��}H#�O��qĻ7H����/:�qx�V��@���ñ�	�N��y�[���vK�2ڔ� p����[�|-Z�b�/�������i6vr-�ɕ˼��d PДn%"�o�9�?h���j�/<w-,�B����Ӭ�/�l���`S~����(�aq8zz�A �[�V��D�ҧ�_�ͱ��~[���	���I�є�Q=v��ȝE&2�~s�Z���� ��R�5$G�Th��_�Y�$��L�S�"��;v������N|s�R�b�Ck�\�b�8@��/.���	&n��g��'�g���6s$��%��vU���!7X��M^�������0�:�v$�s8�����>]���$yv�7�W�BW����!(�m]7�0t'���HN��DY�;�dN���X$Y��nX�a�I��~Q��������9���8u�*�*�	G`��`�,�:#�EB�z�S� ����ډ���RF�O�� �$}�H�\�
�nk.��p�֖$��s?�SiW{Fh^�@��q���z��~��/�<o��8�-	�S��~��)�|�,p�K�������9_��Gzg�wd8��o!�Z=�!KZJ�X�O9
v���G ��Vn)����lF7K��6�%��E�o�=^�^߬�Ms3׸	y��!5Ȫ�7b����u�.�R��8>B+��L�~�=�y� .�����qu2}�@� ��rEP�2�Z�]z[�U�|������0G����\ �t"�ʥ$DK��b��:�:����t�fd���péAjކ*��k�h�D�r�1 l��ɧ�&���
�?���r9��0'�}���`��'��\������������*�t"��[����;�0Tre�rfb�h�{��Yh���a�ҞȠ�PF�.�<�jy)�-ˆ���>��ni�!��%�H_�G����2�=�Q�́ҫ����YQr�q�]��g�}���r�s1
|S�p�e)V��qy��h 35*�a��������e���]%w%����T�ڬBJ�q�^�So��)-�F��x2�i-�4�QU�Ȥm��{����J�&;Ճ��7�2��D^�`@Q~?��\l�°Nv�d�X��j��CŨ{�=�e7�#�nb/��ht�B ��ߐվ�i���yV���J�6w�)��_?NŊ��承dįC��)5!|����?��`J����V�یD��ï�K��R'3�#���ʿ���ԏK=��n� �q妠7�n���φ�������� t����0|��)f�AGڗ���%3�Eq���3A>8S��P[�mcSm����v�[�]��ѩwTS��~�A`�$��z!�g�P��Hk茁a�Iq|�����;��j�VWi$byv�`?aoS�u�l���H���݇L�󫬵��K�Nָ�"u������7�B���������@�L�����E!(jq�4WKK6�Wɼ�OH����"��ɬ.��ϗ2��]%�G�����]�~^����4�pfVh_�B~��N��<�`�L�V�c�9Hv��-��`B�2�2bH�&6h�Z��1a���� �t����|<oTk�婧џ�{�Y&��K��֣����M=�c���6�0�&�o1�0Tы(���al,�v�*�����ÿ=��U8H���	?���ws���]X�Mˋ\?����r���&�U}��g���˙�����G�U�(4�H!AE��)�0e�ѥ����;����}�柆)ӎ��W��`-^o��o��遭gaLGe[�{/!eo��$��NQ�%�Ԕo?|��0�zs��t����At�D^�>L�m��7N�P�������w��M#���1�`j�Hz�� ��0EG>�N���c����^I�oy�V�<��'��l�T�%�n�}�(�b��sC�IH���"�h'��͚,I,�UDA�$R^�Ma� �s1��Lh*�+r^S��v�|@���w��R_�Wn~�V��b�6�ax������9���֙���Q�Po!�ِ �C��ؑ-Á����R�d���4
p]�a�Y�&�5��s��٘x��c�T�wmD�>�%��\A~���K��w��1B�ځ?��j�r%�/U��1�=}J�r6��ˈ+o��#�.�9������.R�<u��q���?\�Y�®}m�1�x�S#m]x1G��A5��|�s ��O����i�.���d��S��'�P�$���q�ZVί̮,�B[�aX^�Y)��V��t��h���
d�l��a^l���av E�a"e0�m
���VJR���t��YèɸR#f��|nU�/��V����&#e���|k`�^���(�� rԭ"d.MZ�����gl��1����j��5�yr���\������jN ��q�i5�훫OR��O,mU6%U�j	OD�p��1xB�B��-Y���Aiyk�~��	<>2�����(h~��<]\<ė)'�n�~<� �0�^�9��D(g�Q���r��[���v���@���9�Z£�-_��E�N6���Q4�.�\~�Ȯֳ����dve\�U���*#9�J/]Y�}� �쾖z90���A[���[��Pyu��Sޝ�n�6�e�U$���HUƴ+Y6"#�d1M�$�K�.x�=�����2�2�zS8P��m��N���2:Rh�G���R��&Jp�"����݅o-�~E��Ӄ�����A�p^Ü��k�O�H�� �v������W���x\ZD�m#���W:(���#��Q�|��nR�W��Zҕ�z#��oHp���0j='� h��jd"�A����-�d��1k�(UM\^梤�`��o5�v�^W?(&��r��tg@8�]<g�~2��ld������ƕ�'�;�ٙ&]������+3X��W%�ݚסO������]�-�Kɲp��v�0�h�ۂ�Vw\0�W;pV|��oiż@������c�1J�%��c97u��A�vio�e�E6�(%�ϡh|hR�`���EU�(G����}"'a&N�j'��U$�i�h�P����3�p�����燷����+7��i�n��ݟ�y�h@�q��=�T���W���k0�t�����A-w|%��Բ��Y����k]����\��E�۳��~<ؾMne���*��|�;��m�&�9ba ���f��sϜB%7��Q�y5�͝s��~�D����QT�ưuu���g\YM�O"��0�*]�,�4t>�r?�nP�ȱ�tU�[�`�L�+s�ą=�0�I��*R�W-�y@h�`EV��@Cp&YZ���=�y�h������`s&0�}��Լd�ݏ��ẍ�{�y2	S�^�5e�� ��ʠ�~"U�k���y*�TW�a��A[}���I��	���R2jRS]�2N/A<6SZ4�y�|2C���ˈ�WƔT���-�~W�3�OIW�ɤ5��UU�Ԯ䣆���,��XL��|��nJ�,?ʋ!�\o���ʙL�oDkyV{�3S���4�0����/O�$�x�^����O�3��(i�`l�x��5i9Yn�e����+t&:4��t�pT�����#�4x�4Fa�,؍�^�m��^"?�#��\&$��{��� o(#1�.�d���粏o0	MV����R�O���)tZ��'<`chL��;s��{�@��o��J���&�N�I��:vOr�\�`Qdn���ωJ�z��^,�w�̐�[+���)��J��H?�kGg�k1�����]���5uK����a�$Cx]\�;�e�ʪ��޶�WI�쩃tJ�oqY�;�u��ڞ/�u�PXD�=S�!�&X��ɛl�2��y��J�u�Q����	�YW�\�����P�}4��f�7�IM�"JPʆ=g�	R��������2V� w(��tR��$�sŕ����{�D�D��w!R~�V�h}���0`�b�-BA�0+j#2�ױ�� �e��!���2H0M�l�4U�0Vt/�Ô�_�d���W\ɭ��� !O��}�Al|�U$�C�@	�UB�~��ZA~ �Sv�}R�0oza�}`�2�� �7j��N��'p]I�+5-��C[��Q�?���OI; �-ۣ�E����0ϐ����W/��B
c���&\n{��ts��#�ؼ#Q%!�ӰH��M�c�����PB[����H�o�X�ET�Ц���ԭh*1ڔ�����l�ڼ�?��$��ۢ����#o�s1z��"���iK�Gй�`MgН~K<�ŧI8@�������]?��m�渕o�GM�B2�K�t3qٟ(���6a;B�G�3�����k[�_�d|�$j�
O�Jz��CH(Ue�J�k�M�eP~J���Ki-J����a�f$��x�~L�u�yu;�՞� �˺5H�we�ɛ]u&��s?J�`k��3U+v��������v��,^:�4�O�
�kXK\L�x�K[��x�_t�a9/�g�7��� �R��9L򡦤yp���i�����B���<�r= j�>���WQշ��KIWA8=�gC�&�����7�.��e���$���(� z�����x#�Sң��B�f�X�G*���N�|���/5�ri��@^ԙ��Є�P����J$(M�w	I���J�YF��e��v�򟫐��5����0�nR�o��%�7��b�o.`{qw��bS���A����E�|MĲ6e�h,��9�ݱz����tl�#���c%�y-tO>ӹ� ���?�	�ֺ����͞����;��ub;Յ{E��#�,g�OI�S���:ѳcu@����W�]�z}y`�M�'��{�B �O��ɖ����|vRoU��=�pH,�/J1�c�����=N���B�*p�O�y���#=3��V� �u��xc}�fy��Iہ�l~���+e���n�g��%�z/.PZX�`G�HO{,�k_��!4zrp�[=*�h���v8?nn�y�������D�n2�ɍ�.�wQKzgp�sm�L��@
��4�ퟔ���~n��N��R,i�q@��a\��w fA�.�KR�`iв�yܕ���h6��`��[rï,�塉�����p~���G͙9��7k���Iw�Fy'CL�+C�������|�y�g�#S����
4܂�>rL���4�-��ϪS�Z���ۛ�t+���4�|��I�ۨ4��%�\�e���t�OyΣ�K1*�P����v_�lw��9r��TQy�^�}DC_Í��3<��.��䙚d��ڼ�%G����d*`m��A�/��������q�JF� �3¤rC�7�ɦ��[�q��Ҹ�?׽I�n0���������C���y�^S�W)滍��b(�T����u�r�7��U{`%�(FQ�)H`��6��]x��V��b����2�	�,�i�¼������E��ʘ)h\Z����.Vy�֍uϚ��Z���&�,���	���;�=��H5t�ނ��$f�f��\	�{\�]���b\;4������%x�X�2>�7�7�_}%�c5d��g���n��P��ɤ�Ƹa�q�N|�g����X:ԛ�O��C��Ѧ��a�]�՗��z�װ��%V�">2�aY�5o/��vy���y��+�<�  �^�z�o(hd���Y�l;5�	���xn�����Tj�H�99d���{�k@`A�ք6�Â8�2.���!B��U���'�z���5{���ǿ�/t@i��ؠ�n�AZ��ȭ3eV��f"��0�����Vo�߰@�Ų�<�.�k�����hAd��#�j?�( �Rn�VW=){*������P���ܯ�Zѐ�"ܥQ	�Q��z���]AH�D�f�� �?k�Vݍ ���l*6瞴~{[�Wx�Z�%����n�%]��+L0K�����B���y�`���(�_�p
6 ���=���H�����<,�1)�����d��TB�HP�}2	T����2Fm�>��8��քR~]�H�*
�AM�^�7�cu4�qR1&�N�ӷǴߝ�,c,@�q���Y�Ye��Ȁ��>1sQ�i������gL[[��(~m=$7h��@}������d8Fv�c<�Wb�J����
r
������@6&���I(����5��h����-w�:�H���3\}���'%s�c?�������)Zq�|��LUDo(~�S�o<�dai���uǩ2�%4x�'�63�Hf/����LQ_a0�zA7�J��d�@��盓է�kPܐ��n/<SH���9���{�0�B�����kZ�&L��K[�G�Kh��_Q�, ��n����&�^+�Ü��[��+���s��&H����gp��툫gYc%mgGX^��QT���#C�ט��k"��h�L,FC^U�\.'�$m����D���գ�5� u�l$��̂�T"<�.ӹsT�D�JV��	��>�C#��#+i��G��z.B_%#�'��R�;[�	d�����Z`��7ANi{�8D��|ĞA��A"v�#�Cѕ1㇦�ż��'�6#��LU?���\��÷i��^�����ӏ���0��2�CN��#��������̏tO5p�T[��DQ�K�o�}�]�U��lC���4g�U1u�9�Ӂ7XnbU��IKh�ۦ��q����*�&��&��uT'�Z�f�$�����Kk�;/K��M���ɦ��Ϗ�D�#>d1��+ˤ�)���)V
�Z�Pћ��AZ�_C�1Q��NN@*����A��1i��5<�WV�QX~�--������[M�/g]@Q�S��M���(F��g��(�}b]�@�.�|\i<]�TC��s�+!sWgS��ҒLA��9((��(.i�����]ʑ�va�<��[�Z�W3�^�r\�Խ���բ�?l��粔�\��P����/��,F3�O�ƽ���]�C�{�����$؎�p����c�b�(҉5�$��v�����)`�Zku�k�D�'	Z�0���4t֞}���PJ!�D�������5�� �j����v�o�n���L,�F������F��`zcV���Ư���T�v�U����{�r����w��X�4�O����q�җe����5�r�����L���5���q2��d; /�Y0-K�n���]%�#��
D��hJ�Z��ɜ8�w=&���� �ۆ8���wM� �ClhW�*r �%g�)v��jJ�oS�x���{h9#�6���jX�"(c�-��{����%P����3���l�?7�7P�g&���Y }�1q�Ch@���x	D�<k><�Z���%�q��Y	�3s��K=�n8� `27xՁ�����/=�9#z�-�]G�h��_���=�x	��e��{���G_����x뮒��/Zר�&N �ϭ&L�'ӥ��IS��;��.�|F�z���Y�������B��a�?\�K'�y�$����x�ry�5�R�U���OԔ�ȹ���8��vФb�	u�&�]���ù��9�:ez뗣C���P��[��C�! ��Kr	 �w��ܤ���Y�ַO�d>h��i�����\��`�9.Β���Z���Y��zz��_��T��v� ��2zGaX���e�O'5�9d����?k{�%�y�̂bKphc���7�Ӽe� �����⬴��=��Y�w�)�i��BqJX&��\_]Mdz»:��=�c\ij������y�K��"��������9LZqL�T���!�4B7�k��g)��bJ}F�H)k�2�jZ'����R�!���p 2~��~s��Q�Z�[ A���!.���s.�F�i�/��{r�M���$ʊ����aWO���Ɏ�t��x�ʛ ^�x�%�06��,0=�p�B�=����
�:Z2�64�d;�t���~�%�ڑ�d�$�YP0%By�GK�q1�0$� ;�V�i>���6.eQ��S*�v�x�Y��{Pg�ȫR�, �Lp��,�;r2k��Z��r%,�F[�V{��	����N�:Z2|���`��{�u��a��DK��}�lTۉ���N&��\G��3�����Z��!(?gC+)Zkҩ�P�ȗ���+�Tx@���mHUYhMπF
�H! �Ĩ�,{��^��ԋ�N���RL�=��I����7���YoE�,F7�万7	����>�b*d�;��@�0О�[��Ω��W���Y~*LI��H�I�Zvt�|*�[F�QN�{��1L7��4ЅT�qJ��������i�C&��G�$%8$C �����@�C�>�}����/�wu4�0���l9,�%� -߰�>T��;T��nq.��]C���%�*'W���Y�J��30yN^�K���y��3��pvߕR}�WQ��W��S_p�v��#��&5I)����i�/ǄC�y��K��b.� �M\��p�|a2��!�ڼ�Θn���Ί��f{+��͢��ya���"��;��#������8�+������ƞ\ْ�{����F����ٵ�u�$���u]��5�'V?��p��"�[�&)}]J<��{LJŤ"�n���͝�L�xO�æ��!�/f�H9����iS_Q��P�[a��G�~Ŋ���*3p�G\qY����L=�%����F�l�fr=�'@��E�����`e�:�^*��
�dZ���a�2��:���_@�RjQ�gxq)c���&��x���������o.Ͻ$��3o��3�'�6Q.X�K`�:�3ktpF`-�f�W��B�������-ON9�Ш�R ���<�������g(SЕWk� ʞF��&�X�)��U;�}��`p|[?e����tB!��}(��\���T����R�����J�2_�y��f�pO���N��<��3��� ��C�uɒX�o¬U/o0sD���䚀ZV�)y� ֋}0��Sر�vo]�̠��#��.m���֐7*׈�g�;���&�Mz�(����ȯ�涞4G���ԥd32=����Z�t�`w���F|��b�����0���]��"f��<�#e�{xw��Ÿ��:BS�%��?���3�Y@�s�o@��'�|�h#�]���j��<������L�#k�{jO����x��;�n/�aw9���t��W�T�&Ȫq~��,a���E/��NN�d^΢W��q�mqt.��	�����	�XuU�O���3��$��YN��ɀ����S�	�{'���#�,�+���j�"u^pUr�ק�Z%�3�u��l�:�*�Y&-hD�D��;���%8��؏9���ɮ�9��W}^����%#)��XC:ʖ�������g�KX �}&D�C�ڟ}@~"ftVf�L8�������
������K������`<C��K�xD��}rIg��]	���?W5L��a0O��4|����C�n�����f3k%.sz�	"���2H�;��v4��驟H���F.5�+&@�ZjX3�E�u Uu(���3+�ΥZ*���[�ŋ��w��[�+Ä?�5�a����5�?��]S��侣a��Z.G\� ���������%4ؿ��}�>���� �&�6
�!�/��ѣ+|��l���6��6�>޵z�Yw�6��rF���5�R:�X(hj��qU�1��P�}F$�aEP���j���9��1�`��2U�B^\t��Ao#�1���9it��(�Y�wis�c_�K�+׽��k�A�S��� 	[�
}L~���;2(P�}�|��(�YS}Nd���hJ�����#~�%ǹǞ��Lo�ޱ23nU��X
�
p��Wvܗ�KB���$����T5!��(��o돮쎘�h����9�ǝ%=X���G\�&�H#ۜ7��!�M���8��G���9�[�����-��:ϕ����-�!��\��8>�����4�H�y���jGcn:��d�:ؖ���w�>�Հ����n}�Zh��'M�O�I�Ó�q��o!��Ϩ;�k��  �O��~u$�p5RF�R逪��D���q�	�{o?n?8��ɿ���H��I�b����^"�'W8èxgհ �
XKF+G��!�KnH�\?,��ly���J._��Y��%m�5�6:BnL�J;��ǌ`1�ė�AB���
P,�c_9�"�?ϻ��_���k�C��w<��e/Ux����5Oxkld��N�"�����9�(��L����G��B����0E���A|\..#��l2�����ϋj�m4>R��s�a�y?'n������)��C%3�	�*�=��`�N͌��j\*���|�*�SO�����ݐ�C&UD�Ҁ�*�g�0_g�`�-�ٹB�(#W	Q¬���G������ ��	O�a/'��?��4h8K���$�_�N*�&���W��{��$D��M/4�4� 	�*�[Іs{���k��Æ�a�v�J�w)���>�s��Y^	T���~î����VZnƄ��Y&����<���&���Y�R�t�X�o>ޱ�0{4>^wO�Ȕ�����̥��a�ߗ�_��$���n�ԣ��(c�,���Q��la�y!ԢU����4�B��R�f�ݴs�ȧł��ڄ�2m _�Ƭ��9"�"܍�`Ey�
21�(I�M���#y;U����M��Q��Z���s�LBd&=T4P\
�����M�<�[�}�I#�����,FA�B�����k��QQ��[j`PQ�!����V�yk�?F7U�j���q�����a�5$n�t	+w�ƕww�fo1/��\�P����#��覐 ��0���"���t53 ?3�gݱp�<k�"�!}Ĕ�W\IE�n�~ўdЍ��� c����W��5����ې�A�7;Ej�榩LQ�i�F���Ǩa��R�H� $����H������ uD,����yx�y�%߶�/l��a���/��~�7kw�z��#ٿ�u��m=��~�.�Hp.�X��>�ly�}�W��1�	~�����*ʑez��`�!�ĬH)��Xp���5��:��Y��K0jH��h�)��V1��*od�_iU���-��a�m]�LI����P|��	��7�����n��#�D�Ū΋fT�����n�M�&Q�����l踧�t�טE�����H�t1m'�����9-ѦYg��ɬ�-��QI���'�.����!H�A>���-D�_�5O�Mf�X�	�Ix����U�D�W $UG�3��#�����b�$�N��|R����+�,[�i?T� ��{H��`" ����b� pO��/c^�R��n~!����W���3[���I��[gq�KNK:��H|K��ϰ�&*.���^𲍨y%��0(��wj�K �O*�6@۲�l�Q�J?ǈ~�N���$��eA[�K�Z�Qm|Ē�o���;����t��U���Zx��Ӈ$ʱ���(8��\���d���p��W�O� :���Q�qY�r�ׅ������?���t6jXW���͂�C�:����G�3Io���g�MS�QM-��{l)1�����ӵ�되-��Դؒ�JB~�ot"�\�^����R���T��h��,e��+�D~���BR 0���m�����ژD/���Ś�U��RV�Z� o���(U����'*��S��w��3Y4�نnd{7b�p�W��
h����U��&
I8���3�}f��7E?V���c/[,t]eHC�ψ��f�80P=w�_�m���l4�w8���������9�8=��_��*��Aw����χ��ی����G���������PK*
T�6�����.w2s�p�h�L����?~��Ҟr�S�wB��@�y�v�=2ת���{s
蹍�f= m�u��JI���`��[Z�h��end %��*�+�k���\cI�՗]����G������X�`�i~G��O�� \���n��l��3�1)�y�w�Օ��`��\�<��pP���Zj�s�Pv�^�o�#�ȧ��q�Ʊ2�K�j��`2�E=H�χ��k��nb�{}`�S�30.
�gwC� SO:)�ҧv����l�&��$,��$0�J�q@0�	����[�o"PO��E��)l�k舉��a.?���k�'�#e�UC�\��8*�̪�*
[�th��{�/йױ���)8�gYy�j��J� QB�..�rc_�dZ�-�ou�q����u�o:�r�[M$pϥjU����p[��VCqc���2�C�
����0J��3�������@�qР��T���"g�O�k{!7g���t^�㩂�g��%	S�P蹵9`�^�^�1A�M6�V�=*��TX��y��ڹ��gw���������̍o�Ħh�T] D&g�v�B��FlqW���V}���������2~P���� ��c��̄U4�sG���U����,�BX~����~V��Cϋ�ʌ������Ċ�u�j5�Ϲ!��Bw��5���9���̬��}9�ǡ̆3��������7�s���*o��i�X����!�η�aw� ��$�B�$�(�8��a� r鷑A�W�\*�-�5	�Y������ᐲ���y���wKn��k���z��I�~��m�n�-#�~�&��@%���w��;�,M#+��P�G��RV�4r��v�9X�N����M�1��+��k�J�K�eY8��<mIB�&�� J�Uݪ�PЗa�:e7��s��atz�@<pO��Y�t��	W>O�5���^0�ŞY�\�t�7u9���3�-p�V���	��	{W/�>-�p�3���]�"�[PD��1�_���W���.T񾼮���-m��~�!����P
��I���j�V�9#���,�s���¹�_?�=���U�N���ʊ�L��3��F�x���"|�?���Y�����,d98����VR:	G�c��=J�t��!�&��ZA%۔���qߧw�_��V*�v���$χ��!��gSr�ph)�>9�����X
|6ܧ����Q�}�r1�b���r�>�����3���)3V	��2��"_K#���ĭ&�i�����Թ���LOF���@7i���fr L�zc�đI<��pL�|��ƈ��H�0Bb1>A������
hC��>�w��ST?H䲷�ڻ�p�z��E��˗���l\#;�j)��*	'�4w4V�u���g���<��l�=D��4<m��v0X��m,%E�)g�
D�|���~Z5�g6/6�T�և��hG����
���~�:(��}�&Ne"/�����0��4[�̅�e�%ܙH�M\Z���ߟ̥��`B7�m,ޛ �r�K�_��F���s*,䩫FD�o�L�n9��
�,'cH�Ϯ�$�4�-.��w��ǋ
5��@���:�ʶ,YO�����dGK���|׺Q0r�UÐPuC�Ǟ��~S?�e�=�`���� rʅ��%�����3��s�i���vg����B����O<`��ö�>��#	��z/W��a!(�N!K}�$!���j%3�g��*�F��U��M_��
��?w���0��<��ux�ָ��s��^��W6�C����6���ޘ�&���ź����[Kh�5�ny��}ۼ%O�S�����[�>n!��5�C�>��D[�FA��O��ԘB��9'8@�C����au�P\-�Y���*��<y���3'��=�g4����������Q�«�_H���!��S���)dd=W7�ܞ<MԬ�C12�TT���:~��Lc�Dj�­�p~�u�S�^�sVL���*t��צ���D�U6�nK�{*��i�u}	��v4p>N�/jV�`���:�� �O�D���j
�)��'���<NY�D;�5j�rb<���z\�-�^�_�1@�z�'�ΝB����z�rWl�o��y������Vb8H����m%U�݂5�y��$+XRz �o]/T_�p[ӥ+��i!۳�k��x�:	_��6�����=b���˒>����B~��J�6xkƞa״��	'T<�Q�FJ8��~�7U#��x�P,�*_w�t5����H�D���������\���������؉��<��Ɵ�'�)��b=��v���"�7$+�c�_�0��������oS�s��J��;A�f�n�a���<��L-4�.q�����1ƨxI��݄7i� .�0�nm�Ա�'4�g�Ax�O��H��Q/2��F�',�y�L����Z5��-��ѵs��={F�-�jC�e�2'�R!��*�b��*����(��$�27�i4�::yN2�o17h���W�,a�[��QS{|�]Z�E��s,�V��\7�0�Ps���dcҦ���Z.����d-��Ԭ�:�3(`��	��6Q�벿"Q߿Ї�wߵB�
e���N~Ώh.�ʹ�韃r���
��Yq��| Q�E�Ae��ݎ\��g3�yp���4{]��uc���ݼ�#�^����+�%�X��*�(9�$�hy�N79Q<6αz~���M7������ً�Ew@��tRen&��#��ֺ	���['R�3 ������O��S�:%�:��Q�ƾYsGn:x�y�D��sGnS�q��ZVu��F3/�Nڴ��Ze�h�1�>]L����P/<�gŦ2��dñZ:���H
���"]�Y�un��Vo���	U
��x ������ �;X�����*��ϔ�s��K���튱���΀�x�s��iO;�����qoY)I;�j\F��T�R�9bޯE����U*\��ÄC#P���Y�5�+Jn=��a����s	��n������z@;=�^D�e�%&��
���ǖ�C^��~H��u�۬�jy�X���JWO��|��bl3!��y>7�$ԙc�W�ix��I�]��0F�fPp���o��ۋ�lh���^/=A��v����K%F��U����+����108�/D�'ſ��M1!p��&��8�P��?:&��m΍��!̴��׾~kg`�=��)�p�0��M��FR��r!f���w�&�/��k?׮���w��#�=q��do�?U���б�
����y�z��#g�����9)�~.��B���%c��n��*�"�~Z���ac�YyD�_�	��PU@��@�8�J�Ɵ{b�UQ���v\�A>��������AT�RwvY\^Gp4(������.�W�SE kj�+�Œ�F��"���-�w�n�Y#_1>P�C���A����O��!7���z��	Xi@��JN�O���'Tr�`�*�u�P[j�Jk��w��$4e	�V!7mzkbpt^���;\|PX��U�fX|0�u֙���M�e�d1UU� �f,�cɲx 3���n��1u\�����cŽ�vԏ�:�'���Y�^.�=Am�iI�_v��@� ڞ^�V��V���l��/��������w��O��BH挋i�h���|]�&�Mt� 9Uv�)N�#��G�";�K���R��$�T�i�q�����K�0���<=�~_G�]ɣ��D�kv���4R��㷋����������`(�{cR�׀Fd��ۚ���}	|�{E�plǠ�&���i�:ތQS6?����3�+9�Oj�ܿm�����E+M<�A��JG�pu6��@N��蘤�.���������τ4�6��"���+v��S����R�u��Ax�c1q���XĚ\�OE�롖��_J�2p�#��~���Ly2��(�q��8�إ�>�b��OʕC��(�c�Ғ�̚k!���gk���ur�M#�t�l���I�����/=]�7{Ȓ��Mqao�����s�q3D�˂	#�K?�4|����mMމL�(r7�L����������z�4�1��BJ��C�g"��[�_��rAQ3�j�d��o�[�I	9��]r��i�D:��K�-w����֠Xޫ�6L��Ql��:��R�c§J\�a��ΑT�p�f��A$�:���2czZ���r�rL���uR��Ҙd?�R�XÆ7��x�B
/y��;��>�ڢ�g��h�8��5t�0�E��kYyOD�[vX��h{��Dao�<��.��z~G�P�Bv�2_^�6���M��c�(�b/��Y�$�ft���bg@'"�| �^g����w�E��e�����A]�2����(���ѡ\M2�R_���7u76��-v3Z��`
�H�U��&�~ٵjҷQ�`���$�z���0-𗞽/F���븣�@KSMGc�I����
s�O�x$,���b4RBX���޾������M
Cl�r��_�2mq&�,����J�4(��o��CcR'��q�`��M��3�4F���5-4d�-��9B�\��jcA�?A�U}��3��p�L�7Eb,��0�~����zc��zۂWa>ȷ:IH��I��Hό��7 �V�Y��'l�R;�=m
��~鶨h�w��ڧ�͆�� �L\��5�C'@c����r�>�����v��ln�Gr폗���c�/�\����N/�V����YR����c���&�O0[�@�aq�;�4W�]8�#l��{)J�$�W-����2���P�Z뢤#'���ǚ�hxrHd>i���U:b�߲��ne/�5~#��:(�<�[Y��%�&����J�1�����w6|��pc
�6w���2k]���C!Q�;��־�x���@�~�K rk��:? z����,��Qgt��g5�H��^��o�Fh-G�F�Z"�^\���i�4(����u�?RF�5��X En�v���Q�4�g��*�����A��Di���rOP��8§�8��4�g�$�ܺ���Aw�q�����e��B�ƶ���W�Q��ϼ+���{�>�(�o�ۼE@�GJq�8x~��?m܏R���q���I��p/  ����G������Ppf/�{�/����@�v������ʰ_�v��ܯ"nۭ�pc�n�t���u�7�͆R
�i'��%s�S���d\TKz~��\�=4���������+N��'"#u�!�N�4��%K�h��}4��%A���Og>F����~���A|b1�v-A��{؛��w����;�w�89X�ҁm�:6�j�k2�6�Η�{�l��0Vp�"U�^7�1�#fLM��z���?� h�!����֑}�
2J�!�/���Ϟ5\�RCI$f7��#N�%��C�š0�=�m���C�
(X���~��j'����q�{cn�}�{��[z���?�Hc��vr�+���,B	�T�T_����*c�q���#h����X��i3��9:�ɇ��OW8�C���qd����%X=�q�3 i�S�����I�-����a�&��a ��r���^
R����iJ�D���Ps	��@a%{pP�a�> t��ݒ�+�'L�֋sY%m_?5��	������s��2f<����@�c�]��/�� F���n�.�K�f�n���Dul���a�8) ���!��?8��`,�ܓ�����I\\���6ڮ�~�e}��/�FGTGk0�$���og��<Q����?f��H�6��k��[��4`���?��ė��Hʔ=3P5�-?����=����qBe#h^�oi"&c<���,[{�}-��!n���R�
��Ƌ� �M�Ѧ����V]��;�,o�EC��nGm6��TI�Dj���d���Hr��O��T����-�aD;��?fcnB#�� �ۊ�@;��z� �X�4�	�'��\'\^�P�\7�~�H��L�j��S&�t��M����2u���H�M�<r�2��L�����u+{��D�;7��V3��Q��\�q�Ȋ�-r�@�}L�-�;�#^�j(�!>��
���<,��gU�aM���X�C^����y���)�D�����PV�5����1��'�M(��@�� Y(��3�\���H��ӄ�B��%FI��8f�a�����{� ������.}�����=c�(*%ס�	n��UJ���9�	�ݬh�h^?f������`���A���M�g5���i�ٲC��Ӗl0VI�U8�.$59*��'������Kl�mF���>�~�MR��@�����Z9�[����Q�=~�:~�HK1���=Q4PK4�'}�0���tE�,�Yë�2��Hp�J����#	�e�Fٷr.fϭL�����N�|�P�Χ�T#��h�I,��W��3�5��"�xj�96�����g�k6��2�H�F�!oߤ�m�Ϥ���}���~җ/��p'�*���m,�a��ݣ��c��|�r\��#��f�.�W@�L�����ĺ����QP���G�[�%�����>�%� 0Y�9���[��mL���R1I�_�f��[<(��(%����C�xW`E����f���#��(��/5����ӻ&ċ��PQ����هa�YF��<�ܚK��4���-��V*>s���j�5������V�b�{��*t*�����ľ,=
�	�,�r�}���x���DI1��<!�x�'�qI���ba-A{�CVt��v�d����'��"�}N	�G�r8S34���7��
�цI��3��΍�c�;�35�	{ �����1V-������5� ��~������Q��L
�ƫ+z���6VDY+Z�q����v��s���M(ʐpw��f�v��_�7U�{B7���ڃ�����;49���mp�:��j;�K��Gg�g��X���J���z8���>�U�n'��c�z��	n�{y��L2��|�tx�McQ�&۲I�V�<�@�}�0�Sp�WxX9$������x��&q�;���T���!B1�-�[4"���5<=_�Y�*�d`��qm�s��=���b�Fe?���o�ߴ̛v��8��{�3����^f�dx��7�dx{�駵S��ɕ}�V�)�o��wOx�R���ĭ>�J���x��Q�ӄ`�lEuX���t�C��jڟB���Ԏ��wn�ǝ��M��5|��c{���4�������Nh]b'@

�`���Z�*�@�j���٢u�lU�ҋ�&�*���X��.u�lx��Fp$e��&�W\ieG�43�Jw`c,a��}���[Y��+�z�~��Zo5U$P$B����q�Ʌ�<= Ry�Ԥ^�u �������vCm������[�������䶋k
�� =���渞xA��	�5}輒�;-��	��6�6n�e<񌪒�����?��-��wCѼj��x�7�S�jM�M��	a�էG�e�2�\�����%n���[J�g��E�8��p�#�OX(� �k=�	�g�C��6"�9flR&b�pc��3:���Lm2�0q2-��#�*��JŀP	�+������#B3ƨ��-�'�k=7q�TIcW��B��q�kĔ\I'S��Z��*��K��j�����6�lȕh��PzvQ��78��f}���Y��?b�y=�4~#h�p��ۨIl�:2H�+e -4F8o�E��{�����a�N�ԣzL�q����R@[чc���!cp�Y���88}im7�6�:����R:f��#����������ִI����6�1.��������׷(=_a)/J	>\���.��US��dV(�M��Hs���h�f��* ooF{��Ev�з���s&z����$�g�4�C'#�0��I�k�OR��BEb/��c���۔NEj��ҊZg��J	�A��X�G��OF\���pz���ι�<�jGs;.��}�!������SK�<%Nq\�u���~0�gٚ��r9���G�ٌ*)���ѪĜ�D�t,fؒp��ls��p2�!�ܤ��hЇ�>�����GZ�`�~�w�O�c^x��lڣUK�̨��k�D��`5�( �- �+��V��(8�_�*��LC�&�0�jw��9-����vN��)e1�� �1��)�'#�����6���{	�ɑ�}i�d�d�ĺ˔����\�ᆰo�V��w[.���㥨��>�F���b�p�(���>/�T�x�� ?o��qYP�_T��� Ow���l��'ΨڳX�� O�g����}�Bs%�fG�c�t"M���c�\�x�27�TY�y�`��:��z�Ȁ�?b�D$�{��a_u�j�>���I�X�����.�����ݎRO�����	BU7���~Q_�����rk�PI���(�"o���'�J[��C�w�go����3��j�  ��ꐃl�<?����k#h!FV�|�o�"�e��?�vs`�-�*>!�������j�����Qc�i~�o�5����S�� ~��>����7��x���匑G~�,<�H�;�͔��N��U�X ���;F]�0�V�jV���>�����C|Y�x��KvX�p)
h���D�~M�����+cdԮ}O<�G1tTG�Lo&���*�-y^o=����7&{X��0� �~-u�XM��QS����	ԏ;J;l� �}f��x����+m�r�Ηr��Y���b\���#lb�5��p���"���*I����C ��K��`zR��xap�C�g1�]�B@�?�I�v9����'

��ڬ���$�֫rِ��qJ�!jp�xD]��uW8���E��t�F<�N�w0P���f��Y3�ݶ �Q�\>�����|_��nk����q�"uSVy�' ���w>���D�_��b��!�Uox����b� ,��~�G[�K8}�UD=�&7�\'1a�0�0���쌄�'}�&���n+'�0O"%g��F�8��Hw�?\Å׼��G�N=���씰�;-��BO�O�q���6��C�3�`d̩Y�L*�(V���LRTM׿�Y�[��qeq�z�&���n>��%���F�R]�����Mz��~[��=f��%'W4��-��2��}2��� ��_o[��m+�3ō"�^��+~p��]�+Ph�v�U/��՟���>+�eO�u2R�C� 0XK�CW��/j6
���U�Kx�@�s�Ղ���{m�T����y��"��і"RÍ�`�k�h�;[iq�����o��j����pl��iA���(;���t��K�o/�@S��[��+N1/'Z�9MQ}���m}�rk2�s ���׍4%~�M�fi�l��<B��A�DCA�K���L6�M�#H�r[�6oN�%���h>�����l��9x3�o�@��Lxz��W��\e@����D�5ə��}9ܔv�l��$-N�|�yPd��"�f>��&�	7�?B�D!ah���q�-8�tA0!��E�3���V�?��a�9����8="=���B2����q�q��n{��Qg���[�
�f:�Z\p?�eVX�)��(���	`�&��=}re/As�ޛ�gOzK,�9X�F��y�oq�5�6'.N�Oq�O��fq��o�\�����И���%��#�ߵ��Vu���n��N��?ǌS��U�>PZ�I(�{�0��ҕ��D�W�!q�&Ը�<��tع�zc��9�nxM��H�Y�{��&M�ε0�����e V�rAy����2��dyo�����u�_5:�M�Ԋ!��E"���
��jKVk�]^�e3�Mki@k}�F�5�=�L�v)9͎�v�*��,���lŰ5��3�o��������Y`+��H"����vrH��|��y��7��2}���k����*�~�^3��[��<Ƽ��581���F��k8M4��m�A����vS=+sg���;��ٰ�p��U�? ~�*�Ɓ	]�-g��Ki��w���� �_O7�d ����<L��-[�؆~ޕ�^*w튆V���",)2�DM?���R^7�ǞғqW�f�c�9������PzLqS�9��G0��������G�J�f��~�R�)�,�0^�F|=��Em����� k[t� �T�h�#'Lq�l�Z.�Ud2���-�O���[4�������|KU=S>7E�BZ��W9,��;Z�	�;%JC|I�LY�G.ↄW�`�E�#9�,N`z��)$�6�P��Y���/\��������٪\�[m�d&;���[�q���z�f�$�3��ψ)�~ΥAe�N�h��>����4/�߰��E��@����HB�wz�Q��G�M+�(�0k����>1co�@#n�@C�򼷦Dd������܀Ǔ�Y�5JLH�N�6d�7IA.�K4t�s�k=���)/��h��@?�O��է�z@�j �+�<�c��Ԓ����+!L��������t�o#���� G||�PZG�2�5'UUT���c�˅��0kw��Ey]+�6��	��[��%���3��}_$��m�Epi�kߝ�c�5�Rє����q��8���gt3&M?�����|���Z3�Ap���nb؋�N>�$��d|��H<ػ�o7���#�;&>�͝$��_YN�^	�_���ԙ�W���i�61eMZO��X�M ��U�tl�9®��k��M8-���	-�Z��S�-x���xv����wND#�#N�_�o�d1#�Pi��P�� Q���������ݞc�;�4܅ߝP��ڭ�+�s�C���������8��f�B�'�9><�	���~@�q�$"��(�T��m )���a��8k�IJ��U:�ĂDj:C$4nh�!RE.���kPu_�+s�Y����R��њf��}Xc�wV������OJ���2I�G�~�[`V'9�Ä� �����֌(Uʌg����TҖz��R��THo�?;��F���$�)k�4�]p)�xJ��9��Gy��go4�y�
wDz�q.m~tw�����&[��:����V�Iy:�e����'�%(�f�/t��bX4������"�5ͷQ�Py�\U��~SM���ָHp6S=U��Ѵ��F��MN�=~%� ű�}��.�߻j��� ww��V?':��:��,��k^��𥉉}���W=8��XN �tΕf!��tB��`m�dhu�O-��~�4[���/�5��)�Be�ޝG�l��?���$kz��)q����&�\D��<)�����I�B\���@s�O�l�w^)��'`(�n����L<m?U�G����*Q�s�,� ݜ�,7,b�^��ж�� ��AWc�X���>?0ڢ
'�5���x��
L�I�l��[��J��	�s4�w6��"�1G��~���b�W��Jb4J�� �U4��W#��9��12��H3z'�}G�1��?��HS��,3Y�M���i)V�
��."�TG���p��N� �y���S^���![%����Y�~JU֫;�rBG4�	g���S���j�լ1ѭx�H���W}>����V��"��xu������Ur�9t��Y�@�Xy_O�N�_�&
�}�p�)��M��I�d�Y����̴���1$=�HSD���%ȇ�M�J�D�(Y�ު��s�o�L'�g�p_%�V�xJDx���)��K�c&n_*���v��17]�7��q�1$qf�8EAM��iR����'�qe�?�6S���6�HOc���y��M�kR����9�^I�x�� �Wy������a|�e�(�A��8����%���P�|�w�NJ˼X�5}�zu�G���q�lh�%E��"�S� ��©I��ZcٝHv���|�V��A��/(O'A���*��>�c�����G(S���C�ۮW ճ�����
��C>�d/�{M����T�\}��Iv�(;Ez�}~Nav�5�$?Ͻ�	��S����p�S���ٷ+w�m��\��rgJB�ݟ_��f��)��s!3���وV>9�
ު.M����%�����"3�[mj�c��?3�ʊ�U�:�t��=�w-����o�~ ��N7]F۾��n=�Y&�yJ_�c{}|���B�{&w]T1���N�z�ց���\���V�@�Pϡ`v��^)�������`�N�C�b2�}h~�G���"��yJ�w�����p���y�/�i;X�%���M�w���ޢ�,ı�k����2������G8.A<��{�u^=]*��Ч��h0P۱0��\%Pϥ,o�f��j�ī%?t�hs�s����Ǻ�6�r6�e�����o�e>��p!뗪�93����<x�9g�#�C	7��s&�'����C=���ra2�SQ�[�4��FgoE=n����h3����R�
���h� 1}�$V(���Ǯ3�
7l��2�Yqy�0���'^�t�����ZX��;̎��>K&G�Z�����**��b�\��B�ã~���{,b�]��Q�R^�٢�+l��V�q�4KN2�%��H��i���fQv��2S�'� R�C�a��.*�<}�Քi/�D�[�l;�`G8�i�ejz-�g�x����i�z5�+��:�o�@�Չ`V2�
�0����C/ο �oG.a�5�"��1>� /-��{�\���T��L��h�i��&�*��v��ဗ�]j�+�Lc�"%R����e��!U�sQLE�aQ+�$�1����@��A���酨��a�
�R���|�Fu�k�P��܏t?9w������df��v�K���߮jw���,���7�|6�5�+Ip���П���*I������� �ͫ���-��K���4Z����k�4K�D�y�P���j�~9�<�%����Q�ԫ�UFH�����+��4���;�z��Z���"���kh'}�� �u�L����Ge�d'�@�={�h{���D���q{M|ע�D^@�U��%E*�R<!��$����#O���6
y���R�6
�q����*9�z|-_L>�%�%�&A%D�=�:ي.��͠�.��ڥ]�KI;�5|�NQӁ�k������0~�ؖ�u �͂
��>��4|O@��k��V���x݅�z�:i���f5���=�%Yn\���fڄ�"䃘R�:d?���jTac��aV�T��{�|A�//�R
N� ���F�/ٹD��|��&�̶r����!Һ�S
���6.�lZuaZ7�ZFW��g"�M�:������������`��R�ǩo}�����pw!�u�fL�p�ږXbX�6���W�����:~hT3�ʹ�A$Óϑ�A1#M�n��9G�0s�M�F�b���������$���?�"�3�or7��D�x��d�F�Њ�BN��N_+�:4����C�*�f�e����1)�`� ��wj6׺�2�d��z��C��;N�WƵ�9�~?���{�Y&���O�l2�(Ks��
�Pp�L� �����y5�*T� �`���� �$�{A�6�7���Ns@�3U�`v[�ݕ�ߐDrmVh���v9�\ۗ��;����B�`�\��ZE}��vO���4g�1i8�|���?��,,7�< �n���Ŧ�z�߸��g`o|xy�gx�k+(���+�;��hb~|��UPZ�K�Fs�(L�*�}��"S1�W#�:1��@
q�8��V��`<|����w�l�<0�*�����&X&*�~9A7��L�O��]#�A�~: #���������*2@!6��M>�����MO;	�7�k'�1�0Ģ?���%<�n!���������n�H3s>+ku����#��x+	�@��-�ɼ�&��{�b���r\�Vw��4��tDCD��<;��� k�Wq��臀�k~
�@ �hE^>.'R=�:�Kw�<α�g�r�m�|ɇ�-����7��;%�.$r��f��Y��b��T���|��!�"A5Ȱ1�mn�zJ�Y�+�K�?Ŕ�����+���bdF�����n�n��RI߱Jw��;����uS��W�4������I`@�nZ*��e���
�6
�$8(�3���s����s�&�!^e�tZeF	{����Xk�Ϥ��c�b.n�
 ��ZUO2T{a$��tJ;8|��fk�# 1�L���8}G�U���]ӹO�<�[}i��5�P�å�TYf�������g�'I�㕱k�5AŜ՗cW`%�L����O�.Lm����@wg����M*H�\��֎ݚ?��\X�"@��W�44�"��ɯ��ڈ,m�� <�w�:�p���]�VC�$��er$!�I����
k����g�Ɲ^��+�7���n8rg"{:�J����Ťx�#�L��}J��td�%X滲��x��r�|/���я	�8[ABE;l�YC��4zJ��pUy-9�E��LR��ԕ�Ǧ7�9bv�$x19��]Rq�?�ʾҿ����^T�#+��q�3}'��ch��`ɬEn�&X�{������E�h�ow�)u^�s:�m��۷;G��-�#���v�u�GI���s:E(�Q_�=���j'5R��� gCimT*zTV�����i�11]��F���?m�a�Bl�֎��AO���������%�H�&
y�s�"�r�3抟<�0qΖg�
��U��������]6��X}����ͫ��J1��Q ;�b.�XC�٨:�� *r�5ga�hݯB����0b���y�JW�����뻨+���2tOģ0��
�(.0��t��N�!�х��Y� ���r&	����+�FjmP���w��<�aD��gr�����]i��W�n��D'y��B�f3ۆ4C�7�^�E��M}39�s�
��"=N/@�h,Ȧ�t���T��̮�x�+.zo@����k�������ͅ���)�ο&(e�U�k��:oh����WRO>^g$| i�YCa�}��>���[H[Q$�lS0��m�^{��^L]����
�J�'��G��d����	a9�J���xi ����P 1�ƪ/r3 �	��/�64	O>%���9���$�����Tm��EVA @�N���IM�y/�tpnI�m�ط4.�|�������+�r��@w���8�֝n�\�`�w��t�4ZOm!����Kc�z��y_0����%�챀�L�?Gd*��Q0f�\y�oɷ��bN�z�h�޷w�_�z���{�Y^��E��Vr���<�'��x�̄64�%˨}_E��|�~�?�y:*�ymc��To�Z�V��T8� e�/�ۜӨ��\t�q2�����s:
�L��e�3`r��!<��ے��,i�o�'������N�OvDEF�$��ڰL�s�����#n�`O�=�����Ѝ�P�a�:��{��V�Vr��`���a��6yp�Z�Y�\�lΌ�p��A�~��	��g�'��(q�[��@���D4{��~i8\.�����3��
��k7��c2�*$�,�֍�><H��p�uh�v<q��8�,���{�lP�~s��%����Wj�hd=r6'>�O;x�B�?|s���ƪ�;kg���˕'�c9=F�ևu�_�#;��P#��6w~[���0��*^/�[|�G����t�z�'�b�T�q3.+�u�6C�%Fslh����T�M#f@r�����Tw����!�" �l�^.@|˯7���x|R�|�Tv/B�V��[�Ϟ�V9��U��5��+w�d�b�<K��|�<�H��Zx$}�#V����țj�7'&{e��,X�T>��%Ӱ\�����Fk�bś��k櫕V�uQ����&��l���,,����S?6�a'�Cp"��k�C�]*��K<<��MgT�9<�Xr_�f��_�
�x	=��]3P>;Ve@{YHr����O�>f__z�i�Peh��S@�0Z�W,2�����K�tmm�.�ئ1��HL|� �k��4�W�'�]�
�A�T[W�ؐ�|/�/t�SF0��Ux�~ږ4
V��Ͻ�����Kkx���iH��&kS����<0�p��)Q:,��9̈lu�Rd�%����A�[w�ݻ�};R�|v&��8"����R��G.6�c�	ct��t�}�o�\�h����4uzQwg�#��w�昨\
��U�2�_���W��g�epy��t�I�J�K1
�_ �3b
����ǂ�`�wmFtZa������{W�������g'c/��*v����OfF���!�]��saS��o����t4|�� Pof.0�����B�< �]�'�Ae8�V�r�g���Ѥ��*cб
�.~c��5R�g�^b�~�\^ǡ��>�4ϖ�s��dJ�Sxv�����կ8�͡��BҊ�E�]lJzN��#�\�K�MJ���H�mB~��J{������EN����(x�vG-N�w٫YWXb���@��}�
�I#��wgS��Heņ˻��&�UP���f��XJ�Ş�GF:�(�ɀH\޲�Y��)�E���b[-i����Y��|�p�S�P��sι��i�7�7ٹک�u,�#�`HLq%M��#Jeu�*fH|���	ly���fy��D�rP�o`uCQo�����L`R;��g��au������N0Y0��đ���,�n�'
��"?�a|FOt@���`fs9ٴo(�O� f��z�� ���}�z��xnQ��Q�9wK��4?S�C�/�z������
9۳K>�,��\�χ�(i+������xC�ïR1����~sؚ���A�e#2�PuN���y���@�\�щ3Xhz.[�
;����%K�|։>Cau��p-�I���b�x�j*K�tFF��9ߘ�4	�Vs��pP�P~��7����Дbl=o�(�B��:B�:�
��L�p#��;M�>B��Z�V�Gs������XjsL�'�&	���fF`�����+�1�� H��6@��ލ������ݯKo��+&�}z�6L�\v�X�Gy��Ugy@��'̲ d'��Jq��YK,�X�M��Ƹ������:O��t�6A��4WH��_����-2e�}&;�����{�(�.[�ce;��5|�� �_d�X��5Pap��Q�+��os�6C"zK%1.���#O��yZ70�2���`���&W��߾�H�_0� �սu�VEi�gW�(d���
_AHG�L��υ��0/������0̊vw��af-�u��c)��؏����-��h�N����v���SBՆ.e Ǉ࣑�J�����K��L�W��	���kڧ��S�~z:�L���q~��f���ck�nmㆇ�(О�&>��^+��R|Fn�ÐK�s�a\�����(��#�blZ��j�	�
ozNg��^'��>3���ʳ��YU&���� �S���Մ(	��Y�J�P�����Kd����J��7Y� �j�CH�[#�~Ďݼ�xTW}��;���^\���n��A".D��v.��H����ī��!��b�ǅ���`� �Rۑ�\�󈱀�L?.�����E�,QZn�3���EA��n����m��U�|�Z��O�D'�@}�fx�.�&oX3l H��K��h1��$>�FNo��H����d�0CR����"�)�qf�����I�Sy�1=�D�ө8{�����������'t�iN�h�v ����r�1n���Y1.fT��r��vTp������31�zv=5��Eo>*�4�ڎ;,M%ʃ�	���vO��E����jO;=zLf�a)�J����v Í�W/sU�=�7���э�5���-+��$[Wk���,��$/w6���uB�m�T��;c,�G�����\��D��:wu��d�7M��Q#� W��R��ʫ���d���V+�(˅g��CA똎���	�ه��?؀
�}
��Q$�)���i6��d�։\�G��3�`�����J�zK���7��
^D��:�����l� ���A[b��+�3�.}_eȗ��Y'ͪ�JԨ��P�����	��+��@v�?uS��R�O�@W��0T�/C�TB��pƾ0˫��Ȏ��ui�9^
���/1�\E�~H�_3��	��-�*���<�V�sT���Z)����|'��ӹ����&��jC�|�]Ҋ��l+0��5���UQL7�����B�7�O�t����&/�I�+��:�2���{hA���EM��/NY�'��<+���a��W*�R��#���NP���!E��7��F	o�Aim��k� �� .`w�_y@(J<�U��п3\���cV�ꋭ�Fɕ3�i�1^���E�㪮M��R�uDM��I`�����u���#�������� e!�HQ[��sޢ��X�N��\��K@�1��y��O�x�<(��[��}�N�1ʀCgJ)I!�9�ΖsH:�2+�^�wU�0��߯KC���`�HB��&�A�|;���	A� *��=�{آ��<����hG-�l����o�{t4��5T��3�}�
w�7"I��R<'������a�~+��兼A�$Ǹ�# �p¡�B�[.i��=Qn���Ϲ��{G�����M˥u�_s�4���e^�#
$I Bw4�e�J�d�l��Zk�裨�F�jg��p�!`%���r_=�oo
�l#���b�WJ	*Hݞ�|���!�S�tyA�E�~U`� �"�Y$��YlH��`L@!\ĸ&�ϖ�^fI������c�-~��Ө�4XA9g����'�(�4c�\`h\D�r緐D��\Ж�#���b��G\,y�.%��%MݲX��=���$e��O�V�W���[ބp�=e%�)���U$6�(�a?K�4ُ]�!�+�7Kl�'ԏ,��@4:�O�(H����PlBt �h�%�s�ދ�p��9�ӭ��+z�Y�<νc�L��D�L\2W�X��pSڞaȉtj�^�M�B��G�U���߃UPQ�K���E��MR��`���3i��|��w�*�޼��e�uL�3��'}�bJ�&�-J��uB^U����mD9�ΘJ�Xn�d253�
���ٱ?y�}��ߨk%uuEG7���iH��4L�|�h3[X8.ŧ~��ቨH�&��6M+�)��5(�uUl��Q��A��S!�Py���Ա]Qգ�W��:�E�vL�T��[�֢�PD�H�-��/�m8F@�4�S�l7��d���I�/���}�x�B�M����N~L�g���+���i�53�
YI*}K�Cd��sq�Wr>?����%�:��-��x�%X�4�T|�>īC���I��Og����.y�Ĥ��.�ŏo�|;������֋�޴[g{�}�z���[G�0l&0���.(���ϛ�Z�����Jz���!�A9^�|�z�[��-�K
.�H�!��6��<W��^���>���$�הjҮ7:�������B88�Ų��q�O���~=h 85\ɪL�ju\�}zř`��5H���Z �l8�I���4P��DS�̢3���:i�;���6�	�Fzr�e��g�M2��I#�Cu�@VGO�B�6�縑s���i���Ѽ�1iv�/c�ߏ���n��sg�Ԫ�2s1��6W�i������_^�]/F���[D���1���$�7l�R\�F��<�t8��N�rݾ�L�h�΋o}_O�J�0��u��CR;[`���aO��b��O�Ë��恃U�T���U	b�1u�ιJ�=]ȣ��8���E��s"��]f��$%`�����~�X��%p��XBpJR&k`�
���q+�F_y�ۊuW�ᥔ���}v����U�T��9�����Hե�6���sL~Ȭ$P.ָQ�/o����&8��'G��@6p?.c�$��]��lf`}��B7h+W��004Y!�J�+��j �ǈ�Xl�E �F�ڻ)�lW>J�}b>���=M�}����B����K���6}��nݓq��[Cj�vŀf���|#�ahd��Q�Ϥ��##�8���%�=���#��K_���m}�M:�P���kO�(pn�¼�K���K���r(�ڄM1˯J��`����X��V���Ib����7l*h2��)]���U���őw���W���o���"��0��%lR5��{� ��J�~ᕓ�W�o�gso+��F�� Pb�Z0t�!Yn�������2Hg���H 	�
'�{���ky��l<TK�;�B��tn�|~n��h�� �T�r�D���;��ʓ�W׻^] �*?U�n�9���4Ƕ�.��!ɃЎ��W?>�y�:%��K�hilI�A���b�������j��:SҜ�=���RL��N���7N��g3�����0�NO�C�����N[�>��֥s�DK��΀ ������l�@��ҡP�R9�����O���K��f\�n�)�Ӂ���?�ç��`���%8��,�NFt�ˋ��~eN�1��E�ވ�ǜ�)��0S�J��$�鵞��8����gjaNѽ�ƶP�E.a�!�uY2YAؓ>c�	(���jX���l�a��B6Ԍ���I�+��z�(��?�>�ڠ�w}���՟��ŇXh�u(s��,�a�2��{�S9�Hi2�(�_�̤ب��,�Oz���z�+.��l/L
�S�U���<#6W�>C7,��Bc8Q�ok�\g��
����U:� 񉠑� ��45?xa�b�Q֜���Q��~�Uo��D|y�lJ(p������I(��]⃊��O����ЂEA[�d��=L�ۇ���nZ�3�	x��/o��d����hC���%?�:L��s�z�r��kN�$�!+�����?�xm7������B\	����!2=JH#K�ǅ�}ۈ��r(O�u�O#���)�K�A�]�~��"�T?��1 M�k�+�ZbWI&�
�ɥ��D�E���'L3w����������b��p(X{ٗM�������T�I���i�<�8q��Ό�o$�o��)�,�1��aǤZ�t};�3O��ίTB�b�+i����xX�c:�P�a�Sں7�?��EN����/��yS�ѭ���7��c�@M���<��GEOЁ��=��k0�+_�(���GV�t����D�f����Y�E$RE1�������@�i���H�~R/}�=�i��m�ꌂm��IJ��"7��`�k���.M3�h��W��J.z؞~�#NAb������3S1����0C�4�.���q�P�?�'68v��'���ټ����qP�z ɺ#*���F�t�#�x{�[�ff�Q�p�s�~+�;�Q���z�T��v>��Oe�Q�	��\T'�V�v�9PC����>�[�F@E��:�}�[�]��P�C�����ߚ̯��ؗ��u�G)%i�����ܧ�oMgC�wc����.���Q�ԕ(�5q�����w��rP��̩_c`@SMd�����;7>h� ��9���Ƒ_;x��B��	K�0G
��+��8R~��D�b��uu�f\�S��+Oט���x�� ���ٗ�Ձp���׆�e�V>�#�r��Y�ț~s���r���o�����$4q�"mN9�T�E��$�f%��
�P���1��ǿ�$��J-��PFlx�3��b7�%����E E#3<ٕ�i�0©�`"x���i5�@���-v��w��D�蒮���l1AG	QR!?."���  �-��拋��,�4�$~�?���b��0guF��"8�'����O�|�RP�nà�k�p(�."u�:��IÏ����K-�S�N+/Yr;���I�Bf��󖐧 ���ứAI3f�Xp6�~��-)h��0�b��{��z��iǍ�8��c'yE1_h�l>t9��#T7��o7�8�c8Տ�f���E��tP���+����=oY�
��xު�Q� r����~�c�Uk��uA�.Oa�ƃP����&��4�v����/�K@�}uYg�"�b��q���%�z`��V	���#���ٍcJ�	��WI(X r;Jm��E�2�E-b�aT��?��~ʎ2��i9<���!��+�q��9�	X�����)��,U��(a��86��>;7�Z[�1&jkOU��J�$���F:�l {�s���|�2	S���.��"á�� ��͸�B\�WFƁy��Y
���ئ��-�d��Cg?��]C�ж�9�-�Mȡ�Jۧ��xmڈ؂�44
����qK�����/��0����-�6�H����kF�����	b`�G`�+[ix*�p��מ�p��I?Y�P�;��FF�[��'h��͐�W"�0����i���d(v�+f�����h~�`ï�qT������@��C�Mt$硘�R@�b���\��I��YX���#Y�f6p����B��m餙&�/R/v�s��w`D�[�v/�Y�m{R�#��-��//�	M���v�0,���9�+�;��J�:7o�;Kn�۹<�(��$gb�Lc�3�@��i���^�g�ڂ�2w�*�t���ل���7�����~���i�
��*ةA����c%�o��p��d�.�g���p�@����:_&>���LZ��&������1%?������C�������R��~Ѳh���L��(��_(�NK����>���������{�.ߑ��h���1s��
�<����j�PQC�?5�:>�x���q/#�ְ�P���*$*rh�׈]�bQ1u�ݗ������R9ꃣS"�M���m$߯0¯d�l�^�����k����V��Х�	��^ci�����TT��$���/m2�X<��87Ɏ��3,���F�e��#�4���v��;�;��o�W3#����7V(�C��� |W�\FBY'w��Yo�P�b�bEْ)GƄ$TX�������.>�	A��6��=��Yv*�6H��e��:b݉i���V]Q� �p)�Cz~��r���գ����E�OB�O�1%+w3��{�|6�F&܀O�4F�I����7+R���[:5�6�z���i�m��ц:^@�GeҠ/���V߾0D�1a�;(�m.����%-)˯��L�0@�y��{3K���궣1��7�Of�_��l����$K��~>�����)��_�.33to�v��Z�E`��BJ�9d�u�9S����JY_��5TI��O"ԝ3[�%����	�6�
�g��Z�TD�"�V�V^�@W5�t��k2f(��C	q��oI��t�!����p�0ݵ�LV�d�d�.6��s�F�v��Ek�S�h��g�A��I�@��o@6�M�f��V����ߕ�B���W��<D8��#6E��i{����q���G��)�3�״nG��x ����J�v��V2y�X��#��i�l�����R��f1'5G�S�_"��6
/V�]*�$�W+��b��H�?�J�wʽ�ByjO�;����_ە��w��4y9�l�K��,-�Zuv�tV\�Cu�k��#+�R&�0��1ʼ����@�vT[o��q�G[�����KO�_�:X�g�$��x�7�3��ඝ�Ys���|6�d|:������D�(|��O�eM�!�16�|^��=i�T���B���i��ƫ�1$X�����ͻ�n�lޏ��R�ÿ�Bx����Kp��\���G�v���y"Hv.�+�KJŎ0ʨ�U^��9��yG� ���z�9���'0�;�|)F*�aY�O�620��I�|�[
�M�x�@�
j߰�x�U�?%�S(nZ���
ŝn��!wA�Hb��KD����z��J�誱y�8N��˅P}��TN�j` |:/Y�~�i��5��#R�D���s��_Q��<�x�J4�f���:7�{uh�G�`v
�o�_� 0��� ��@�0v�`�<Ÿ^�t�Z#�4�v�U'��Ӧ�KCbV�@�"�pD��} ̳� �H.Ϗp͔k��%\��غ`<�3�;�a(8{�e����[B�p�p,��\��h�`���gIy/��\����������yT"\��SsXcxa���]���ØFF4��ܐ��. 3V��3|UA�h��M�\�S��wƪ,S��!Cyn��[���=������	"£��g=s,���^��h��c)��r�:��d�D��4~����)��@2�B����LZ|�ۢG3>ڛ�n�m:�;ū݋XJ[fe}D6X�=3�v�.�	��P�s��+�L�S+%U������%\��uw�����У��nj��^鲷p�=\/�X�r�w���%[��=�����(5ui�˄�H���tšP��ID��r-���d�]�	�d�&���9gJ��[t��cyQØ`w*b�mF��D�����V�@�A�w-�;$�W�s�p�Qu�A��������P ���u�D��/+,���+h}����#�7��sP�@�o���|�k7w.JGk]��kM���_�?�$e�hǼͯ/*ĲB���$�a�:#�S%���d	�go�4��LΓf�%:���]�����9[�Q�7�[�K"�1��N㫨�0�@w��X�jݦ�O[e�M9Mޞq
VЯ�״�/n=��A^sk�u��	�BژX��O
���Xzk?�o��CJe3�]e�`�4��_����U���éx�\X���5-�t��`#�i��t���e����{����.9�|�3u+����bz����dϫ�I�/숙�e���g.��r��M�/#1�ꃯ�~�!�=��r�ncI��O��1��D�{y"BF�[p6��?V�e��h��)p�"E��.�"��j��"�i�؇�s���0e����E_��Q����]��Ro�Ma90!-���0�ӹ�҄j�8�"?��#����r��}'\��o.��b��{���(l�KK� F\�þ�{|PxgQ$C�)!qmv�P@/��
y����Z�dc��s��N&uV��ם�)ǳ�&l��o�/%�h����C���!lS��w�a?/4�[�㸍�y4]\�lm��G+JV���F��5���&�;XR��@����:*v�=و��n��wd* q��.���D�6��-u1_�
T�t`x_�gp��9��{���w.y��Uʥ]�ڨ���Fp�����'`Ltю���嶫#�_E��S$D��K,i��Ge�m�h��g�9-��Z�엋��K]vj۲�QM;�Ъ���#X,s��v��d��R\A������gO<��#����3���<�#B����|t�uX^J���
���� d�7P�����fI
��F8Py=�J��U�5�4�a�]N�hY.9wɦJ��7���Bol{��+��T��y�^����2g�p�G�sε?�:ۘ�?t�����L�r?�PU-F�M�?���K�o�2X�W�5������$C:F��QB۳����³��ȹM�h��T��I��v+����=��?Β�y�^�`{d��^�%��I�M]�!�r�OsHظj�\�.Ŭ>�)����/]�I�q>铎��9gQ�\l_Pc�h�����i�M-\��������~K�+ݯ�l� �{��Mܝ��\ӡ����8��3�t-�t?��e�מ S���DvX��M�b����z�Uί*r\ٍ� ��oտ�K�?F=��ܽch��H�`'R�엤k����B�j�{�|���ϔ#k�b��e���M|���SR���)8���a�U�g����@�zؓg�(ˌ���wfq'8�v��&�/o �h���?3B��اh*)_�Ҫ�nz�K���}d���Y�}��`6"�%$�@$rj;�`	�=M���FwEЯ�F=�.a��D�8eD�ؔ���5hU�/|�HuF�\�!ϛԶp�.ݯ?QcYN��k�O�P	�
�͉�����
t��Ƈ�L{��s��#˯�ވ ������?V��NonІ����vS��~��0��R�EpI �V�C7�f
ja�x���d�8�:���RV̄N3B�W4�U}53�����j�9[(6��26�Vm�����&���k��YN>PC���+
d3��	�g�{�� �At�p�^%c� [��E�*�o�ٻ��2�e�ڦ�{�c��M�f�7z�a��r�l���\�5o��Ь� �,�s;��Z8��h;ld��3��-��<~�N�`q����F.��:��1���/��!4&�h-v=��\�t��PE���h�_�F��S�2ɺ�؄�� �̔��1����	n�9�T�t�@�i`�+7g���F��R��X3;Bt��:�8���wY�X�0k�q��T�<��A��]����t���\#�L�vI�c#���F�[�C�P��gg*�TW�����(%���8�W�E?�%h3�u��q��>87��}
5�n���|�����	�����,on�8�w͐6r��Nx�7��5i�k\5�u�	m����zxaO��֩jN��˛~d���w��4���� �.�a����H/���5�R�����X6�y��"���꼕����)����V�Pu��Q���5�D^��2��/OR��r��TKe@=��������d����+!2$6�m�1`I�ߺk�_}����C���#T�4����]���ԏ��U�Tc�=uBs5A3Z@��mc5�ՑB��3+��[9=X����nL��',���ˆg��PRj��	�b��:ŋ�|!�Q�Y�@�]���h[�c�-Y�|U��@��N�@q^����m򤸏�H�LC�$�)VF��}�z��H@w㘊%��W
R��xqOfo�I:��՘��Q�M���顜���r嬴u���P�7a��#��z@1��)Y6��L��i��ءj��^��-�<^�s�g��^��t�_��gV��A�NK��:�\g+��V2��񕹭#�4�W�����!�+Qn�P�lF�Mލ��1�1^t#ן	&B�P[�33�� � �����3lB_��t]���ɭ�̞0K&<��*��n;��;��1;�g�#�V�.�j��/�@���y����<�cL<�
�����q��Mȝz�$��d�MOi/�v6�]ո����K��R��&)�xb��E��+&Հd�\;��
��o�|+�cF����w9I�(*cɚ��a����y=%s��>��p�θhذ�O~�Ķ��w����Qt�l:C��Р��%A0����̅�����?���x�Q�d����%��b�Z]�ɝ�I�l�
�,i�9N�%3�4�ѨW�B���@,��M**��:�Ρ�˂V�����*ulR��Z���J���!���b {!�4�O��f��Ȼ}�
�������G�����0Μ;~�p��.���M�#<d�V���z?U���BE$�a��TIML}�t�W�g��/N�Ӓ��K��ӔOpj���kK�d��@W1�~@]L��#�M�_&��a5��cU���k-�Y�}��[G�����}eE�S�Qw�� ����\�^a��!�O�v(�NNH��ݵP�bNd��]�EAo
��ޫ!\��חթuqF���E{X��*�|�:��H+"6�]�^c^�3���EM�K�Iʹu���0�H�C�ϫ64�1�2�n�'d����#��&]W�@�Y�\�9�Ǿ@�ޏ^�n���ِ�;d��]Q���Pe�g�wF�1ھ� �uA��"`TQl��]<bY0lno��.y�GJ�,9�p,�:��J!䋩+����n�ޞ��
fY�ȣ��Vw����E�SO�+yӨ��y��ʹw�AyN0zo����!���ܧj������r:F�G� �>vB^�3S��D�D�)]���b2r�ZR1&F�R�U)FꚘ7�yw2�$�X�������T��O�.�k�($WF�e���߬��㚴^�Gݮ���ɴ���w�nʔ��ue�w����  �)�
^����30��ڗwMz�Ҝ��d��B���C��[�d��\w��yb��FHB���4gA���>E$��+�"I�y:������,S�����������+ZVP\������R&�B�ſV#/��%�������3q^���S0_5y%��U�EvhN��`�-Ǚ��><� E(�o�\�ѪB2~����#M"@�!��D��hF�Y�>�Y��M�V�E�X� r>�f��m�B�D�e�d�95�Ug/_4Vu�����|s�h8��T����z��7�);u��Sۧ��ݲ��e���
�n xIKa2d��IZ1�~�6��!����ךE�.r�ƹC�|�C��D<ʹJ�K�pGn:6>|RUN�*ْ�u~������[쥽H(=M.��I1�j����k�GʩwY[�������%�������D6s:]
P��F�%,E}g���l���x�,I+���~B%�}��D↽�g�̶b��%{�e��H���3xс|�aoV6=|���޽�j��aR�*~I49�k��&���`�ᅵ	G�Ǐ��Sl�paH�1!'��X����t������pJ��̠6��ۓ��?���[_�4^f����j��[ t����r8�c��L>끵��r� X�� Du781�xi�������g�GF+)j{W� KN�j+�+/w�2rj���[}/[�@K��)�4t��y����{Iab�m��L�{��Q�6�gmO�Cq��\�|Z��h��P��dK��_���0��?����,�
���*�C?�0�ƼČ��H���]j������v�kt	�J�E��5>J��
x�i�����\*W*��?��!��{������a�[�B�۷�K�P�-���䠂!3v���#�mb��[���Ϭ�E��-+��ag2 Ql�j*q�]���l:+U82��@T�l6���ݿ��ӂ��ba5إ;��n�җ?�G,v�m������q�P'Z��~�((���bD<��)q�����2q���1�WCI�P�������@ Ѝb�T���|P���;��C�AD�?�N�vܔ��/���b�mGa���-�>��r+]Jh��$�k�(�cBu�'�*�����:�4ڎ�FR/wk�>�3�c+$[`����( �[?�i`����L���Gu�I	{�C"�aۡ]�mW��Y]�*WJ��%4����i.b�ܪ��D�9'�Z{�ә��c�$z����
�/�ty��M*� �h{�㐤��J]X<{�U3N�a�N�F����b�:��͵�=eP��O��P�?�*��s���/{4B�e Ō���c�j��
�X~�YjqN7IVj��� Df53���x=~�Vͧ7P��T�6Fu%3`�Ah]�lW�@��i]4E�9�B`-���#*�b�߫Iȴ�����<�3�S����ݣ�Ic� �}���]~�ң�AN��Y@`���9O]X$&I�גߨ<�}&��|Q3q�a�g�&�}������{D0��ʼKWCE��e:wLx��]4�%���A0)}5��0K0��]=��6�`e�½_e��U\��U�{oHk:�½O��0㧦�V*�0k���4��h'ޡ(q�Q��Y`@;�)|*g̚$=��T%����G��}8+�M2x �#�RE��궏�U�X��B�l�W��Q�����ĭG�ge�w�0��8�M{����T�M��ANf&.i�F_W@�U�R�'��s���h8+���)L9^�Y�p�~`H��Q%�4�99	}��>�]�s�Q:��  �PۏO\����@�C�u���!���=�_:�4��A5y�4ҿ����u�#��kUꞠ�xh�m�ߨ��~�N��is @���W����<V�EB(Ψ�3&��U�h��[�(M��bx���~�n�)�� ��$T��1UN�����7"o+��k&XX\4Ὂ�G.�����.�p'��J��AN�X�����y$��Pw��t)�Sh!R�ဂO����D�Rv�.�}�[$@��'+����d��J(Ɵ
�z�0z��'ᚓRCg� 9l�E8ŧ��f	�h�KIeM�3ʦo��D:!��7�TUq(�ԩPv�j"��Bg�Fi1��#���AQc����U��'�������#[�fPl�
������ʉM�ˆPȤ�e$�� ��6��n��#�N]¸^r���9�9]�P	_Yg��hBn���t�-�'�T�r�7H���R3���]�����<X�V�AS����r>�u�|^>�T*���[�a��^⏵d��s�wL�V¬ٟ5Av'�M�lʯ�i��QQX����B�A��2?��t�i�gji��
�6+uA`��ñX�̍�k��9�?Fo�E`Q(���#�J[�yck��H��BQ{{�T^d<� [���`����*����L�&�I�h��2�9jb���e��Bq`RXҚ�-j��g
�?�{��/�걼k��D )My��-�/.�6��'�X�i��1�,.
��Y�'y�>�e��q?*�܄����@����� u��YL�&.���6�{�ά���RE�����J#�g`�"�[c�S�#�<�D�
�:{ݎ����$U6(�|��ec�N��o�wj��ʍ����g��Y]�߫g"�7`J����Ά� <gs�c��-A��Z�Tp����[��5N��
�';*��	
n&��D$�=y��E���ᇘn�v2�｟����+B+~��������Ϻd�Q��QA���F��Ut])h��K��ݷ�n;Lc�/-����q��/�XD�~������)�>�2Vo|�_�*6`��ٔK#������>�J`ط�E�iB�^�3�ϩ ⡮8�2��Q�G�k�k���T����I�E������D�n����V޴b��������^L���.�t0��7]�%�(4ՕQqD��� C���~��X����P/��o���� ���j��Ҧ��~��Y���e���5���7�B�n�W�3(n6�pP�`��:)��N�˴x]7�}�7g+3��0���W��Plɗ�}fv8�p��E�4��0iK���h�w1�	����"	�f'J��ھ-�ޡ����s��(�J���TU����Z��,����,RN���bF�^�9�cc�ECuΙI_#���� ������W"AC65������t_~`�F�D��8�h%9��rkW���`�_>���4E5��\�b��l�����Z��_L�2�V�k�c�fk6�`�WXPHPu�,["_�K��aD��Ér(��.�D;�ٙ��	/PԿ9�Bׂ\����1cv�jKE���|�1����K�P����h���j�Mj�ۤӐ���6�9�Ȅd ��1�P҈�`�Sb�c����/�6��5Lؕ&.d|Gy`���"�2���q%k�-��w��)=�n{�P�x��g��FPѷ
�ՀQܨ��gS)���ӫVɪΔ�v�G�_��9��q �#�0Y�W�^�5�� (;4w;��YzT)h�k+˽|,��@5ʝ��ȫ#m��C�X�>���	œ���U��{rы���:�w�W��B�T�?��9@o�H�`n��f�x����Y�l�֐3[ "��~Ϫ��{�GR�鮡pu-��mşM	����n�͋*V9B<0ɐ@��+^M��7�������X�]�cϕ�Ŷ��$,���].b\9�$�Nqԋ��?(�2�^�W]t��U�2������x�-kDS���b�������{8��q�IX���6�rLr��}�m[���χ	aϼCh&]�'��P����+��&D�y>7�ώ�L{~�rr�>2�%�(}o`t�y�\�+�����%|�!n�O��_
H��L���������B���#D�[m�P�F"Z*��A)%���p��)�5�H�d^YoSc>ݘ�3����%m[��A+8j�s��S�y�c�y�������'�i��q\��\a��M(�xn��Ǧ�;��ܕ��_��&{�� C$O�R.��i�{{&�䡢�s�uր���1���B�;��_k	a��,R���)��ibJ ˴��?̀��%�J=\��#9��JCԐ9Z�
$v�p ������L��a%�6.W���R���5����<���s;�
8�3i�2	��Z�5ݍi��ѝkvܺp�mj}�io?�)��K(lA�J�|nF���5��{8��=�����dw�QR�徽�s��[!<��OT �ٲpI�p�U�߰Ӕ�Hn:7"?�4`��{��A��8�ήh}?��R:qWA�|跼G��B׬cs�d� ���X�߸B��{'�,��+�{%�ďR
��[�l�*Э����ZZF��qaH	x|��(4ډ�}�� 6�N���b����1��f����C2�G=�q~b����5�K��V�4y���С���o!�U�W�� �gTg��f�+x���P	���]Z	��Ф+W	ٲ^�M�T��W�4W��t�U�=h����-+N1ogci�褎"�ɝw�o\L�
�}B��� ُwa���q��L�����o:8���i/OB2-�GGT}�9�.Ş񈘪{���- �p�11?�X���A�[�p�
�2�	Z��G���g��������V�
��� �|���j���o��X��.UAM2'���/�f���t� �"D�D��V�կ=�:�]F�$%U���YV�c��S4�ȣb[{����&�EF,�l���M�L�e�J��ۧ~)�y���@N�3>ʒ6=rl����ʊ���}��W���D 	k�M�Vpl�6�8�դP�!/��&���#׆�P�?0؅�&�?䙬�V����`F`���,]���]��4�MaQ�u��ߣU��E?���2IZ���[��ah���Օ���d6�>"�)F%Y���W��0�\�Y��hC�fy���n%�WD���*����N�;��DO��H��|���k������Q�@aO�v�}�7=謤Pov���ćc������f���@9x�[ ���U���`5^�0��(��uCV�����c��2�7([~�{�v�����܍�� ��9[��η0���Re�+�-��Ȧ��7���ȏ*��[|2�E��3��^�G«D�b���k�����UQ�(_��u�&���u^A���-e�݋��b�+���^�+S�u:��"�ޭ����R���e��*�ޘ���7$F��g���	����h�M���5S٭� k;6�WC�R7T��6)45G�C�W*L��u��q'��Br"��Q 8��u����hܻvK�z�m�*���H�m��qKK墡'4�5��tNk��? [��GR�6v[teEn$0��7<_�G	3����޿0�S
���0���+�W��o\���Ыr]�K��ǫ�������a��W�'2�JHm35A��%QC��-��<�K�t���&�${  ��ٕy�}�@l	��X�r<�#����ρ��Ӝo��m���\r�\)tr��$O��x���"
�!�DI;�4VM���B���W�uO���r� �o(BW�Y����^�w��Q��O�~@_��4�Ŧ��Q��@A[���r��ڴ|��o��� 3�9�p.b��)��$��<����)V2�[�����3턜rWLX�ײ�`h��BU@1 �ڻR&Xl��^{�X	�9k�O;3�<����Zsk�'��t�IZj��l��o�Sk��kA�!Yd�d[����k�DA��Fx�7"T&��Kߧm��,�ת��N3m��W�4� sf�g�����5��y���x�]��=�D�R�(�&��0!| f����n\`'���~��C�&M����{S��x;2�5f��a P�!���������,��:WZ��g�;�ו>G�g$�(�k("��D.^�M��^t��b�s�B/�������f�pԙ�|eS.D�/��� &�ǫ���¹��=�2b1d�.��Gly/ҽ�U������^��(L짤� `�ٯ���FX��C����4Ha�����b��2r�I�=4}1]X��}�H�u-d�˕��B}��tٿ�8pE�x�N>iTp	���=����sK��.U�F�������X5��֑ y�������(�: <��3����~�Բ3�3�����m#�czh���P�1h��\�I���hp� �z�`8s¥)�ko����Uh����$B��+�Ϻ���?��>
����A�ǆ1���a��鴾D��Φ�3"Q��cN��R�����p��z���t��.����e,x�
��*����DoɆ��oJ����Y{1�eB��p�Dc8��u�ˈpng/��0���̄�����.1ڗ3Cn���CG����j� ��Zi@��"R�*v1�k�t��+<Yq�@��^�kV���������{�̡�m������Dr�6j����b%)A�}����`$�W�>m}!7�/�d� ��"�
lk�!\aa���}�#�&��(�b!KJ�h�yԜ�+-��0���Q��1�SU1	7�+���H�C��T���-(���$KW�Ԅs���^��z�9��Z�\���j���R� �L)�_�&r��n�L)�jdݍ�I�e���:�S���?/�#��-�d]� �Qb^W-}>�p�թ|/>�1��{�FP覫n:�U�����^���kI ����;���#j�a�I�y�L�=I�E|��E�Mj�5F)G`��C����>㻲4Ţ��ȿ�om'\C�
 ߪ�s蜆7���C�6|�b�#W�~b`H =Ӛ����;iѼ�ЯR�cƋ�JÏ�o��\y�4�1�:���F,B�>���v��X^�ɋ�2V����A�sp�ܘ�cifk �����h�U�Ծ$G��c�7͵gdW���������	v�1;��ϐ$C`9r�����VqO����9�ݓ��:�ti���BG˘��s 2J�uʝ�8 ����@VU�E�e$�"<A�A6��z�lPo`�n�W-��{��dô�nl;Q=�SR���=��v���j���]�n*�g#�
qZϓ���٫�#I���"�?��9FA*�ĦR��0�E�ؕ�ԫ=��k��{�Kw7��$��T^g�nO-&u�d�,F��L��PG�>�,�	曀WC�6�2��:K ��$��aF�*;�w�)J���>Ղ!����Źù0W�hFI�a�.�K��虞�����}�>XW�պ���N��� � r�1��Vdn�
���2��M�]C�pAt��mෞ�t��VNbD(<�aK`����c�8�U���~����c)��#'Kn��=BJx[7[!+hh؂^���ǒ��#�(�v��.��c�o���..���� �eT95`�74��N1-��N��ca����'f�ޗ�y�,��H��.,�˭L�a$bb�7z�W��aO�1���zX��p8'���>�����Ly���pVS��{�����=�8F�uA�w㨳p�+-��M��-���U��=w�
�����}+O��ˎX������FT���]"gu����L�����we��N��Էk*ׅ�LN~S,�!AhRT^w���֔��lR���GN����!�N^G	ڋ��VX�Y���j&�&���<���>�jܧF �]�N��2������3d��3�֦c����6A�i2`����_��=%L Q���~U���!�g�����)�y���J!W��%*�
����Dw�VjYw8#
��H�~�8�W�ozs|0'PY���n�u���H'9���"�m�@1�f)�c	����uM�A�6L~yt`�k ����7e��*�Oક�����-a�b[[�Ɂf�G���$
��^�6��0�Q'}3>F�������A�q���6�a�Ɯ���Ǩ��|�+7�ǀhQ����a��Ļ���͸�����˼k7���	bÃn����e�vh<s�q����'���/��0��M��[YL_�$������J {xy�TWk��A���]��>��)/�����G����_��	��V�>��	|�R@�ߣvP=�k5��%���;w#B>�����r	����t3����yFuEm/K!�n;�#�����z:��Ե��e�N�����fn���|��x���I��B�w��ʤ���$X� a�0�H;[�ĳ{ ���%P�+��I��$�A\V��m�/#q�0���؎�]�睤�N���7�k
�$J�j�;�v��W^���a����Զ�֪}��)�0�/_�u�tJTv�p�z�����t�%a���z����o_�nOux�X�Ȟ�/&�8-H�ɟ��ʱ��n���K�ҳ?��@æ��մ�qC5�7�I�H;���� ә��]c�4o�\��ι`���1���5R�i���5�M��13����mPK��Y#�����e�lqc�/�{���j�C#z�oØ�����fz͢��U������|97�v�Q&.��������/H��K�M�h�*UΓθ&�]�s���ccK=�~��Vnp/���/�V��X!̘��$�`��#L���Ȟ���/_fh����I�`;}:C5g��0���sxd��R n/�*ew��M�m)cVWM��_���y)����׏���
7߹(�`���� p[yV$�O��gL��7��^1���	�бH挻cR����j�.�p]���D�|��j��L�F����~0�ǆF�I�W	/�E�Vڰk���E����	����7������E����t�[J���{K߱�>���J���������]�ਦ��յ��|�� �[n�j�v���(��Im\�FJ��� �I9�f�h��J���m�XA.��j��R���)`�	g�0PC���%7n�=�I��7wg����+����� y�q\��Q�R�c��۫���D������/r��6x�TQn���Wd�ѧ@ؽ3^�j�r�]1t!�P���1Z������_��mf��j
r��e�4i��=fC7�O��fP��G5����[Uu���X���^KU�e
�A��T���ţZ�5�ؗ@ͩ�Sx��[��� @���~Y�^���]�hW�N-,ݧ�F:��z�� T���RXU���zfJ�9���� /�y���y�Pw�M�H��F[�C�9��"�k]�N�Ӈ��R�h��a����K_�s�{�f����,t��>�� Ψ�I���>�ն�n�Xq ����7�v�1���GM>{*}`�)Gr#r��BOmu4G���@܅���n�\pSҗXvnM�.h�.;�ճ���Ÿe�q�S����<�MV�����}�	��dY��`�9N,����h{��YK�p�v���gN�S}*D鷔L�*sȊb�.Aچ��νq���$��L�&�����/����E	j�%zu���Q�q���˻�����`5
UT?�7X�[���8�q��Q*�V�*�Om�[k��o�0u�b�傮TU��}����<t6z�`����`	�2���{U~�S�#�nj�Z�)�ޝ�(K���9A���tW �G���S�����WJ3�/_�ƥI��������Ogb��z'�D/����ڇ~~ .�����|��/R��,${��+�a8���qSS��
b�^Uy3�M��n��0χP_4�x����pcs;|��㮽Av٪��L�~��U)V.9�8�;�ǽ���T���{w� D8$�N�W}�e�bc�\��A֮�)_K�2�|+�"3���s��pO.�b��ɯ[��B����]�]E��a���"�7��Ac֭�>���. �M����:��H�¹F�D�,�(n�I�q͜�2�_����|�Ҫ��=���蟭_�?�̰c��n��<�Dn�	�Gٺ�ck\c(�^�ꃙ�X�T8�Rnױ�`��Z
ID�ς�<�~�����1~��

ޱq"��[��>�>z*W�� �%lYo�ecdpM��z��m�`#�������'P�yނ\^��� �h�4��}�)�k����i˗�s���81f\N軇n�X��w\tK�	��?����Wp���	:��#9��������*ð% :S[�՟~����ra{�')���.�rWKwG��=D�q�Ր���<s�O�Q�u)�)�Kd���\ƄZ�q>$��T�ω�&"ԍԆPe��U�>���������ᧃ�9�� %���ٗ���ޞ OK�����п%�m�7�$ٿ_VG�rßb�w(4&�y׬�lxIQ�j�T4һ����&���ͩ��b(E�>�wH�˚��c!YגV6�a�=J��!u�}`�m&� ���5�F�g�Q׾#��c�D���g�4ů����8�8�R��ɑ1�s�ԅ��)E�F��[�7���2�ug��=��u�ev�7W�K��Z>�zwF�i� �n,[�\��%"���6�v�\�r��:U���M�=9Ћ��w)��~��k�5=+���p*���uo��odX<����+sCv�iX�ه!�5��K�[]�s޺t�yy]�^�6�Ǳ��U��i��q2���g��MnPDZH�6��= Y�"ȇ��z��2�N�b=Z��@G�v!����S��H����?�6f�9>���jژ?��OevRr<c�PIxӯ�-n_����;�7`��s�dB�n�Y^�;Xɢ�ϵ�oղQ>�aEɖ��e#�4����<A=g��(d�6ۻц�n'{a&Ho:b�L�>�*�~��~��ȭ1�d�J�iB]�W��&�U��כ���+�
�*��:
��(0�~�4�t�Ce>�:9GK����9�u�KB��1h�Õ��.������W7�-��=X�ݜ%�Xes�e& &���M2��އcӉ�+�3��4�\��]jpԨ��%��P4��!����Ͷ��d�H 4`��f�1)y*OR8��� k��l��"P��̙0���?�z���ENClR#A_��/����x�y�CR�̐7|b.��`pu\��V����g��96 ���}���n^z�,o�Ddaق��*ѹOIz�$�d�{0a��NxS��I��)Z_M�'Hl7U7���T����\>�EI�Zn"P�5y�G`��sq�t�O�J��l���� 	ak��MS����B�^�|�d�ka'Th�:�8"lh��ѵ�6�T�'��q�����P�O�R�Q%,Y]�����J���_�퐔n+�������ͼ{�+�:�M�>S� ��ڊ�����o��6�C�KJ��S�W��w{�WA��oM��{u�'Q�������t����3�MTٕzaGT��CHz�u�W�!�(�$��=�Nv��l�ь(�j$\���0�8��BW ����}���%>����c1����E�(�q8<0�Nm�l&,X\�Ť|h�ryrj�͵�3���j��zG(AsJHv�W�'��m��0L���E��O�kRyp&�-Z[���^E��l�',�/�<)�8���S��ߐo�ؐ_v)�=Zdg6�~��%�I����$#��8�Ƌi��:������Ķ��A�a}$YL)�A��wM�i�B@"k}�#�=1�7G�R�V��*u��(}(�DO�Z��":����*!��B��U�����q�;}�"
A�=|�.�{�Lp;����ZH�m%��1��m�؅�<�����M%%j���#���o�}��u�wA>	��v��^�8�����1����˺/Er�����*$��	��b��,�W����!Ԭ��X�����0l~"�`�$�8\��nT(�3:�sR&!���gH��@��]�����k�+�?��iP{))�񝼭�u�E�^�}��cE^4�A�_~7����+!cB�@z&���KHĥ3H
�Vݷ�^W��5�Y��RQ@�N�]�ȳT_y��!���I�sF�'rpɨ�S0:��D�a[�T��U^R{���<ۃ���S0��k�[N�����
"ch�����Q�pvZ��lÍ9n��vz@"Ӈ��O0RK��GH�/�\�ɳJ�t�&�_��vWk	t�M���Y���W�y�R@͏���r>�=2�풡��8x�P3�c�#eK��?�>���=�U@[o��P	�&0�V��.��?o%�hb��M`�K�跩�+��98�q�+ٯ�~9��t޿G�4ѷ�Ͳ�p�3��vm{�&i90G���Yǵ3�!����z^�8^�����8����������m?�@c�:�Q&��˜��:�>�����=.��Ј5̌�T[���T2��g��)}{p�c����V!	ϧ4!��xe���D�s��O�7E�Q't�ϗ�ND��� ����k��UV�'��o\6�w	R;�>�"� /�Q�U�*٠�s��&L� ��O�b���c���q�n���)��9�+�x������4%
h���]Ą�����/8uNJ%�M��ג'nGhR1��=U�Yj3��u�+_e�:�Q�C܍���n��j�x��̇]�֨HF?/�
u��Im�"�j���wm��S�"o��X���N����B	E�p�;��k1Oi
�{�g�}��7n2�L�Ih�iG@3�B㰟���'b�	�6���ȤŁeY?��,Ypc�I;�a��3�֛�(�t��Eo�y՜Ŭ�P�͟�*aT�nq:,k�K�O���U�t���9yS�|A���}X�Vz�q۩�k����9wL���4X
̈D�|��~n�Q9�*�l�{��N��y�lR���0���2��QZ�������O�$h2#oဪ�`-� X���zE�7���ˍ	1����N=�`q;|׃R��j*3�+v�+._�i�ى?�:�����q��Z�À�z��r}m�EN�D�n���s;l��O�xgB�u����%o�T8��ݬFK��P4!�����Ww�@g`�@�-C�9�;QAD�q��?���X��NA��0g����L�m��{�e��/�i-
�0{ aX���0���Mi]� �N���Kf'��:}"Aȥ�<��;)���e�����c(A��Yڢ]�#0(>܉?�	G�e#~�hZL����:�x��Y��T����
�sB�r����ybc#��{�q���ې�Cv��G��|x��s��q��1�p������QQn!�{�>��1�:� �q�=�Z�� a8%MPc�����D���m���a7*~�(�,D�yɝL�V,S�kU�����t߹Y;���0_}���h��	 ����l��er���W�e�/�����)�Q���nhZ&�/]�!����7s�ѓm��E�ѻb���O��j� 7��
�J3�-<��?��7*�rc�e2-���*p8�� �Z�1F�9���3e�V�C]"9���0�N����uRH�J5Ȧ����n��>��m�k��׷��^LxP���꫼��Ed7�d�F-Ku �"ZcQ ���UJ�EI���t�	��a�F[��#v�1`*�^����J��4;���������Gx�[*�φ�1�I+ئ�6s�(���:"�1�6H孢���7���,���c����tr/����!ZS�f-��@��l�Hz�Uā&\c�FpВ+�p�l��H����6Ʉ��̉߀���a��hЕ�\V)O�������	���o0A������c/Ic�n��N�8,j���H�����T�E����\[�����|��a��v��i���=m�Zi�m�6���5؎��3r�M��,OM��,�P�;_���Q����f\x�?�K�gĿ�d{$*���ą��S,Q:�>�o�,K1��gs�$���?��_���P*N'ҿ�� C���#�����R�G�HC��L@�]h�=�oYİ{|A��e���2Bܸf��t�|���|��*������^����>hh�e�c����+��$DE�;�������Yd N�;�&�+���A%�
��}>�[R� ��op�(uZ�y�p��3��G۪3�'I'���^���E����ft�5��3��X"�7��zF����푫+7�PnϷ�D�}�a�s.�3���#=u3	���X��I��� �$9;J�z�S����Qq��{�zz��%2�\��Ƚ=aEU��U�教&���������T|ƾ+�ꠗJ��sW+�ސc[;��r�re�]1��>��@����3�[�l#w����B�E1�T�Rj�m�*���4k��3�?������̡��:9�"E p��Tj���T�'cJ���59 ���������ς�PX� \1�����a�4>���K�����ֶGj�?Z�� �������1��������}ƍ�Fb*�81�f4Ug`�8�`�;vn���)"S��{��z\ՙ�5��9OAS*e%�'��Yk��ɤs9*ch�KK�9��V��]��O}NF$���h���	���1��v�`^�;�,��(�4�fTQ�͕��������-�/$����z���� �p�3�Mth�ۆ��� $O%�b�V2?̯G+x].��e�K9A�C�R>�H����V��A�����P���M�Yf��TXk~��P4�("2��\ID�Xvw� �zi+�����>Bg���7`:|�𪔮V5�N��t�X� ��U��c����.��0j��7��b��+	K��Z�e6���X$5�̥Ad��q��a�w�ɂj�?�*|���=| q�+���
Ԩu�$5�wZ�^�Q��T�����zTi���ٸ��y!�]5ß�=��۫I�c,�⬰���	E<�n[;�W�	�*��πo��u����M�Ö#����K^Z�Uz1����#�Q�e��3t��z��e�2n���~b`ԅUTEBŎ��,�w�]4Q��%!
?>�H�i� �_�li��"��zB�;�2S���X�ы��1kF��2غg
{R��p9�"1���a���wsT���>�U��yZ�����J+<��qz�b"����Ԏ����X�jŽǐ�� w�<������}�W�v������Wk���4��7x9^�,�un�JG��؀�Ղ����D'���2`�/�~����&n�ޕY���qN��4@�x�"�3,Yu{F2R�pB���g~g�E��!�ѕ)[���Zav7��ue���aj;��I1W(w�J}�U/Þ���Z����_�N�<���3�m\�`�갞r����e
�-ub�G��Y��G��\��T�R8���gP:�/L�9x���8f���g�_h�-m�
���j*��B�1��t�7qG ���?����y�!@SƟL7����pfH��y/= G�����|�.�K������`��yJΐ5�I�? |����h�I��Z����V�h>���g{u٩I����pZ�X�:, �pq�A���&����Y�C����f���{��"��T�(�ZVd�3M��gC��\�i�GV,y����E�� o:��7�D�����09��:N������Pqgi��sń�sİ�s������ɋfzۯ�y�j�/a����a��9{e�dbh�Y�-��E��(�j��ò�EEce6'SC1̮$�����I��� lv0U��7����/YI������u]Ҡ;�H
$ߋ��X�&M{�v�XMOCxw<Qh���V��H�=2� zL@��X��*�у�V���[(�׊^}��ak2a��{�Z[�9���,N��q߆qb}�!�FN@��8�͹�BssSnR�ڜ��B��z	G���w�u�$"6�/�}9�-��8��]���^��u(ʦF3"���d�*�}B�`R�l���WH$Z��IƤ�e�J>�0O�P���'}^�'~:"6��<�}Ɇ-< vd�[;����h��c�@E~z��kG�Va������.�̺�H�j|�f9����"�sM��G��GJ��;�Y��:۫0��=����-xh5̮�?�83��������!�G��1$��|���"��j�h�9C�x���&Nl�$�F������DW�`��py�`��bӇP_��H�p�U�!_W�,��/(R�y�c0u�l}���,?q��)��E�J����f '�߮ �{�Q����p��]��?۞w�h�D� �d��>�M�L�f.k�f���dQ�/�NʬD��"9^�sB��0>[�Q���&Ѿ��`�y�Ͱ�~v�[�s�S�s�F)$Olp~�` k)Z��3�%3\}g
�A�?��ª��EQOд�,�G|2˔�g6֋�|�n��y���E��|��7�a����o[��s�k0���gF��$��6�F�}�id�X�X~�C,!����5xI��G3M��c��d�j]DdM�H�B�~���kvʄ�TW��.�wm�̵H�������8ۄ���(� l��)�qU�<u��g"_���<5��Q�t3l���`�յ�H��H�c�cP��CT��3��Y�<+�A���#ؑ�)�j�^?֐җ#��-@���<N5��Ȃ��Z�S�i�>�/&�)e�S�j� ��
5e�m(z���z�0r8l�2̈́k����I�1�(f	'h������%��%1���;���-�*�Հ���j���5���#%s�]�qPMf�B�������ǕE���'n��Rz��RѨZn133b|O�hP�΃5������d%�g-��e
q�B<�~��R�s5{W.:X�&Ls��]a����"%Sv3��7�X&�g�E��B�a��t�t�$��h��Y5�2�!4�OD/@s���*w]��wO��q�L��"����엥��w���9 �j��H���څ���.���(ۀ�DXE�1������)"�Zp�����祝�2��.�<{�;ô�%��*n�ŵ���"�gY/MP���6_=��D�EE2x���7��9J��Ra>ܡ�wv��E����%A9,�3�m���5�"�!�Z��a�߃�,��
���ٛè�.��쭟����Z���4�6�5pe�,J!�p����#H_J�Cc|���fM��\�{锑h��w�1E��Ik���gR��a���D���i�je�cz+�򗃂8�����J�5|G�y~�$;W����Xd⊐S[|An�z��h�F�A�q����D%<�>m����d�3T"�ͅ�rP���ӟ�)�b�^���[KD��1�"��9D�(�o���w_Zp�	���O�b���e��������	���� �C"��]�I���ܣ(�$)��^���5S����������͉����8�;��ɑ��2�u��y;��}1�A�ט��F�$��c�Ƀj�ǁm�E�AG�����͕��旼,�kJ�E�A%�P>ɐ�ã�0������T�qi����J�ԅ��M�i�jִ�(�i��E���e)�F�82AY<�*y ��Wp��݉�k��((A�s57[<�&+́A��+�R;��pQs���l-V턂���.유���])�d�� �e����=��|���F�TC���M�(��������vK]�=MYO2l�H`�.�d 6dֻ2^���$����Z;H�H��j�{LQ�N �8�F�ϮDH�3T7X89j��s���3O+;̫�R���9�%��V.) �U`|*{����T�;�g�5���_�p���fט磀T�~���+��I!S����H3���&��߉Ɲ�OpG�g?���A0�\>>� ���;�ޜ�|�,���n��l���[�WH� 9͕,Qϙ�F3�[�����6>.׳G_9ſ�ɜ�G �?�a�|�`1[Q2��}Z���d9�vVH��������*[�>���CA���0�'��	w<�PID�!��PB�j���v�(�c2����	�֬��ۊ(��A��+�Tej�m�FJh2����Ź ��?�v�� �e��C����m h� ��m`��^%|ъ,�L ���(t����$����KJ�;�{B*"�]�i#TA�t��U	4,�3p�L�����������'��\���2��M�6``_�Fi��
�Ir�2</���Qk;����q�#ם�:�=h����mܔ��x��xo.�S���Y[e O��>U�{�B�B�@���v�i�y���LX�y��DdmiSۉ�Դ��o8��):=׶M�ʱ?7�A�w0�x��P����d/R�X��j펌�S��Qz��Q-s��J絔�93���xP~�jLEM� lc=4�x��-Y�Ro���$��w��F#�����c�[����(�����x܆:�쉡�<&:�\�?ZLr���I�Ts�~�`�T�-l(�+ [�Hj�&�[��
������*���Q--�~�h=�.v`�b[�ף�p5I��{{B���Y�et�3�ރ��&"���r]� �a�9=�Fd��{�Wi��Д� [��`�I��vA���A���G������Ҵ�V�SA�$p쭙��qR������[��ab���CT�y�����%os7w�w�<�;RF������-I�N��[s�&�M�U�-�'�*ܿ��z�"�9.��y�@b�NS����3CP<o�t���(d�ܖ�M��Ы\�G��UK��5S^EL3I��i��h
�A��` �$bgl�_].��k_D�)@0��ϒ�eIIX�EI: ��W�&�D�ݻ�}q
���c[c�\��Vt�'��ϴ��/d���l��6^J˲��Fw����f�1�hڂ�g���' ��<�S7"� �+O�?�'�� �o~7S�	�X�U:m�e�;�W^ש8j��o�}WnR@�D�n_I#2:�����e"4N�G�eVgl����B�N���������|2;�8���~��G���٠rW�J��蠇s�گHf#�~�G�D�>�00�gu��b���`]�i>�S~�2�x6�w��P>ur�v�v*@A�*�a��:��"�����e�eߴ����������.I���X�6��Sb���{�5Jfna�� �m�s=��:1J�@I.E'��#u1X
>�/�<��ȓ<�`�=����.���մ���o�E��1���@y=a�| �(;��A?��ֶ�5�jҀ�&�?��iH�K���A��m���}M}P��ߦ��ƶ�)vU��:ŭ @�Nl�Q�<��f����BnV��F�&	w40+�"�����%1z�{������iҿ.��.t�Ҥ�w�n�����X��������Q��KvR������O
?�j�A�ZȈ+7.�d��L����O���7��ms�����a@&rlwz�9����r,V���`�6e[q1�w[դk�w�� ��c.�'�yr��i��5��Լ���}�h�����ɊM&X9,:�JP�M,N��7�U�J��a�b�N�ٺ�uo��
�{b�@�)����@o�8������NY�h�d<�޵�u6�_��߄�Ś ����uiЕ�+a0����<���"c���@˷�f#>>�q�Ju��x��]͵����=xd`�|��":J��M�q�cE�&���p�nն��/o�{ea�NF�x&�6�D9\#{�]��p_�A���D .p�Ĵ��[I`����6�����*�ime?��N=h [Α�Ҕ�vw^��V���W���F�nx��cS��?����L���xS����QR�q,4�|?�n��FG�13χ����슗�� 2��[8M�E9���@�Ƃ �P���t��xٔۙ[���g���Y�.ڱs�SZ��Q��ߪ��\-;D
͓<'�����'�p1�0m�z��_�h�vU$����*����*�X�kG�{9�0ғ׀�X���Q�Å�Į�t���F�~x�|�qq��P��z�=x5.�Ëe��wMqr�\��p���G��"�Ʌx(������K}0:�/t�!��&��t�,6�rVcz�����Xy�+{����G�� ���n~sc8����ȉ�
���B���ᦀ���(��Ě���#f�P���
;:V[����U�n��N�̵@��b���_v]�������e�r�S�	L����_Ɠ����Q �o�;���&�Q���c���^��gv:�N��k3S�L
YY<�{�Y���L^������'�
�\@��D"'`�T�`��Q�W�ϊB%0Ћ�����Zƍ�/���p��6��DK�.��U�Aa�)����-�9j�K [�V�T`w�g�l��cY�e4��X�d�M/�?N gl�Ԇ��8�z���9/�,H�)�&�P(ʋt��@�������h��sdH����]�6xy��?>��4��ӣ��͒^�j!�6��Bȼ������&[7�v=�I�X��� �b����#�Z�G� �0�.�Dg9��Q�(�65��&�%�m������:��3���o���Z�;!(Qj�A�I �O"-g� �*�xφ9U�`d��̹�(%���۲�i����-A�kA���������&��0ak����
���3L�AM�����r��B�<�6��#s���䏁�_� z}%�g"��<O�B0�2�4�������J�Fƃ��0�:���w^��޳&C�A��i�҂�Oi��nE({ü���-&��_�G��,*�����Ul	/-��p��\��;
�������~���(�^�Pʻ��o��C���=,����s��1�t��f�K�����1L�f�s�Uf^���Wg�Re�)Yg��yw�sJq[p���ZM����t�߲��$������YY�纫�m[$�؄���������}�@�o"�����/��'9]�*�>N���2���+�k����h��B�Y�EΉ���^� �<��F>�4Nv���,@����)G�7��XE��Y�/&��U�']����ۘ��5�N�@o�q�ж������&��Z�p�(��l� �I���@˃�#��D��kXˢEf�,y�$�3]Ƽc��t"�9x�����C��K(���>�w8+R�x��_�K��`D�*���C��g�F"غ����%�z���ݥ }���bWo�+�8<���NWSJ����������Se�IZK���_�C�EV����c�y�y�yT�ͧ˴b-��>O��������Ӌ#h��5.T����q	�q<f�<�_Jg�'���� �+�˃�<�c7���OR`����Ns��'��M�/s7ɽ�{����\qQ-5�ء(4�+��/�-S�˥�P]����-�~�YЁ�#(� �s�2�q�2�3�K��,�$7ۧ�����i�u�|�gԮ���p�b�%��X)E�|�����nc�i��d��sL:%��h(@\'�j@2d�#QH&:V��������ڔ����aU+s׌�u���^|Fd��ZcN�8^���zG�K7��'Zź�� GHs�M�h��rVM��'V���''�xR	#Sgm�^Ĵ&�J���3��&��6ù�Pll9�M�lJ�<�@޹��l����c�~.=7>�HPD��*�^A_8ӥԌ�qo�m|Փ��)� ͇����/�ƛ�����J|{�������C����G!�ci�p
Q6����(����l�6��)G��r���9{tO����#�ciBK���jbo��2�)*��U�	�R���Wŏ>��I?��M[�,�%T�z��|��I1E�S�/�m�~E���~�--�z��*[
�jǛy�L +=����e�n5�UҎ��o���|��������Y��c}"^O�vJء�\��k�@�D�K���\Ywf-;v���i�Gfv¸!�Z�W^�3Eh;:��`�{N�������5��F@�����nw6�3�3GM'���i�t%��|MGt�4����R8�v4%Dg~$��ut�P[]���K�w!�ou���z*���=�I��wTͻp)/^�]�C�b�o!�M,�ㆻ���UG9�B�e�0{U̒}%9ȐZ�/��ҰC̞�IZ������
Mgt�L�Y�C"B�7Y隺�AG�Ȏ���ʁ�Z�U�0�My:O�����+7�^�B��{��ͥ�:� ���<�*�L,]bd\�ga,~��O~�|g��p�����𲢎�I�n��8/��T�`P�Sz�{�1	,3�t�l8�i�l���!I	%;��/T��(�񛶢*w�� ��g���q^�t�==��T�uv1��K�g0������/��q�̦#��-���=��"�g[� ��������k���7N�-�7p���oU�e\�]��H�B����t�1�m�z�T�I��<����?aN�e�@7_�tT�V7[!�:�]��0���ok,!0MO���<�v�(SA��޶^@�N�sO�2P$���:,+�]J�<G]�D�@Nd'��b�]���Gh��=z����{k���x�T�"��o �A��)��a#T\���¿3�=Mh��vnS�:}ja\�U�l��R:Y�j����unM������PB�3�YF��[�f�u���P�%�(se{��&�&���n"~Z�)��$Y$3СS,+K?�P�>ޖlq�WЬ��z`� ,�D'ò��D3�Q���d�����Ĩ���*��Ke����A,;�����5ʈ�k������tv��#��X��!g����ᏻEh��U�(���G�9RBH��W��
���LW]��i��fB�m�-,(�b�؂�N\=���)>������V�p7	��/:mxv*60_
��RXMM���i72:����`��x�����:�QS��9O���b� ��f���ֳ��$��z�-��]M�Zߴ�����b`�ƫ&n��UP>��\L��?�F��������Mpݨ�W"!l>������/���Y�OK��Ӏ�Ħ�sZ$VhO���p�Bc���d
P�
�sDAjg�d@e�<��<[��m��D�����~iv�4ds��(�����B��%�&����'��Hj~B�hQ���x�K�,/׀�mc������+���<���~5 ��u�lZVq}
�h�nXG��u��Ɍ=�{L�N�Cd���]��cX�>��}�Y	ϖ���<_������e��}E%������,NwI~r>�T�&��7� ٌB�֖�B��=�Ƹ���ͽx��*ɪ������y޿�#Xn�[Gx�T9��;ʝ�4���PJA/gm�ZA��Z�.Q�6��%P��
�'�wC�[�v���ҵ!���b9Lm�qg\r�I�p��&S�r�wj�]����%R�WRh�ol�j�4 4�dI�@�^a��䁗�w@$b�����p�sE�?�T�d���}��q���D�2�x��6!�F9)b��%��y�����V����ݰ��:�ե�9C<�a��9�w�Yl2C �Ǆ�y��+w��0'.��X��m ��ZZ�6��,�p�H �\��Ѥ/o$?.ܴ1Z�dG��@�r�MyeU�ٖ�yq\����A:%{���^s��}]�Q+뾅�J���Q�0Z�D�b$���d��{L5�)�$�A�KO�l%q0c�8v���>!{���f����V���I�k��5fP��Z�9ƞx�V�>���h*���q�5>6M��j{x���Z�Z��[�EJ,v��G����ǺrE�_E�$D�����%�T�O|�ބ��c���L/Fu�b]A�H(&������y3����o�fT �ǥ�~�:l<ڙ�x�e�)!�����2�U�)�}���Q���j�j/��i��N�R���
�pk�<�>}I�.��q�o�_����UB8XSii�iJ�b�����v���̇Ł,p��ܔ���1DKҕ��;5c5�XC�~"��62�[�"�a�,�����[��E��#�[yH�V����'�Y�
R�k��GD�A��h�/�$�ە׎����jWdq���Q(K�Fq��$WW ˟i 2Z�����D�.-�����~��h�z��8�ΆAH7��%C�q����:�
Ye��QL[y�I��Yx������:❚�#�.G�^a������ALG"h���7�K�s^���fjdo +
��c�[���,�̋��7�+���������Z�i����vL��ݎ���B+���J���27[c�֔b�@*v�W-�꟱�]���M% 5J-��p/a5�����&�Ȗ��0��{�Aa��úe��>GTi��3��1��Y��qB7qf������V+���d$g�*N5ȭ$���{o�9@O�ԧǿ�v0o(q������1�����%<pI�� @���6�3ۥs�X��7�#c&'%������9E��BD�Q,ag�?VP�7z�:�HXN�׷��i����|{�AH�|��2�G�!䓗��t T�R���������ȹ^,Q[�������p�l�Ҝ�����\�%xQE}ky�LZ���<	���N�J�N_^��*�eR�~zqww�<�
�Z7�? q͈ ���aCJ"�(qh|q���~��ģ(E��C�n&>���fׇ�kt=ЖN	�<51��Ǌئ��|�R��e7�H�Z�MT;�?YryU�����{ye�C��p���1��nOR���P�3ٷ��f-�a���Ҷ���B�/-�i\�d��-uf�����wEeWe�ɢƼ{�o^V K%��"��ܸ����"���g�C�>!�ϖ��������G�ꅙK�Qr���a>��y�-H��P�
jgk���FvY9�1���|p���f��Z7  �/���IG+N�;y2/��@�d7flL�CEЏ�z22�}����g�ed>S�+�&A�#!��9*@ZTގO$f�'K���J�ڊ%
����ѿ��Uc�M�C��@�}�W �	@r׏x�����aw����_����v�U�D��� �9����zkF��� q�$[|�)�^? ������jU_�8��ӌ=�_���;��o�yW���&-�t��Xr����hr ���F�n��Ӎ4|��r5�����'F��QG p<�Ԛ�"ɻ�>���fXf�e��;��M���Ĳ���Ɏ\���.���ܙ3�Ԍ5�bZ��$wa�SrڇZDR6__�`�jO��mb9����`�%����>�U�/��9�1ߛ��q׊�D���3[G�a��6W��� �LO7�s��ߥ�/s�Ry��_f�)�+�Nj�������Ƨ��,��߭�� x%]�4�>y���%Ի&hJ�;���b'!	��ѡ����'ISd��r�]�|bo:�%�7����{/���cw��`�O���ʲ�[���*��T
%�����#��.�6U�3��8��п�EhKi��y<&���(�sŅ�%���$z�,@�ꭠ��(l���#ͥ�գl!B&N��eQj����UA��Y��9
Xej?�8�e�1*�����
e�5^����|����/���,z�Β!���:WhJV/ �6f���?P���g��bj羽�dU�Ri�{�� ����@�� ��m:���O!)�>KS�F���k*T�?S^z��}ݞs�zۄ3�Iذk�Qt:|\�8}Ԕ�բ����u�6��C��Ǟ��¦U���0�K��H�?㟢���5({|�ZYT�8P6�I�����F�ЎmY�]9dKu�gd*n{�0Oa�HW�b�C5�u즢ێ�4�K�J�į��4&�؉D��<��BD�sd��*P����0����]�Z�;r��5t��K�s�M���`�k���|irlBA�8.�Ʃ�q�a")�,+��h������r��M{�&�Ԝ�ߎ�A0�g29�j���li��ɖ�V���k�O7���1�k�Q���+�.��h��
T�B��G7.��O�Z�N؍~cH�Ӭ{�JR7�m�����Ub�$���_��}��J�M��)���{��f�3��C^�|ɜ�ڡB��)��^�����"����MGh�!���.�f �U^�S��'a�Ml��@�����1���z� �{��l5����cMH��fwL�v`/N��k�f�ا��|/'�Md��s-�\�?{���b.��#�w �+5hq�5���8Q+��SDo�~-PO,���\�]�?��^�ય!Ѭ�:'����cq�/����Ox�;�f�p�o[�l,�GH��Z�l	�_O�}f6gFO��	�'�����p�_�^s��^��Sf.	��x�E���wrH+(���fG���^�g�F���kx�4%G��F�x�*X|��1x����GR&|f�g �s����`cgJy�y�jk:1_k �SlP���jTeN���Y�C�%�%�ge�`�]s�C9��j����U����3�RKN��n������	����<���?�����+���N-�TJd�1�ͺ��+�����$	=��H"�&��@b��n5�Z?H�_��d�<J�p�%7���L~�m�l�2�=�����sW�狡-�@^f�"�Of��H�&�gp����1�/��+W�1�9����N��J�%���cA�/�i)CS��G��q8�o����k&������Խ|�<��%��9�^߲��/b*u�4��ۍk�שּׂ��"�r[ry)�1�a~�S,���h����k�_�e`ڇ'�X�l1�. �C7m��>}���uq�����I�2q�sV�8%���d�O.�z���~џx��FSS�7.&>��)�� ~�6��S�X�-c���_4�C���`Ȼ$���;YDԇ$tֻ[QX���z#k;�ϣ�®9e��9�����Z
�=��G*�Jk�M���`q_��A�BO��Y�W�e���t2s��E7Ri�Ť3M��\����
#��^��X�j�s��U9�����(-�[�C1~Ę�}��	gG���W�{���'Rn}n���B|��B�٥�� �AY���i�J�����7D�].�NH��%G����)���|Z����;�B�����$�F�-���;0ᅾF#����R�������09�0>@mMP9HWFv�m9K���k7*�4=߷��z�l�6�fD+���x�U�4���C�!�V����[�R2�7*�q�у�V/��<��|���}�ܞOьə����9��y���#"J8P{���]W�2v� U��k�ߝH��F{�؃��B�9����s�����K�������ʝ�#��GX�e�q�H�i��N�a⛻WA���Tͭ��݆�`�Ө�r����W��t�An�6�44����
St�$�@S
���U(�	�sw�������k9}��NQ-��q�"}�6���\6cA��,��)�\]��z~�	��+���[���$���m���h��x�D�q���~���}�$J���RcG��D��  p��^�|7f�z�:��\�0*7��݃��$h����?������M�9o�?n�F�|dDғ�QɊG�3QSA���58y];��;��:�:����<9�^-���̔�/�tN��l�����/��y)��eO�i�K�a&�R�2n�֕ء4�ZJ�M$y젭�����i���D߹-1v�s�^K�V�_X�~}wf���9����z<P^�	�Svՙ5�?�:���\�o��]@�B������ڍo�V��ӋUi,|�s��c��fÙ�1}M��y�J>�v]ĠlУ�K����)'�j`HGYx$��xs��1̻X�L8�}�<��ұs��5�Gon�	H��U���& ��r�o��rp�*o���E���>�}��RzT�{�RET ٯ��<�2a�7[БdH,�|T��ia�?'b8����A�w�Sj8	T)H��a�v�VHL��qCB��W���T����7b�1\�<�t��vu�n�	�wԽ�w��.���%fF��^{���U���X~d��n��r4 �O�T�bM��V�F`7�ˉUxatF���(X��'lt��En:'ф6ۧ����5v����y�I���I�9�����2&��*An��F|Y��K/��L�}Y<���3L�;q3��b�?1 ([�ݡ�����.2Z�����W=��Z���AI�2�c|.�E��K�bȪ�|L 7�ݼ�7�J�:@�,E����e�'��W��$h��H�j�l�ࠁ!�����Mt����������ŏD%1���=n�x��~Qo�ZK���	.R�%�db���9�Ys�-u�^�2(PTj/W\�������u��:F���Q��R[Qs�[����P�^;t��m�/�|�j�l6�_��g��l�b;==��VQG���(3N���3'�p�۵�MOd�f���!Z�F:��=��#��s�����%$C�ZC���f�q]	͟��X���D;��N��������!d__����+�*�8��(��~���I�7�9Qfj���
PXl���w�=M����?�q|�f�lR�3~�</��`�_�!����%_��",���͹�
�0�w���b�XRv���òv�z7I���Ыc�k
-��D5�g�)Ϸ\+>�ॸ�!Ͷ��ȃԑ/��p�] �zgQ�4d��r�0�oQq>�=`f�>��j�R���,򄷪�X}��?�1�41(�=��g�1Ax�V�Vhڅ�(���dyAu+�d��S��#�4uლ�0G
���]���^�j9�@C���N(��mN����.��pDϬV�BQ�o&���%���J�2Gm���6(�Ĵ_����T(5|�s�`;�ϋ!�8��㗞[����@�K>�x�ll"˯B��Z�[�U��`9��Uٔ��ެE\Bѻ	u�Tw1ŀ�=�m��w�Z�'�3��32��a�0�+���:ѯ�D�\^���D���}�0I^<E���4֥U�1�O���?(�����s\̊���U��ɛ�Dδ�j>�k�k�D����@���E�k�?���w�����b�3)��rt�-뉑��p�x�N����M��u$?C�H_&t�``|p��
��`��_��[\3V�t/k�o'�=Br�IV�W|����%ʓʝ���P�!�3�#F1�e�,�; �)\S��q�~�V�Ვ���?���l], {}��Ø$ML���r�]���k�a�L�P���~�*�K���y�������'��@�p	���F����hHL"6�k�l��<���j�XAlB]��CoZF�B#~d+��q��5��٪��nU���Y�O`H��6�ԆY������٭<�p��a
�����9���	�ʸ�0�H��T\]������m���V�B�õ�Z�Ć��nqGb�Jjz�BUqV�x���W����UǮT��w2�8�&���z�=0� 0]Ԁ�N-شbH!��7�n�q�ok���y2���|� �%�I��[ְ_^�{c�9�Y�����A���uڲ\��P���ػ:�f~�l
[����=�	�L<�\�O�a�k���'�ؙ�eh�9���[��O[�I��i����b�����K��F��(z�k���ǹRTn%���=�b�`I�,b�BD����4]����ӑ��!�$s��/�D�8'�Re_��T��r��h͇���Ǎ.�Y�xT2owo�Uyq�0�VJ+H�=|S���߱H�T�Y6ػʴ�r�u�f���L��"��s��|�rс��"��ws�s�^X�榧{��2Q"�A��Bj5"��sI�c�A���N�s��N�:�~�6���ʬ"�n/&ZF�G�0/0�a��SÝ" �7}"hL���W�U
�p�ƍQ�np�jk=،��@��9���aE
�^��])��2��v��u�K:�q�0}�֝�KN�n^sw���<�CO�%���5|3@%.٢��p�̍0��P�a�Ն��M��*�U���p�h�葔��<��{?DZ�d��V2�Ă��� �qa��d���<��	e�4U�G����������5��K͵U�>��>��7��f,#����d���s��vB^�uu���~�_&hOWjB�;�$I��G^q]�O�k��&��NH��a�#Ps�%�"E�
��>a��<y�����~ 	�pp����e��S�&j� ]������5�8/!
�K�Z6��?F~��%�Kz匈<�"�3@�m�W��0�5�O��p��{��s�w(��CGL:+u㪠����`�*z�%\�a\��[�\ͩi��I���g�0>9���v!�
h�1��9>��\k#�?}{+��6��)���RN�{�rx��I��-O2?��G�@[�+�3e��tKf���|C�Iߠy'�������6�KE�7߲�4j������56�PֲH(���X�ߍ�c��,�vRv&V�-LG'[��%_T�~D�WU�t)�%^�G�����ף�)KH}�x�)K D9����c�18c���S2�\H��g>e"u)�>� ��n�I�yw1����M (� R�v�Gq�`�Ez
h�<��;����8|�:�g��2�6_^���+�kWs��o�s�6R�X�.M�TY\�~!D�4�¼NӸ�*���~B��f�r���Y��8�w�i�8�� ��]��S/-��<��ٹ���^���_�eo�Ľ
&��:8�wx�;�����;;�L�K�+9e�騵��A����H�
�%�����!�`��0,��qh7���8����N���m����06�󫀃g��s��Zn�I�_V��Q\����5Txq�$v0��ḁ�@V��DKR���(��V�&������i����iEe�"d�0)G�Ux��0��� ��O���xy��U���:=�E��~)��I�1\aF'ʵ�9��q�B�./p۟Z�����a5e��]!ʯ�2�{�����F�L&�cm��+^ywڬA��C'ݔ�*r�ha�;�r5d-�|�b^j$�('3�����a�uI6	w�xG������vyQ�NN�IuX����<`B�2�����[���E���j�	Z���-m:a݆G�My����L�e���TŇ�cwx� /��� +���w�J���P	E���4�;k ����1��:���g��K��cdy��x�Ġ��%��}=X�N����P��d�ꦫJ�fP:��
aȥ�K�g���9�=� 4-\6��+U;��
2K�$��Ko�m�>xҖ�9|$!O��t��S�I]*?��77hH�!\kR�h��q��Q��)u�l��+���l��j����O�.�J>����пWR>��K������|7V�ơpSH�J=�C(�֭+�"�wm��,\;�>�7��Px^���ѭ�ٽ��0v�?��ޡz��A��w��2쏇�3��)]�g/���������#m�y	��}'�Li�ϲO�X����H�����]>��p	~���O(]���So����'��lN�h뿪 i7E>�Ɓ����&���c�Ta���n ���
�7?Ǫ��l��~i&�4�j_ٯ��-N����V�b� P[�� n�@�s����<}e�M���ϩp� <���[>4Aё�Kev��
�&�r8]%9�^͘x�鮣��(�QYJ�"SJ6kN�����qF"r���k���{����m��4K��� �Z ���e����5�*���ϫ��i�F��sf ��2��*~b��N�چ( ߂�F)��Ϧ��sf9
�I����(E.�/ʽ���q�w�q���e詮�~~��&8_�cy���Pw�F�0f�*��ye45�Y�/�N�_����1���qC�Y/곎ݫe�8�	���ӛ_|�x��G�F�ME7JwN۵,�X��굴C��5�{Z�a����_A�r\���=`ekgrE��&��S��R��*��[2�\.�>Q<
�p�ߋ�G��}�-�B}�FṞ{	����+|��¬�C��К�������� =z���d
��Y�n�f8e�7cz:2��I�K�\%Sd�.:�t�y�e�� RϷjѠ��W�ؾ���X�N�U'����%���e~�Hѱ���(w�J��������.y^��0���W��{���
Y�58��������J�ь=���|�NK�8�O.���lC0�tj��
d�;o�9W��+�m�p>����p_lZ]*jX��g�K%(Â
���5x�;�o^�.��_|��ef����W���*I�h��!�Ycr��t��n�/+��s,+)�&^ >����n����`u�'�l�*"y%1��`+3�9��ܠ�]w��*������Ţ���$�Q蛬g�Y=������U���p����[LT>�K;��]]���W2�d�i��������1i�P��ʹ!��V��?.Vi{�`\Z.0)}?I�L8Yr�|*����=��|���+$^>��7>�K��X鄄�9枿��<��
��i�<��pW�	䪳0	Ģ���*J`쓭N�ob���J�-�I��7옵*�	��������M�Nr���C��gL��e�i���:�d�tָA���j@��F%��W� ����HM����Rx���%WXެa,*��,CO��Qo�&T��} �dU{8���?:�s𯊕7��3_��� �b�+ks��yaQ?ߎN���8��4�W�>ǤKd��d5s�;yv����%@�9UTL���
��L^��]
��	y�q�*�vJ)'���9���$�,�.�ҁ8�K[`�G��8fg���6�H!\�yC�DT,8��&��CTV=����A쎿��L-�H���b_\�mo8&�z*G���lA�?��?%�����`��b�җ?��`=Ě�iO�,7�{�kD��E�L��΂j* ߜꕑ�TW���*`"���G�=}@~$a�JM	?���a�b�y����9!n���I� �\�9F^�i�n�Q-
� �լ�t���#�?J��c����k���F5�T�iV�Zl�~�]w����`�G5����M��YԘ=�K�%��qt��0��JB�_ߦ�3�b/�X �����".T�lWBv����ZP�Tnft|uS0N������,a��!�����ʚNy�r��&�z����O� 坙J�
*�� a�.D,В�*�4�DX�k+�ư�A/d*΍j}g��}�����ۧ+,R����%�J�I�I{G�_+������2FR�J`a$���,y#b&��Dlb�7���D���e_������|��V{���Gd!�1��jqvB�[�^B=���S�`~��i��rHw^ u\��d�f2�Sx����5�4v7#�L�1�q���o�
�N[!��̸JȢ�Mf&����� ���~�_K�y�&Ɛif!>�0�	Uy��
������r�W|X��u��P���~�#���w����1~��������\��e�nբ��&�>�w�l���O�M�m�|\(d�oc���[�x�\�+FccD#��Ŭ���׃�hs
�K��\ҙ������X�'q�o��+6_�qI�G�ȿj�/2Rvd�`琬�T?`�h�����-`m�F�����o"��I.ᡙ6pA42I2&i��T,0À�`��-� k��6ʿ�oh�E�������*=Z [���ꏮPG^܂���nt�ﯫ�~�o;��p����N�I�*\���t[-�	.�$�u�PG���&�eF�K%3�%�1�f�����n��5`����z�|�S|���}�@>�S]2�p��h�@�c�2�Ƭ7��!�W����"��Wc;L����c^
(��/m��9	 OY�S�����<q��B"��J0�;�I���;!%�w�4���\�A�����1i�W$���ܑGi��a�V�\�� � :�m�'J�_�g���m��|�bQ�8B�?r<����ki����nP�ywKh�'�D���]��ݑKYc{/�xN��8E�?�O\��@��< ��,b�������Fe&�BP	����jQWT���gP��m�|�S��tlc@+��N�9:��EY�]�ĉ�j5�HZ�E�O��S:��'�I�Lq��GQ���8������	��hW��m��7ƌc�B���{���XL��j;����6�V����W�S-���x��&�y��X�Z�V:M�R}͆�q`A�7�Y,5i�8��O�?i8�B��}7�z�}H��KL�O[�O\%�[��2"�тJn�H�e����4f�Z�ؒ�ru�H�y�Z3V�aAx"ѧ��:9׸��;6L�u0@�<���"�j����1ଋ��H�Ƶ"�dt7DɄU��(�G���SWr��R��8���4�@{�4%��x�����F�휼ey��X<���$��jPzM�\�`��ٖ�^��ǎ�E��k���<c��w�����B@�u�7��&�J��y��]�2��V���i�r]����:��)C ^��� ^t�Z8�v�J���q���M����O�Yw�]��:X&{�,�J�y§?z�$�;�F�Xs�H�fSTv�da(>�ѯS�!�W��Ue��=�� ��u��O�촡t�;����ʨ��њ��G�S�F�D����j$:�rY꽈�L�ߞ�-�mq��K�TAި�w̜����ch7�2��'H�t!^l�a�����Qb�+R�uZ�n*p��T���|�BI�%]u誊O+�����LI���K�4i���7g�H
Ne/�������[v�qq��z�7�����یd5���Φ	t�ǖ��0{�զP�772�4����z�"�^%��8N��9�\�h�B�_��>���ݞJ�q�q�Gkۼa�R�;�*i��qw�e(����Vq$���!�E40�"�S]?k]k7��[0"��w>�zd߬�z!ϟfC�0�Fu��{.�A�H�+�}u�F�O��c���ŕ�=�y+��$��~2m0�}�hʥsp�����C��2�f�!6���WbX�^��y�Q��s�Sȸ�T�T{�t�YD�Q%��7vՉ:�P�C[P<i���ydj�%�U价��:� �@=��:��n�T�(��3�_Szy2��@�D7�$Pę!������Vw�3�8�6Iڣ)�u�޼�4A�j���n��u����,������6�C��I(	���@���eb4>�"s'��%V�e���6_ ��P��9�FS� Zy�3�����k���zC��%a�\��4%�}���=���vW��x#�!�o,Q���]��E@w��'(k�f����h8)a'g_�$����Y�]�����K@��1�9=q]O����U;�I�J������e���N�:N�²$4y��\�K���(�-������!{� H�>�@�/vR]U�%d�w�-w��϶/��MQx�b��U��� ���s���4�5�����*�mM�{1a��s�Ԥ9c8s�h��P���	,�by����g��Q�I2X�Q���H���zVȔ���u�1 �����j����)�zU,k�u��&����sD����͉���ib��brz�Y�'�����B_����tZۨ	�d )f�l{'�+-֗e�)SI�PjY�w]�p<�<#����4o����(7�U8Tt����4�~、�@O&����FXN�c�f�_�WKɣ.�	�_�z����E�>�&�Y�JB�H�a d���y�=�O0_C�4]��6(C�Pߠe�
`v��d/�T��|$�	$�fe;s܅ʕl���(P�)����o�Z��e� ���5d� <'���mm�3ِ��g0�Kf���P8��(ؗj�R�
a�ݍWk�7���H���y|_"gZ�Sr<<OQ�r:��y��$J�]Bj�}k��˅�OZ��~E��	�{���>�L3���Mr��⣧^@�JP��n���;7]\/�Of�KEfs��g��7x�B�>��rQN���]/�*��Q�Qp���n�0�j�X�j\�%��r)ٛ����hE��d��_(�������7�z�"�6�%�_�E�v��3x�/)�<�A���KlΡ-ڗ��&f�cs7YKV����ȬS\+�|��{�K�e-����%5x�r�'�!$!�;u4�yz��0�H��>�9O��+T����e�ZJe*vpLM�!���x��-,��EB7��Ah����X��R�^�v(u��t���X0_��U8�{y<Pg���_��p̦:wcD�������cށpc�B�Xִ�v��^�]9e�8lsK�m��RAS�tX���o���C��_StNۜ<)��ȴ��甥W�P�;V!�Ͷ��4�~a>��_}=�;KGھ�J���[ʱ?�ҞV�9mnq�e��c�m�%��b�m�q<��=�.F,�Ji��G|i�T����vc��0�JV�C}B{�rx,r�B����U8���S�����P֌��ɧ8���0���h�(�+���P��u�&��q\R�:�g����cE���ڑm���?@ ��J�W�ⷄyX�����Ȇ4`V�!�ِ��<�L��&��u9�H�4��,�����L!�� n���&�[������d	���.N5��c�~���p�zT�{��;������E��іz�!���`�ǜ�h�a1�<��=�Z�mS��,gQ���r��br �[3�R��d���tU'�d'E�LMzb�e��f�	�[R�"�O=$ⴴ#(p�*O�75��hwW�#�r߮$D�����ĭ}CM^F��#���<?##:�}͖�&4�e��{��{�&*��M�չ�2en�:ΝK[�.`������jJ)W�9^���){7e��y �����Jb�ͫ�-�VJ)/-�n_)=�$���L����vU�ƪ�|���A��t>�:_wBL�v꼞Ę����Bi;WO���i��遊�#�]�mSr����$��xb�]H��>��#�������NO? ���h��u�g�����ه~&(1��L�|��Ey���:��)�"���x�OyA�7��S�1�����ܻ���.�pdw������c��
�6ĉ�De�/a*����M`@P�G_`-�^ᙎfU�?c��U��&�ȸ�v�/�M�
̺i���]�MB��`V�.* �0�$v!�GgM��}��uj�/������	��B{P^�`�B��7~2F�6�b���Tv���u���R�����T�C�VT�v]H
G�����RA�RM�Z��z#��P�	���쭴!d�v����4��w�4�''-S؟� ���_䴃�t�;3��MQ�
�k�aŇ$���;���r;GŊ�2�>�daT�ģ�w�����2,�Li������y1Z��Q�_4�gІ�c�N](�x�M���H�����zt��߾l�Ft�^%܍�]𴝭s;�	@`���^�2�F�<OyX�`5X�.ڳ�,�cJ���F��B�d�H���y&��;֩%���akřt}m�(���[<�oG�l�aA1�HO�Z~�/,�&'`(]�Ph�ؒ!K�V�O压�+�~���s̱!�Z؛��4�������N��\'���LUP���Zh���&�l�i�(oH�|u�[k�0K[]���/}�����t%b �x��;�|+
���^6�\W	��jr���b�
jRc���2MqL���{+���t�5ɨ�UE��,~O�P�_��7%�1E���3�).�;�pH����*����+�O���d�.�7-���`4G��5P�[��Xr��ũ&������'Ja e���e��˩����w�@�a������'�g%���]�@���n������mZtg��3�ͺxD�*$�m�0��hUF�B��*d��a�������e����D[��<��F���&���4lщET�w�G+#��9|�[x��m��%W6�=����^%#�#��Ւ(\���-?u{!�"�$�ن�&��K�ƴ�fKEj����"V��`���~z(�=EM�/�l�+��8�t��fLNFڪ6m��X��R��
���7����l�aY�VU�G��,�G,@.�Fw����Wev���vYc��:6�Y�½>0�e�>�	�"�k����^�3��.��\�wO;�\yb�R5��9�4��^#��b\\'a	�0b{�Sa[�\	�̥
5"(TW��n�W�L�Ql��Rf"�~S�|3´��%����k�_��!
J̐�{���3h�ԗ>^aJ�I:P���l�0�Y�&�oЖc��xL�w�߭d,���5&B�/�Y(�S)���B-N��k��H�V�	x77cJ9��m�J�>�1��W���0\��C5d�g���V���_�	S�b�A��"�Je�dɅ/~Է��pF_�!��D��:�=�hѪ�p<%�EϜ�Tᬰ�w5�؛J�4��a	��~�j�U}�~o���]��A�f.e�7I�X^�����X�����>R�,���ͮ���$4�*п���W��ڢZr)4[u��?hV��HUx�1�JX��׏4�����WR���4�!9�u�Z��?9gܾǴ4i�]i�}��2!�����PHX�����pJՉ^^6MK#�0�F�}�����8��"t(	Cm����3���Ng!�P�|%�&pn�[����O�A�ZvX�`	�E̗��	5�l�m�����i먯�X�ߍ�9���Ͷ�e�����gKV�@�ڈ�ۜA����xly 3�#��Xr��=�EN'K�i�!f ��
���v�|������^۾��:����Z���V�!V>Ε�y�яgZa��'R��V
��h����o��B���|�˂�.�Q�: �����l|�3)�~H�+&L/�z?[��i�4�'1�V
5Es1�A���G�y%� ���qi.ֳo���,F�^�O����6�T�W}���Dj���;��ג�~V�AH'�fZ�Z[�YS�%���k¸����0L�ɽ�d�Z!��W�6=-a�\��?�t��E�c���� ���@Ԛ�fi�����(Y09�Ⱦ/ ፝G"N�ͦ'�L�������|9�Ĝ�ᙔ3�`7���D\;RS�th�Y�* �����+��0_'�R?���P{a�ܮ�R�ׂ��F�4)f�U60۬Z����o&W�|���
�-bs��(�:��H���&n��I�Դn�� 6��|��)��8i=ɀhɴ�����[e˕��v����od�<��;tf�����@����-,��
����z� �@r������.����ȕX+���n��M�j�Ɖ�i �-����j�c
.D��G�kZZF>�ӛA��ěƳVn�y_ϼ�2k!5�Y.|�����L5�q��s�7���-)A��vs���,9S0���ڽ��ǌt`4����\���(Ƥo���u��'&��X��l�c��Sm�?����&��o�O@�; U�2�s�t����L�@�x(<��M����D�e#wr���f>&
��s^��%:��R-� �
҂2� D,єԜ6�s��o����	��C{+����DSI�iN1�!�=<q�{
2��$m9kAy��g�W/� UbZ�P����ʜg�xz��X���a���.'�07�(I�|����0~r58t�?m�ɤ�x ��\o�1�er�o��T��E�u���q$�:ܚ�"|�H��O�����,Ce��:y۠�����6���x��$s/�Љ9L+���2�_�X��f��kS��@X���;�Y��5`I*J��Oү�r(� �p��ޖ]9��~*�+v�l6=�G�|�3�x�T�n���3�/��&�2|���P��p��ơ��k�.���}s����=V�#�6���&��2���b�h-�V��ɾ�쨆V�)7\�5����rK9(W]��P�f���݄At/���A@�g��,�QK�xa�*�;I���͘�9%��#4�q�'9�����F��ڥ��~��*Y]@A��Qi�����i��h��t��ٙ���q��_�@��[��}��s18�fZ:h��řm���4,�fN� "�*C�M�&l��3-)+�Kf�T�f=������{j�9S�:C��J��ŀ�f�.m�K&�>9{}ط�dܧ�X��Ê��]Xi%ܙ"
��O��w���4�Tx��I��� pŴT��T�����O��C��"{M�U���N8(C�'�=,	LQ��ٿ����C�����)M���^ �:4�z�O���N�{�^���CF<��!i裒�x��J�*9J�Wm\�(>���
�h�tsɩSj��f=kf�6۹Zv�s!�/��4�!kw��@텔8:O#Y(��`��f��]�O�CތVZER�Ѥ������v���v��?��d�� ��6��qs��ތ�%P�K�9x��T��z��TC�T^|صڦ'��'5��ds
��DN[%��#���EX3$���e�P�MAa&+�TԨ�vxNMу)���b�>˄}����W\�0�׋����c�0�pG`��3���V�yш�J]Ly�@:��i��%za2��R��c��� �1f��@��a�F!aux`5�j�@�|����^���F���*Z	�O�z��-�Y�pְ�u�kKp�ܮo=vV��V}�}�$�`mZ:�=�O��`�\)�(���*�I���
�?lJ���]��r>����L }�!�:zG9�x�ބ���Y�ך t��|�9��"$Gw�O�&~�?���|�8�Հeo��-������'�^e����
+��W��LT�E��CV�?f�=��?Τ_�x���q�+���I�έ<ߜ67��;UJ�z���!�x�N�9+B~L�5�+>���2�ּԧ���/�N�������l�(�6_���ć:bgѦ�9OT#F<���(A 
5��	Sb�Ȭ�j�x5*�� ��Ag�C��R@�]H���ik5�;�)p��]��u�Ζӧ�4K�E��/Č޽�	��hiDz<��ƃs ���l�+w�0� .��0Tr�v�]��>+�@U�c��X��8vm[��<R��	fR�����.��Y� F]���'������tO�|��pE=e^�L���셜^F%M@[V�8Q<�/\!��ަO�R�r��g/�ko��W]ݽ)�
 B?�B� �1�/��eS�Yb�>�6ב��S�Q�9�1L�#G��b[tAT��|J_�r��7D$ݹ!X��c�8�j&I ��6��Q��	����
��YF�c ���N.9���
���S���\�9����T���27��h�IC<L���F8*4�WR�RN���	�e
AT����f!߽��@%���[��l�K���˔"b0���8��æd����\ 6n�E�"�Ga����3�����a��<],���O ��w�1�`�9�\�nt�?��N��L`O���n����I�B�A�&�d���F���%�>=C'1�4�L�ĵKI�N��k=`j�dǥ�����<�����]��9h=�$gZ]������I���	.��|��^*h�D쉜���&]z��X=q�~��s�3d��6��� Ū�u8�+��6r1��B���lș�q�m�d���@#�ʂŪEa�C�@?���n�����;��+����~��6��E��C���)��j�a�+�4�K�m�����yd (qD� G_*w�\�e�� ��*x����V<hu\XuH�`(�>Q2�%I�j.x��C�;5�,a��r� ��4��2��ob�K5$df[G^�7�k�����r���F�ۉ�`�Ps�ڐU�y<��Z,���k/��S�Ro��b > ͢(���Nwd�[�i(��'F�ڦ�&��(�8�ivf2� ����@���F�3%^�Z��l��Yk��l\�9���0x������]}�沎sg$�?�v��	9AEM�J�Q��.��n��짅pX���u����n��	�]e��1�CQ�D�k�7D�!Zu7�9�u�X���l��6�4��29�]�����I6E�%h�s&(��L[O�$��2D!�'/�)Q�˚������X������%kʙ-�X����p���1̆�dg���R��'.�JkF��KW˅���/l���I/�i�ϰ]Q?3�$M�^�-�}�S�ד�ǡ��ͷ���RF�k�4�)��*�{�"3 ��o�s�9���	7b����J�����dH��`������� ��UcT����l6�0�Ե��;qO]b]�����70��#S��#,E�JT��O l�:�,��rf�zʤ�tZ���h��P'�� ��	�d����i@�U מ���)��� 1���[���!V4�8xu6D.}��C9�ؒƻ���t�Ku�3|��&��W��6Ot��B��Cf�Db��]�3�ygF[�~�
�]���e��SO��h�/8�H,��{��(���|?��n�.����2#%��F,�a�5ًb@���$�O'���~j�ºO
�=��H��ry�`n��]?`\=v���(�r��<|���G_Mk(=$C��8VW�'�o+�!ɟ�H�f��j/���{�{��A����ELaZ��r,Hn*�y��H�+^h�� ���0ZM��[* =� �TYsY�ƿ���Ry`oz(e�<jo���! �N41�"TC���c~8��筷��~(73��׳����2be�OQ�0_?�HU�P����g�$m���ۤ����&�PĄs4�pCd��u���EA�sTE�u��QK �Q&�������|��Ȉ�|M-�n��:�ߢ��^���k\�����V�2&�0��r�q?��ȇb��;���$�6p�u������3s1H5����.K�� ݃�!.��3��
��C�ͱ��m�'��*�Jk��V�=����f���E^F#��E��2��U�}1RE�O�ud�b=z#���B���{^�y@��E��sq�_PO��WǨŶ�2v� A�S3<ƃ{1R��B���^�ܶǘ�n�vl�Ԏ�ms�Iv̻?�hAi��G��pzA�ff����ѡ�H�H�5�J
��0����ot���8��Y��L�ˤ�0����iĺד���F֜��R������E���,�Ziջ�W�?���z�+�7r@�0ȼN`f^�2Y����!�®]���6B9�4j;5��&gHG.�6�gϒE���t7����A
G�e��%�o���y ��>VƝ�#�J�9 ���Ż�yη�)�yl��:/jD�A����=)$���B�>�eKO��S`G�[ ~>��������Cov,߇h��A����h�\3�@=.��ɏ&G`یo
2�2� /����45�aI`�HH�S�ouv�9�ؖ��"��Z��OC���vf�i�!��U~��6]����vrE��Km��K�=*ӝ�q׵�m�E呇��E�)�`���=d����j	|=�$�%��	K���l�^�s��5�g�����`��j�4�
��fw���"2�8����S��C�;�s
r$ ;��Ү>h�	�X�\���?�k��~b�O�ldp-�&�	@��?�W����b������>V��|�L���T�W�,]��S�.�F�M�v���!=��C`BBv�Fn��$H�ğ!L����#�s?ӆ����lBo��4�X���-t��)+_˘3�z��gUI�2�H��a�{�wm��x��M�P
�hb�KfŚ��x�4wY��p���ݦ�+��$��f�k&`���#[<�|�59~}|�����,C��|�S7�ݸ�2�6����;
{1fۨ_�1Ղ�]$<�o�z
-&�/R��5@Q��:��pg�����qJP���/3�H�t���I�]:�o�l���Y9F�����'���T��v��cL�"T}#�\����U��@uvb��sEf>�u�
�q�#'�ik�I����x�_�Ҫ�y��dܲ�@
8`�:-��ēő�k�W6c������*(J��{�#m��F`S���αhPǀ�-7э��%z�+3=Hw�6�<(+������*B��Dǩ����@��1cln�/x���jNSЄϻ�Q;#o��>ʔv��[��`��3�>�}�s�������H�׎��Pa��;sL��F̉(�چ4"K��,?���?�.'}�	sر�:)�$�q�R+��Du	���Px�H �6����t��iX�Α���8h��*��1�'���y�@����7j���/8�V�C4�J%_�V®IWS誁�ߡH ��z����>�`>�<fA���A��=:�Z����W��b�6�%���q3L���:�r}n�m��s�8�/^d��������k��7o�}̓	,��{���g ���{*/���] "r��2M�N��'�#eA��w�F ��Q,�+����8��C#�4���{|
��y���Y��mY���z.�9w"V޽?�X�B�����mŜl![ �8���ݙ�c���8��#ڴ�K0Tܥ?%4�4\U\��)��y[Ƶ��!9H�?��İh2����u���n�)i�
欋�D#��SO���>���%9���<�h��l[�`W4p��w���|��B����A��r4�Qd�y�i�u<�ci�y\qs�f��� �1�E=�(��h�y����xh��h��5ҫx��\&��_����.�%�Dv�J�)��|_{�*�.������m�9h�mY	L�yKF�@A�I]L�c��l����hUNۭ� C0��2g�t;_�0~5�_�����X���O��W���E�lZdT8��S��&�S���Df=���=XOV�����X���@()<�t.�'�aEP?㊮�P,_�4E�ġXsk�㕾�V͒�����F��Z�!�#ޥ����+/�N\رE儵�5�Uw^��ÝY�养�@��]g��
)&������xܼZ<i2}�4����r��k��1�����8��Z-��W0Y���"�)�b^�Jh�c�"0���Kti����+��W(F��ǫZ�h(4�G ����(��BN��=�������q3���c*=2��|+SR�ױç�D�W�Cy��ߠG,�G/��+�l���[&b��%B�Y� F�J.���7�t�+&�Ly\� �k����M��m^����$5D�����7�.�#��OMi�13m<YE��|�����������H��z,�Fm�l���Hd����'��a��С���EqM�,�]6P�M�'4_6Y��<�X�Ӽ��r,>�i��Nc���dy�[�>��ݧ��}�G�d��U��	UyA!���7���$0er$�*�]�L���e�IԐ���߂N6�h|Ӵl�6~zr7Q �~���f��)����tlr&U�o��E	d��꘡��@�V~�'a��[v��tv��m��*���� ���I
�N̲|��>v7Ll��u�e��򥻿��V�I �r��'�e����K.���k^VA }�^� D�h�;8o�F��-��w^_���Mg�K�U�NO�"�_{�����m�F$�c �9�;����rgӻ��M��k*òe��'��"����6�����!H��N0��F_:^_�K���2
Qe�?^��k�{k5"bP��t>�ֱ�,���u,Ȫ�Ek�;��(X� �I�!A�8Y����c2,�u\`S���4�D����� /�P�eԝ�n `�ц�A<�1� *u>�۷�r��C�bX�鰷 �������8��6�r���HV ǖ$%��(Fow0���3����g�qJ�^�ߕ8;����Ӫp "�j��ϳEe�j䶗po� �@T#W�ѭ��d�<�p=�::��#��,����c84��W��M3��p�V�Z(�B���oļT�S�3bk]�ٟ��a�E�#���AC@�%�;�=	���ɭ�E~x�[x|�g�����(�('��3��s�a<�r�Q�K�Ձi6f���z�������M5oM=��׀nX
ߊ���DO����ˀ����r ���4��
����:����A/1�. �����-�L��1~ �� ������%y&f�z�9��̔�N7+����H�N�T��%�N�wb�J����X�"���Vm��~FD��;q
 N?(�C\Ra��*H�	�|��Ct-d!��	����^4�������Hա��@��߈܇��/-b��XT����J�،��u �Ϥ*w���q��������^l�g-�����%b	:~��a����Hm�����ȟ��c��ո6 x��f+�}B9��bi&>��E�ݍz���G�AA�z��hƭk!�}rr�S�zY������x����<#����"=½�q��`A?1�%z+\�k�3a�g>�|%�fk� ��ɹ�n���
��Τ�9����؛vu�����k���.c6�H��sˠ����K��h��B%n��a��_���T9�ؽ�r��`/�2>��JO������:F3��!��\� ��QY�|��d���\��m�?���Z&x(�÷�1��+=b�R���. r=@�LBx�'���p��d�h��U.D
��1^�[�=R��,�]r�=SI�۹�D��w=�6@�lmV���O�t�I�C>����֨�\�1�͏o�i9��Y�����I%�v�?�[FI�㻾����U<һD�G-��K�`P�P��\A�8�~O!�D�Z�;j� x��,�M��m
s��|��r�N��H�ĕ���32bɗ�.�\X� O�BKfA:iK�!�ҝ�!��G�F��I-���k2��M~S�Z��|�7�	��t����^���-��8���ך�>o<U��}���%�%��[��C���6v�����~(�K0��W� i��Z��P���$�|[Nu}V�
�N+V�R#9rj�ܛ]�$�}��B����B����X �c���>�{����q�b�Ec��i�&�O��~J�X��@q�Q��j�a��l���H��C�W��fT��/L�_�<��[���wh��Jr�z$�Em��jp�^���98�����:��P-k�aQ��:g��0{8s�4rw�mᾨ	�E��	)@j G���>����@u�lG�4�W�N�+��'B���n����l`+�&>o�Ȗ��x}���O���VQ�����Hq�zA�^S�7�w�ʜүh�&�w�Ulf�����p�*Sd#������I������X������y���� �uW��E淚8p��!�iP^��/��:^��3X(?�R�e�y�J-9�w趥�.�	4?�裂�B�Y�׎A�-4aB+���@V�!D�܂�|2O�vc��O^���T�l���C�<;�2'�!�=�l47�Ӣ�_�GP��uC)��sRng���3�I�RM�5���cW�f��w������&�Pg#6S����]�R��d	�6j`�+�=���Fpѯ
�x��g��v�	4|�7���jB���Ga�%�ё��(wĵf#��T��{"�P���$r�0v���p�i]�Q��s�ߘ�$�e�����@UDg�YQ�J0��@�d1,]! "���L�+>-�L%���^��V�j���5�8�mG�{���#m�����.Ya*&��#Œ��X�����~�a'�bW9y����ɀmk�:��p70Q����yt�c3���a�7�1�Q-�٢ �;,�JY��VC�C�Dt�rI������5����f�>;�&_���� i�[p�7I�v��TJ�/.]�zw�;�q��ǅ6p��ޮ�C�A<�w��p�6fDH��V�#v~)I]5`h�6��͝,�J&��T�����̍�SQ!}�`��p��z��-�
�4p����O��u ͩTJ�3�Q=*��#F�'�]j�3R�\��*1��o�@2�<�NU�d�����	'��_�7%�x�h�qi����.�C�F���n�(�#~B�d�	�+��H��h�鲃�9�n���+
���ԭ���ǰ�����X���� ӵ�V�(��Z��)m6�����д���E���¬:��	�N>��ߞv�u����t!_q\\Y�N������s��C�� �,G}x���X�V��>A.��XL�B�h;�0Z%����-(��w���5��.���Yg�>9�i� �~y0�%S���4$��3���ˤ�x ����7xYs~:a4��1�j���Ա�i��λ�5��*�І^p�YVƀ1�������$dBD�3H�T$6$�x��z#��1����ŝy�}>2y�D���2�_{�6O�ǋRJ��o��2�j��=�Iy@�tL뵄qhW��v��բ��gN��k5A��r�`���b}�ק�c@<�w�`-Aj@?��w�-E�W�|7���J�@�у0��%T�_�����-6�H�G$M���Ni�y)Q �& ņ1�	`Gt�Ga��r��3�C<���V7t�C��yQ��o�h�^��>dI��������x������ѹw���m!�W?&�8#��DaHI��[�M~�<����ak���Z�iz�W)�~���61�c�J��po�_p3�w�Z;C���@[f+B~��K�'� w��\�'��z/�Ù��X\|�(Y�1�a���V(����H>��g�]�	�]�?�&�����B$�]����jS�=��(��k��-s&�-�u��b�=�.��cV�\��F���ӜsN�܈L�*E�b��h�C�j�d�k��j�dO��by����i��S Ʀf�n���b�v��nxͩ�ݢl�U��ֳ(=�"&B�ü%h�`ng�449p�ת�/�&Mr�T��x�+�� � ��)�i�V�