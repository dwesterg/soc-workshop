��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���'gW�ӊ�m�K�&ϐ3���&Ee�8d�p��FB�|~�t^�T����E���"%Qn�Y��.�nR�$U3l�6���O��<���n����ze�'�{��4��O�b���p|��D
NK�?ZQ/6T@�c��
Z�<�y��y�2 D�g%^�G�BP�~��$�.s�S[�d;�����������2���1{���#3j4!ʇ��k���n	�g<$|-q�H=�L��E��*jgS_�X�xa�/���oϯ=��$�w
�+��c�r�n�t��vK�捉�_v؅����OS]�WZ�(\�^r*�,�&m��W�ZŽї����v`X�������\�� ���0�NtM���������A�x����j+[b��k4�B�B�b��nϞ��(�2��W"�b֝V�q�3��2�=���"�ع��Y&��
8�v����5�����x�D�����S%=NC���:ت=��d�qk�O���y6�C��%N�hi6�����.��5�R+�C�?=2�!	�4("���[CA�{�.��8g}fI�V�7;��U�O[��Sv8Ō�3eH�>0h�m�^c��ߣ��@�g�g��0�ǵ݈�Y��4���zC&�R||�Hj���L4� ��z��Q�ŉE���\���npo���EUwp�S�t�8���A�xl�L�BɳhM�{?8G�=�=���P�h�C���kQ�r�zk��0
JUi?Cњ�n���a���x���Á�7�	��\�;�:}��X����L�J�:���Zt����3R�zѷh �~u��Ȧ7������[���0�� >1ת;�{۠�V~0r_`�Y>\`�I�T�'F}1G^�I�K w��V��j�*L�#��#�wq
��Ӹ6���AۦfI���	D\��i���<���b80��֯�$��N�Ʈwj�	?�5�Do���RP��?��/������>����`���a� �f�gUXvH�`����YF\�wNa�*Z3���HC\��������������.A9Q���;�5�c77İ����:ns[���6�_��{�yڈA.�2��#�lS��k�ط�+�H��	:
 kN��4 �=��nЩ6P0J�W�2ễ**!1��
=6Dc�ʽ�|}�1�_�b�0<�Uϟ���{�U�P�uF�d_Gv�/x�?3cw�w�tj�R޿���{� �����ʢ�Wʄ8WPs����R<O�	(�7�� XÜђf�ļ@�ż���y����/k|�x8���.�*[�֕��.�{xW�>ߋmŅ騯5���X��N6(m���6����:�Zђf�S�G���û0�Q�p��*d(r�Ru��3e;e�1�^�vy�M�e��5��'(��8�mΒ��E�k�l=��<Ͻ�Y��<���>9�{<���|����:1��6]�<�ج+���
��أ����Bw7@�m�xrF�����v�+�ؑuY���s�A?["��˧%��t��a!�QgQ�w��,h�Svn��蓋�j�峢�50�I���B>֯����C�HϜ������'��|Dkܯ3�*Eo��!�.T�ƿ /p7��窙XW��<�M/zzy����Ȼ[N�VqN����!_i6��,�De�Q���<�	q�9>>(jDh�yG8[��$h�[|H_�J�����=����V��_;=�M+T�(��If�����wIru �������[����8�r���`=�2uw��َ�����Z�)���6{������A�q�*�I�t ��tR'k�ӣv��Ņ�|���x��a�K7��8h�X�D�f
+T(��r��:���R�C�!p���5L���u�׼a��Ee��<=�\>fH#iZ��6��A�uy0�,�iw�&�:/������,�M�.�В�{����@�P_e��Gb�X��R�i��y�碵��]*�8��Hb�*Q�9���Z��-�`?���>�GQ����І�O�=
��[%ϟ#೷8�_�]�f� ؏��nYR��k���W�M���ad��M]oT��t�a?D�!gp�[O�[^�C�B��^[#ź-ԇ������w���W9���#��+������ H��2\`P<��m�	<PWӲO���ԏV����a�=J&�[� )��d�b���U	H���vJ���8��0�/\�ɘ��q��.�/,ґ��:��{*�݋Ia�;�$Q��q*$Xg0M���[OgW%k���V�Npu����J$cq^X�ֽ��V����k>9�>���P�eM��.&��(Ã��L!���?&��]�ׂVc1�ih;W؞�J�,�#>̩�N`�߈��2���
�6�ga���fbǟf��pߔ/*�=O}0�(f'��t����J�E)/��(U�x?�F(�KS.A�3�*�U l�<p�� ��������b�`Γ�4ݬ��E|.�?���!OMd�y�0|f�&�<��>j��W��L$N:����'�c�UΎ$lY����-i���xzH�ƭ��8zIxR��sp����S�ʿCO�m�����#������Ijٝ�o�=d]g�����b�)G@�"DH�{�3vU+q��W�Z�EU�"T�R��\��t� ��(�#[R
P��i�����ݕ&��K������_���m��~Չ[�:Z�B<b	�g�:��:>��9�d$�ܯ-L�U�l�ȃ�>�V��MF#�����^�Õ�ʐ�D��vA�Jr/f;

9*L_��B,����y0a��:fͱ��M	�����vG�PPd�)N\�wz$]Y7\���}t���u��ҷ}0�x����o_'��+xO�cVmqo�	�~��xrJhŚ�T�҉��L��v�EV<�6�g5��N �!�t�2�̓S�ȥ��3#��_��1&RIr��En�G �@��&'ϴ�Z;:�S%!��ٕ��}�deX�ˑ�黪J��9k���C����R׹�QC��Б^x� ����8�/��(�Σ�l��OZK�e�u���9 hNϤMdv��XW���WB˄�R+;��wⷶ��du���@��./�R�۸�ߊ&��չ�HQ���=^\�+���.�'A+-���'�B
|�5>UgܽNK�.Qt��@Az�\GnQ��q5F���G�E����(V���9� �9��J��6T�s�s5}j6��Z��1�'ܞ� ���Q��PN|K�
ĥ��p������`+�����ٵ�1��l� ���ꔄbe.�	����ZkE'�ɏ����
�� A<<��.��^vM����ࢦ9�T�����3���HӤ��Qq��Hϙ�&@�:I*i7!K���\FR	j�.@Cx��bR��C�}_x��v�qz��mR=)�SC7�@�E�$e�o�*%���ؿi)�re;U�z���K�$p$Zc�c;�;�>xFwk�:�]��N�2R[χ�u0=�d2O���_[(<0d_)ac�]����۱��Fp�����a
s��f����"Ft�t���ZP���I�/�*�;���k��^���I����8��~�㗏%!�6C�xX��㙯`��v�t˺�9)����kK�Bzܯ.�;��K"�q��ׇ������
�L��]�m�Z�%6�����R��΅��ӹB���ca�F��`Z�.{�\4'�xOo	c��AJ$�]���QW�*x2ޙNռϘF*c8^G��+c�հ%�:*K(�0��:����u�KD`ю���>�N������c�9J��ChT^�hʇ!���Ua��H}	T��S)a$�.źѵa��҇f�˒{�GE^&����EHS�X��L�y�4H�N�Bde���RPM�s6�x�m7f���}�U�C��\�]�%;� �L���M��k�����nh�'	L�4�v�s��-!�4�ѿ\�����;E������;~"g!�Tj�֖�-{mЫ�M!��E :e3O��ԊO��J�=�[�pƦ��ژ�:>�Y�;�:L��'�5�![�?���t���Ԍ����lr�/��Ǹb/
w��}20������������s"~F�#x��������ne��V�c�)Y��m"R�s�5؀	�L�8�$�:-9���]^���?d�&0<(����J][�-����?�j�6�WM���^,Owo��X�
�ʊɂ�S�.��S�wd�>��������;��)�{��eW8��Ғ�WWrq��4����豞�P�>P��s:�e̗G93�7���cQ���'���[X�m!_V,׏��
~V���A�J4�ޫ�(x5����>BP�W�K�/ʾ���0�@��fC��X�֤����>�'�C�*<n�l:]��U�p���2p1����G�	�I�ʃ��}����5F�rp4�+��LݘW�z�?�\{!�}�`+�2�x;�b*"y�6�Nv`8��{�MP�j���h����Hv+�9R1�0X��ƆV��l�Bn��=[�#�fD�jN���^��0"07��E`@oYD�i��F��{/�>t�W���,��0����'y�PR�q�����^b�G�	TH�h@o�����ig�H�� ��G��� *��MY��y��9���!>U<D�0e��zJu����Wob�#	�-�oC,b$]X���p<��Yx�����o���*��T��m>��a�1�`v��n�/X"��RۆwZ!�U��+<bm��k�o�7I��T���j�I��Z�ӤBD��D �-��"�Ipl�_����{�����2�=�.�&}��"�l.\���X%�*od�)�c#SE
#Θ�W�'�j}K�:���e��������y��Q��9Lj��,�����}��c�-�j>��5��v�^W��oi���es��K�oT�4�FB�,�1����"}�4ABÂ	��č��C�iR��m�τ=ŵ��P���Y&zo^]W{qѧ�����4�qVP�{7�|��w����X��XquI���eĝ�!�k�T|�|��\�<�o�����/���cc����3��ivR�ZF<A���_\��Y�e�C��Dm�r})b'D2���e�c��bM1��A�
�|���^wʇeg��ɮC��W;jJ� Edb(�u�D�����҃b��l|��ؠF��ͤ1a�f���R0���>;�c_�y�7ʜ}��s�oe9�%�Bm�}�y���E���7��M��]V�Z)x_V���l�É�x���+�µ�UM���s`��w-����-u�p���8�kܼ�^��8��o�/��m���)�9��PVh��]�UAf*�ϵVS͡%XVU��f;-`}Z�#	�J?�*)ẉ����1��cf���p>�
�^�Ŋ�z�U�����)��Fӻd	�!�to�^���%ה�3R3�$y�V�Y0ۑ��ً�0��\��ܘ)�k�!�������JM&�o��N���T�(���s�g�5t��Of�2�t��w�ʽ��%B�n��p�<�C���>��"�Y�h�~*Rk��¨*����QҨSU�P��m�c�~X�z���$��m���CD������֩"C�C�B��d��a�����WýI�i�ϭ1
��lp֍�G޷B��P�T��\���+���F�=t�y�7&ߎ����<c�f/6n��I�7����sK��R��#��h^��Wh4w�Y�7fJ�ɐ�Qi�$�ɜCBbe}k��tF5�f�Z3���A�����o�kz�7޵����ǯ�Z&D�8A�r�K/�W��XT�����fC-�����n��Ux��o��s��Wm�i��5}J�g���:�I0�y��cY�u�ɫ�o�"gv2 �[m.0�ժ5�-y� �B��QJ!��F�P��j��b2�ǀ��t�D��b��1l��ϔǭ�"'��B��m�����ꃀI��zך��fؐi���#����sE |�27�J�>tJ���i����@���>�5:�,_�z�v6]A��M���s��i��:� �[�s��h�?��Z7����Զd�����6�*�Qy��n�y��%�6_7(˅�}mH�!z�9��$��V]*�eC������۷�'.N[kҬP��&�� `�����TDE�j�v"O�[C��`��t!92Ld�z�
�i�5�U[�87����X���a�C������yG?�D�7lM�Jz/4D�Fg��o����YM!��Cפ͟,��4�ڶ��m̃���!&|H��|G���#8��\�*
:�J��w>
,")g�-��k%9�� C�E�,ny��A���(%@:NҀ�xk�̫��7�7���'���,��� .ޖ�[�8!6\̫q�Њ��"�]X�3��G1�2_��Y�����ɣ}�p�D�c#��D��d�g���+��V<)�S=���d# �����{o8��U�:����w<���(��/"lxfF�oR�PN�A2˒�����lN�"�
R����pr�Q���ӄY��`c;�Ղ�&q¿���R���)5���͇����H�6��h ��u��O]v�g�Vo�,-��lz2ܟ�Ǩ�ݔ����r�]���SFB���qK����# �YH$t�0����ϗ��rֱ��J�K)��7�h�Qi��D�U��%>�3��]^�Z����l4�� 5FrQׅ���@mлz�
a��a��:>a4c�k�Nf'x��gohL�A�r~����ItQ�g`OF����&�Ӣ),`r����=���o�!�+�m��ά�̠�Q
]�g=O;`�[ T?�@�hw�.X3�==��p#��O�d�2K��u˚|���x�G�aD�c�����c8�hDT�BZ_��\�V��� e>_��t�c��'�a5�&�o}����I|t�<�(�)�8�%��i��P��t�Y��%6os�қ��������\�j���80��'5r�C�]y���z(ҁ�z�JzD7���.K���G��NnM�Q�2,6��4�˿t�>����J��	�딪�j��JFQ�ܕP���eOB��,{StK���)silXl�G�X�逬��߲�ׅ�eL�ZR	��wO���P�x/��"�I�x;�n��x��M3��_ϖ����crſm�OS������B�2��7�%c6AQ?���	\��n�B3'�Y�}�!������a �:�l��tù*�C�F�P�cL>e!�K1�����ݼ�˼�B��d�A�Gׯ�'@�)5��P
��t�8�5��j�Ĕi�{|�C:C�*�߇�Tk�,�f�J�e7�3/tO��l�Gp�C���A9Z�0!�E2�k�S�B��Ӈ��t�3آti�+����Q+���Y[n�oN�A�,]�1�"���:z�񦆝NmS=Ž���tY1}��	�%���B
$�DЦF�ɡ�.QJ�zTۜNzZ�	rs�3��m��\��bg�.���:�J��0�M �;^F�1"���Q
.X@ǋqK��i��A�Y�p&o4L�$��J���^�g(��L�݉��[��I4�9AI�75fC	K�c�R<L���:�P[Cىt��\���9K��e���V:*W��l�P�{x�{]�W)z/	��	� e��2Q)\~^��f{��~�e ��hl���V�f�0���Fz�E\W�o�MЧ@����d�u���rE�z��_X���#�*�h�%Ҭ�<��nx::=hҍKn)��i*�<�eʁ��Q3�:E�58$�'���p������R�ު��S=[5X���s�)��8v��b^��Ai���cЁIv#a�w�h#��(>oCGxuf�,��j���P�~ac4�t�|��rox�cQP'4M�e�/Y��q;��s��0�!ר�����^�*m���*�C�������[��O;�3�u#iP�#}���2^t�6���}f��pv�ӭ��+�����Ip��p�q�����Rdos�k\zay�ؙTPA��"CIWJͿ4�"�W�ho@z*��3%��!q�G-ņPJ;MsE� y�ѿ�i|ow��O��v�,�Nl%�_�q;��5E*W��[~K�2b�di� �p��ɂM�1q���f���<8$s��Qm{�-n =Yn��ĳ�ph;���
 �����,�t�oX�pr�>����[�tJ+(��Z9e�U�Q�#8�;�E�L�>��
��d��5w�,���Ш�r�]G�Q�N��?UM�t�Z2�B^x�g�eP�ql�A�����L{��
�7>�t!�(o���}�F�Ao�]5_H���FP�2���ۉ�⮍T*|��ُ\b#PӒ���fB�ۢ��t�Գ����vP�Fg�]�c6V&��޴��NbA/�iO�}��]h~q�Lx��P�N@�A��ߡg�
��8����Q+��5����6��=_��q'��D=�%�����n��7-�̥�ģq�BVSS���&��0䙰�t;:{%�I�h�:�Ϸ*��W'R|�`=�L��6=�Gt78v"��Ƞ�-�3��ɑWT\�a�oE��z�"�a�Ī��{�2M��7���\�Ćk�<��a���y�v�O��<|�vfՄ�he�?E�-�������Cto "�I7z����p���=F���DZn:,�=c�!(���:jv@	�_�^� �b|����Yt7b��R�@N��uVK�}��L�,
�i������{*���D��!i%1h�7�}��s�F��{�9��|��+0�Y�t��7G��6D�\ܵ3?�o3��������<!p�!�g	��0Re�Ĭ�y���%��r�a�+^�+���{�W�}��euF)Y�K,�fM �uekﶔd��