��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8«k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7�vG	.� ,�=�K��6o3э8{'q��''��}��%��6`tٮ�b�C��?8f�Vn����t {ZLp����b$�EИ��<h�~�"���d�����7���j&7���������N�#��O�yh� �fB�jy>�6�0"�lP���7���V����`�ʻ�2�Gɸ�*�H��{qQ|�J=V�NC���2�e�pV�<R�-R��;�����ۯ�t\�Z]NZ=->�_�}��y4ڬO�6C�6���m�e���`�k�ʏ�V�+��>ek��k�ˁ�]����Ӱ�k���Cs�ޅ.���#)Y�.�\GH&j�ʳ�!�[��P�;����m���T��5zΟ���ק�Ԕ���*�,�w#����l�e��/����"�|�7���q~L�|(zF���Ы�:��p�Ɵ��M��1ܨ�&�-8��J������M)�=�8��GED���_���+6���h��Y�ʻ�t�Y#�<��M��
�&L�56������!e��C�a���޿�N&�لy�>3���x���Q-hW���f;͌��Y��zu��˩C�L]��WnGD���뙏����P���m�c3��=Ǌ����O�'J[�R�Z�ZM^���cR�16;�y�ϖ#�B��_Y���$�6AҠ@�!�k���;M�	��u�K�i��U����z_�4tz��[��q7L��e)�'��F��x�H���S���l!S�>G���::4!�-ؕrM2,�wX�cE�|n��:����@�t����d/�Q�	��M����%�
��~�#7��ɿ�' �o�gl�գpǎ���7� �h��B&Y"uZ�³~�)����(�1��;�ӚS�i�I���+\�8�( X��?����+�[dg�ˡ5/�˖h���<���J>�����v��V0s�x��]Z���j<��/�:j�ܤ��	���U$�:Q:��ET&��+@�a7�!��KDl����Pd���;3��kM�1'�\ĞM�'�/��ji`)��D�1�]hX�j�S���g�vj.�!}ii�>ʡ2!�~�º΋ԍ��o|��t��l�]
j�^������z��s��h�m]����{�i�^BQ�\^��U=I�.��3`�� ��#f9���v�ܪH�xS�D�YtS��'�d~kP�͉���9�󣿠9�~4O9��Rϋ>;>50/[�,�R��-T�I5
�M�n�v�˚���W|�6O���n[�jM�l�3SrR練Щ���αt���x�am?��z)W�B��,��_A�$검�f�$pDl���]����՘�j�F�#�4�1;�R��h\��*�^0��2񇒁b�sbQw͆�U9s��-�5N�ڂd�&�� -�YD�Kq���[u�nX��/i싫@B��P�(��x��9���H�\�T�j7	{��s����Q�K��Ӹ�^��.��5`i�F��HpLϱ���?H������:n�x�ܗY~A��X��F��=x�PM_��R�,�P+��s�G�0�C'����(������"�V�����=í<+%p�+�T�A������ ������]-�/Ȟb(����}��*�J�	���t9}�}i�L]H��gLJe�:���}-j�p�J�w뻑�=~,lx����^kw����g%��q+�<��������)fJ�x�S���&{��đtyS���e�c�U�&<ֽO�tSs(	�����P�D3������Y�mST�yp�P�4fd.}�y-��΋#�a�6Z�<U�R��>8w��3��v6��6�j������0m{82��JB;ז��о[a恵MY4E���jt�N
���L�/W��}nT���p�o �_�͜�|4в`w`'FT�1�y�� ���6Kbb�V�M2*d�刷������a�*���~4����LݷY~���_�j�53/��������):E��~��0
x���N�F���Af���M�O8�y��s��-�b(�-����MM���i��3)}*����d�Ѿ�b�x"��^1}D�C,-����1��rߊ����$߄���Jg��p�z9T��R�*=�����Z�P�H��T��Bs��h�f
�8�u�+!���ްT�E�/E]��/�����ļ�\V���0r�/yd)a�1�ؖ�ӈ��K��h��E���E�M�h
�ks[	1S��M��YR���Lp�}�j��4�6:	>�>A��;wgG�zd=Y��;�9e����XU`5W
��7]7��^��t �Mp�R��6�����Q�q�|�c���:o��V�4ܠ��ȶg�K���V�uں!�_�1��ZO(��1�0���RZr��	��^�SO�)Ե�����@"��X,ȗd�P��'�R)��"���OR��?6�H;Gm`��DXq�%���ێ�xO���NM�N򉀱�O{��ߚ��^�\m��2��Q$��	f@�u k6�&k�+����v�qkPE���ٽ �3� :}-��M߫�VƳn�Vyl�-4�߱�K��d��ͭ�"�O���np��F+I ��q�tZˡ�յ�X�e������q�|,�#�jxA)=	���Ic�hE�� ��E���|cY�"�+|��q6r��t������B�_�P�F
"��+�٦�$؏�ʐnƛ�VQ��e�/P@;$3�'���4���j�+����н�s�I�4̉�c���8Q�q��;�5a���z�Y����B�;�Q��!���j�d%8ڨ�qE��'�n,�Y)�
U��xQ�\�"�Тdּ����W����O_'ʛ@�cb^%M�\�|%^J]�C�D�����q$��ZH2���9��d#�����\�rp�X��S��W��bV����;�5w7���&槷#�Lg��.��!϶I�G�%[������;��R+^D�|xO0��+b)����Q5��ώ,rѢ'���		c&R����1h\�9�-�t�'����BY}tpe!K���τ�"ݸC�|[~zu��Y�g3�w�&t��
7� 6,X[@�-F���^1͆�$��h���T�Ռ�A �]a�������]4��P��u�fϞ�� �Ku�(Ik���H~�r8g��z����dڝs��"�،-^��nt��2��.��&QЍ�
ܩ���ջ�+>=��q�5W	�fX�X+0Cy�ހ��G�ͻ�w��K'�1���ɫjeƾ�PX]7�}�P- Z����Z��L�9��"��_���~�rO�㐳����헕�w����\1���p�s����w.?���6y�oV^O������K&9�8Jŋ��)W�?��b)(��� �5�	aH���_L��8{)C�)��!�̃��mr�%��h˖?�K��sr�F�ǃ��j���� ���i��u���El�'9|Qgd�YYgSYc�����@#?���F>���ނ`p��1?� �jO�1������\��H�ʖ���m��m]�Z.(�y�}��Xj��{c��Զ �g�|e�X)҉���s:�d宕��(7�-^\���!�w��%�r�qX&��Q0�Hv��4�)�;��q� ��ٛ�F������W�Թ�t��C�y�tM��ܽz�p�ϕ�m�q�}ı�?xDW�v�xY\Y���q�=�54������<|��������?���,�	*6)��XY�s�|��%���kC�{�|��P5�.�ю$��?.�M�9|
������1�,dM�Ɔ<(8$��hb�읓o�;�$���<�������;��	6V���B욗��e
�%�9jA���\:J:�}6�D����ʠ����D�7�t*��141�&��m"�nFbrDGY���oo j�$����e����2�Bj�<��p��yq��k�x�j��Pi��á�� ��ʉ��6�j�?�m~����)�ā�e#A���k��
狎.7�.̔�B�]x�>~�Ȟ$�u���3V�B���eKܱ� !�H�d�TcXjRid^�K������"�=ϵ擞� (T�O}�~l�۠��H��%I� ���'oQ��=Y�a=��L荇fO��{Ҥ�I�C�n1��O[5�p#���J)oÝ�.�D�ek��
���S��7�e�2��
����Ϝ����d��� l ��T������q��y�M'c�qOY��=�N�����������$|��@s(bڝH���oG��$�#i�?��}@h��D��h���!��}������)D��{0����
i	���pHߪ�h��-}ٟ��Hq�#�J�k��O*�E�+d�x�����+-=2�H��e�p�`���EA��9l4I%���D��N R�ʋ�P�4���?EqO�}v�v�B� gJ�~�cc�绥,�0���ٶV�����L@��ٹp0%m)9�7]?[+�͝����A��e���j,v������0���}�wNB�=b�C��/�x3t�xTH�֎pX�MmF��3�6�׮{�a+�erӕ۟�{d�����K��9ѱ����߰}���PAHU�;�̛r!�Ǡ�W��h��xXh�	N���i�l ��Z2�ҕ