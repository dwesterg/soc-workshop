��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8¢�}E0�Ķ��V@�~y�x�1M.�=���}�g�.(���T��O�6��<(&{�;a��=Z�����h6}��w6,��F�="W�l�r�L�lCU�|�`�v����y�6�7�xV��^,��^y���љ.��\� �����Q�����1`���!Y'���m"�.�JBFxSW������e'�����Si��'7�� �7������mrԳmM�̨��yĕ���L�6S��RO�l��)WV\߷�1a�MDL�	5��✭�	������ʗ���G;D3�����?~�OK�b��q��qؽv}�9^O�;~T��rH�9\1V�ī��5�]�ga)�<��.��p�H��1�я2Z�]+��CD��Ϲ�Q��a�G �iQ 2(ğԑ���#��.Vo�M-6!��!�-�V�o�w�dvat,Z.�sp�)�̰ Si^�����l̜mg,��b�Z�)��k<��檲��L���w��s�n�S{�K������x�:!��'���>���d��l��-��y�u/��av㈗���/�c�O��;8S9�r�[���+Q���,."�-�����m����F��q1<�x�φ^Bs�B��ˁ2"�H� �s���1r��F�DL�N�0�}k�`z�}�4�'��OȤ!`s9a��O�T�q^]�m�Y���'�>�F�ǰQe���>�	�X���E%��� &U��Μݗ�`��7zgF�{�v�Vo�78y5<�($��7�Al��R���ʹ��.��3�hSKc��O�]�H�����o�"�`Ћj�ÚVkG��R�&���A��o��M�/Cv����?oǁM��oe���A ��l~���<O�O������).L��s����� ~�����pz�{�\�:�[f �o
=:t��i�O7�+�a�5�P�,��aJ����q���:��24�%�XJ�����ά���XY��š��@v��&r��Uv��M�f�m��VCh�?�}�Ux��+S"k��n(v�99�����L�6r�:a�:����J��`���pH^��F�k�Z-����$IN�T��-}��W���&c���c؎�{0O��0�D���L��.Uդ[�,
�������j��H�X&�"#�vrW�������.>Y�C���L�wVu5�:��KZ�8��jL�C�	�K���L�� �BK0"��՟K�=,;���i"��g��vm;D�t¤�~���Gu�`/8�i ���WۖkDp�1ڠO�_0�`]+B�	�Yi�jO^f�@��_|S�o���0��*���:�Bcɪޭ����H��p���,MJ|�1Z��� iQi��7y�t��i��-<�y3뮧���y�6�&]��%.sJс֕���-�f��~�	!�g�o�M���V���^�d�T6��^�s�v�_>�d�_��#2$�]����g�q)V�O@��x2å���tw�Af�X��q�U�u�t������R��e��!��S�8��m�+� <a�
�������!�$F�S6��w�7�vIv���m����ߟ���w�m�=Ê�!u�Ln�9�m$�e?�[Y�xS����3P8�	�L�,��m"�� ���T�.�JL�5H�g;�a�h��7�o<Qx�^x.h�7��д���B6<<����,=/j��}:��dT-��l��$KE&�ڗĔ��|Zt|�z���z@fͺ��(�Н���F���)�� . �$k�)�ْ2�.'�}��~PnE�q���M������U�V�C0��C�0{3{S<sp�u�F�N09ߕ&u}fB�#�R׳���e���7�z�jGDd�5�9y�2s8J��d����"�ʹ��j|��?�t�q�ItÇ���(4�ak����IﭙL��P���)&h:ۋ��r'���v/����sձM��ӄ�z�b#a
��h��mŤ���oh�%N Jr�9�Ab���52����V:�15�~B%Ej���tEݞ�Wx��4��j��+�:�'G3y��d+9�� �wrz�+�f��s��4� �`����FswV#��]_�O��6P��Æ(��t"ͦV�=Y��̫�ۦ'��C}�� D�xr�(eC]q�8h��?�Td��(�9���t���e�C���:Kw��ϐT��N��N��&�}s����Q����Z�]~N"�Pz!�`$]�~9E�確�����M��w��	~�F{S"Wzk��ْS��sL�=���1��4Pd���:�X�����~�#���ɵ,�0 ����O�zkG47� ][���}�y��eL&S)�o�2�aHy�.�MFl���L���	�����N��蕧�o�|���j�d�2��~ꛑ+;��>0��ϟC��m�"�y�#����A�*�ú��/!l�# �(T*�w Im�B����C`�՟�A7zK�ZC�O��1������?L�@�����O6�
"x��� H8�H���o,.��'%��6xW��x�XW��ј�woaH��L[��A��Ce+����9D��)'j`7�k���"�k����?D`�a`��������/�8P��/W���AYE���&�5�O���k��x��3!�P����U�JH�v�M�O�w~6�4��m3�:�y��LF�_�+�-��$�k7�7Y��] PI&P�c$~���-�V�
��L��X�F���3,�RTF�cjx���b}���F���	Јe\�]��V����a.k�m�eaw��nJ���ḏ��u:�@4���.F�w���O����4�F���3r�4�yZ��_��po>H �.{�x��5q�]�k�����)�=0u�@�Y���R�����xy2�<M߶<ud�~�>��Xy�=K2x�Ɲ�l�G�j��q9�{6#D���]dj˰V�l����6yx�\��͕�ܒo��</��X*�K`G�`qy+B����/>87���V�y}��9���O�{g�$���" $3�ҕ�ƙ�Gl6��pm���޲�����XFĤE<c�r�jw��#�;+e���,Y��+O��`��'On�C�YJL+�C��N����m