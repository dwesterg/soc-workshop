��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd���4	IV3 i�^�&3Ts��P���=�/*;�bʑ0`U���bB�@��dy.�f�-PC�:�u6��YP�9��w<`�=��B�;-�Dp�Wr��e�E��&���h���������r2$�|��G���cw,��B�
~�+�U����I�.��ǅV�.O�e9�� �Dh�;F��b$��F)4<�/��O�b��&����y}�׽G���nh�*@�{c�e4�R�R)��LnC"��y*~�ad��*R?��u:;��^.= �ӶV�v9G�c��R�c�}���4F�S�`����}eN-v�R�R�t�C��s4�q0�^
F˯Kz�KR]Y�x��?<l��Xm����2B��� �J�����?4RI�J������0���\�B�[^B�g��˴N�B�͞�U�mI|NP�R����#�rdu�� ��
��E߷ÏW&6���6���:~xM]�@3S��m[�.���qn��xd��+���C'�;͒o�1�����+�ע�S�N!s��D��:^�Q�2���b���Ԅ�,ٷ�?�֣OX��2�./Cs�P���l�`M�0Z�d|#2�XՃ%o����qX�09��J
��'�[���S_(lA�����Y��9�E^0	&?��3� t��.�Jѐ��Ρ������:�~�����r,o[���7��w$���n����l��Zf�m-2����h�u)+��z����k��Ei���E6��кHLo�Qr�f�؆s��
�2����8��ʚT_�^���=쮳���O�%�$Ͳ��͐i��X�)�
�s�'W�˵�y:�p���J!ё\my@�͓���I=:U@��m]��%��`�fs������Nz�~[]�@������+�N���Y�*�ˍ����Q�C��9��1��Z�j��g��h����=b�F@���ެ'N�g3&����]r͆�BTl���LYWF3�Vx�/1
W�r��gyg��� ��N�%6�����O�[���ș��@��mR�%���ߜ;
�H����,:i��������)�%�ƸNm=li�ڠ��m �>�t��p����VΫ�dL?x>� ����o�!��G���Q�X�o�m��_&8��XTF,�"�n`W������y�S7�~?wl	��U�6����p�s.�m^����o�sk�,et�<��U����y�ns{��w���^��8HBC1A"���P��wn���d͎F��`�K��O,�cjݹn%��Yya�X��Jy�N�����z��/�A5����=��s��%����`�sļy�қ�j��$�宇���j {�Šv�Tp�W6Hl���\�>>|b�ѻokCpzӢ�&�5�^�6ͩ'��ôo�]Tv_��̚�aM+������qu��\�N6̉��Y��H\�A���Z�ʅE;��ӳ������-t�%y�5�S�F�b�����t�.*��ڞ��.d��}���-�L%���zd��ӭ�ޙ�t�tH"�MY[X�C�a>�u��c�C�Pq)&[�c�����{����
	�8i��Ρ[�<��"���0��=26���BPG9^O���M�V������p%������&�Pq��PR�;:3�.�s��"U;2V�g��4�(܃@��G$p~��)�T��%Y#����]��R�Z�)A�48bf����7�5�D~���嶻��l�Kff�O��(7�1
E\?Y��/�����a&�~�&�<���{���<�;v��ɛ��*����M��Ϣl�:eN�Bg"�26f�%����>�_V�W�95D�g荃�j�0�c���І�4�<r]oP���6�~Q�?�s��x�2UP-��\��+��d�N7L}˿��kJ����<��C��'�^	b[�