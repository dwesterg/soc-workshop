��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t��-Ok��S��Xr^�
#ƜaE� �����&�f���8��K�+;y5�n�ޕ,/��˃P�.D�>�6�»�ݬ�lnUK�Aq��)u"C2k%��u1����G�IB_��9�S����<�7�OnH	�A禠6U8E)�uDRV�^K����k���"���e�G]����*�0d��!"�)$mm;|�ZWM��{�µ$�ll?���]�P��p�LV�U������±���8x���oL�hB��#@m.�>WK�.�&L;���K��cS�5m�Z~�zR��{<�.j��uGs����bhv��s�-�ϊO�B���fs������K$���u铦��X�zs
S�Y����d͑��p��]w���s���A0$Z�?ڙ�竾-e9�;� �B�w���tM�$f�x���q�gke���ySh<&@�o���v�~������  �@�8�EQN��͏2Zr�eף'��&>���y�r�W�USd_��q���%䥓�����ܛ��#�:	Wd�~0N�9�v��':�_z�b܆�~GF��*�˙��V��V*���=��5S!ev��R�m�id��4�ө窼�E�-b�����"���(��艞P�I�/����N�=��_��Bx#܂l���O����J�{V����\y�<b�[��+f��M�>�z4"�Lw%�iUߠ0a,���PP�,��/\��,���yG/�L��������7���9l5���_��n�����M����;���;��Byֹ7��",UI�=m��)�6�E�ki�����uR@���jK��5lX��ke.ه�X"bޛ-@�N#	q?Ղ!m����S<P��*��-A�dP�~���?f���t/�E���>��6�noHeL-E˶w/V=��CZ���t'��kx�@�.8̃� ^�'�=���J�aq5x46'�(�hI��Cv�(��[�@7��[0�x}��\`Q�&cm�B2��9�|~+^���/2�SO��:38��x�D������US��nP�M�%77���g�؄���/*�W��� \w�:�)���+'U@@vg��Ar�DC1�~ۖ��k{1�a0���şKsJB�	h�'`�	��uU��\N�g�M*]��BF�f���X,T��wZy>7ҁ]�~����[����bjn�q)R���x�`��o:����1ՃzK�XY�t�Gܸ��xsX��ղ��aS�%I�Z�}��ʓR�'��@ʋ�b��Ź�t�^��ʩ�!mM���Rk4)&9����=�yGf�!V���=�P��s����ך3�Er��R���a��_�����њb��G*������yU�5���G		S��ӂh��~�{�<��E�+'��u"�Ih|����]�)H��j�G�Lz��}���<V���v��_U(�I��w3�?r��6���jl�����1�J+u	�Qw�d�L0� ��<+���-��T��ٖǪ<7n�vK��cN�7·���.�i�z���D^TQ�x�G�I�;��u�.�z�)�'.��l�,K0Mh7ߤf�ڝs7����ͧ�+U����SP�B`�J�D�g��vۃ.�g�����J{���f^����D����gL�7�b�ћv�킌�9���Vy���zw�WrA�β(��Qs����ws=���Or]f&tF�ͥF��X�4�#Э3����B?����H�1t�;�iIM/V�${�E
���T��L�F��Ұ�ߋGA��/��H|������?�$�S�B���P��a�����&v���R�.�E�[W�]��|�]��%J)U�AS�)�zZ�>��D�@��] Q�m�R�,V�kA;Z~�O�@�5@|d`���	+h���&�%ǉ�u��}����rTZn�bsWW,�Em��Y�����
��*��t�g1š�S��~/g��߸�c�c?�Vn�;��=k�{&@z�EB���#ĕ��ګ�P�CCl�$� ��%Y�����ג���	lv;hǷ^���p����;�Z�zp�jgo�����J���7)6r"�M_{;S���0��R5�~����وlb:^>�3c4C��VA�D����ăڙ�w���g�"F�� ��[�P��-���-2����]2�#˵f2�I��݂���Y�R'�pJ�k�_��kq5��0qm�D��7}�8�U����{�0̕TV�X��­�O��܆���> ��C�tqQ(�ι>�O��R��[�4��}N��K}#n�`;ff�i,�gG�Jp��q����)w�խ"�1v��a{"[b�G�
$M�%�3+B����C�2��%`��}Z�i�%1���Dc��;�N"��=��I T���&{�%��S]	�`���ե'W����)��OK��2_�:k��F������sTQ�>=�U��16H>Z�A�0A�j5l�� )�6',�K���@pt"1w��we��!2�d��g�e�%�=p�P^݉z�;F]05,>9P#ǚ7�Cc}����8�V���;������`���<7�D��iK�]����I,(��xօ��ĉN���(�Y��=-�r�j�?�z0�+��"����i�^'��rw���i,@\���̅�U����&dx��j;����(Qh�"%0\疩�2�5�����s�tѷ�bw!����Xק��\H��l�IWv�������U-�}F
.�=��Md;���#�#�Ky~`������s��0��
FZ>1]�.r�D�U�l���F�� �A~�S�D��-
0 �����R7�Һ��|>QZW,�^=RQ�7^K��?��C��	�
�����b��ƈ��:�Q�5���*Թ_���F�-�S��?������DoF���~�]�]X��V��S@�B�ʙ� v6/����k���@a���q-�&>F�t,\��z��ԋ��ij"d�bh��`8�˕����$����dMNE�W���-�������w�BV�)�W��#"�)*y������nV�҃Oy�'���'W
��U^$+���A��sޞ>3�1"�$I���*��D��m��IRΜHl�Ex�1%�c���t�9�Q��#J�����Qd�Z?Y������FP��x��(���E��d^�k��8�u��}Pҵ�>[�]Le�b{� �b�Zy�|��c8t����Ϊ��sB<�"��ϹN	N��dÍY�.���޵Ĉ��-�jw��a8;���;�!��X�b=��`�l�Gۑ����l�G�x�,嘷s�q�\B�+�K63�_���oVU�r���
O.�?��7�Q��n0��Z�N�6�Y�l���:�]�FāC	��^9�E���(н�U>z���E��/b�T>�DS_b/Yu�G�����n�[[��;n��#�X�v9�8����L����`�$�U/�we#H�j�Ѫ��� b'z>2:����ds?g)���V�<�|�}�a�(�^ �r(]������*�%�c�B"WR �/�Rs�ѕ=f��7�p*>�{�a�B�B��1�Ev�u ��\�}��!e>R�Q� U��sn<�6�>����讍����.�0�	,�~�7T����Ć���o.I��x�{�B*p��'L�RW��>n���q�+���'I1��D�./[89����ݔ��t��Q�<��y:P��}d�˴(��. �VL6W��JO�6ד��t��+(�-��g���`�S3�N�n��VZ�?�����6CJ���u��ѭȱe��Ӝc��i���:�A#��|!֣=y��p57�VaPY�[����ȃ�'p������Ǧ��1j`{j�aHn�]yj

�Uk
l ]	V�5 c�R�>�ɐP��nvk}�� �CfxVW��G٠��aY��ً)��/a�pO%n�b�U��ʇ����:�Yg��S��P�j���(��x%�b�;�-负�j�*:��IQʌ� -$	�v�T�%�>�#�
�t� ��l���V��������Cd���ۭ0��C�M�� 1����A�K�f*����t���a6�|�s�������R�jc��U��Y�@�7i�K�ȱlf��7k�O�����C3�����_�)��H #]!HY"how1��n
v�	,<��JS��l�]�ֆp��y����� m~��n���n%�5��`UĮ��٣!B>�/��>l;'�h���w�S��u�G%>����p`���4C-�R���^�Q�����bB>e����b"�ӏ�,G��.ִ�+K�3�=�9�Y���4��K�C�D6�U�1_"A=5G3P��i�f0Cc�+qqC���5�G�j[}�^�"M�;��Q�9��]G�-E�a�=�NY��6�1�@E\�l�:��P\�������S�ܧ�:�8ɚ7��(���X=�ҳ�Po��K�e>^3w�*�y�zeVE���ºF���<A��[�^�D-�jl-,{���G�<�w��X�מ�r�mK ˥K��ŭ,�;�#��;� ���	�8H���%��0�;Z��;;~�:D���]�l��c��U���rlA����ӓP���l7�RɞiY<���
3B	ќҜ��a���m�K���3뮽c:^�9`T/ c�s���:�tm�!>y&���3�#�Z�����ƓGG����Ur��b|@�6��R	��:�� |k �,�uhn*��J�z�3��V��g�4��P˛U�gP��lʊ�T�*H��`���a2+Y	9�g-��#�P�J"A����6�4�Dꆪ�҈��v�VY�*����I��Y��L8A�ּvb� �`��7�I�y��싖��Tz��D���'|��O���* M�ca�S�7���~������Y�m����o�B�E������{���,��+���%��N6��3]�|����X�ž���E7$��-�U�1�x�M�SK�G�j}��hq�;��y�˞���t���ٱԩ5+>-��ZtTD�v��LjI{ͯ#^(�p��ј�(
,�ɥ�S*B3�+v]�	�:���"�#j�����[Z ��3�=Հ8�h�4�u�-����9���X�61*����G�<k2߽�������#O��K�n`��%�@����Z'��ZЭzh,I�����A�{/�_��C-��/�.ſ��@��!���T���&�u����T����T"�^w�f�5*�8�Te�:8�4̕�Y	&t>{s���8P �4Tk�f��I�&��,��� d��s�K�+U�4
�gy��;Z�����^�Pu4��>C? ��>}�d����Ѥ9�6���fo�O4d7�J�1��Sy+)o��j�5J&شN���3�t�#s�� �1P�� '�~b�vv�K�~�
�Ev��nߍ�b��mFF6vcb%��9' ����wĿ�Ŝh](q|�Ӑah��^��_1��+��p�6��6W>\l��Jf����J�ta�����"���*�H��l�>A0<}}�״����{�js���Hг"�큣J��"V��y2�U1;Pb�Wx �$K�`��?��@&��Oe��碝�-&[xX*��>}�8oX"K�P����ϙ$�h¨aq���g&��[
mB���O8��7�ngԗ��'����i�ɟ� |��9��W�WY������XD+�0FI d��'�t &U7K��m�0���r�e�'lr-
J��5���PS���9�+7ru�D�j�����۷crG��V�NN�si7+������Mt�4��k��pl��uJ�o�}���J�мz%(-7�u�f�%[u�J
�j�r��Jj���<Ѻy���'��:
/����k9�HW�����i�_�����!E�7��w�٥���(���~�Q��;���"�m����o�E�ID֐���)9��a(T �y]�)<�t�_���^���k�����o���� ����,'}���E(����&aH9�(��`��/i`���ft~���Ȓ5��V����l1?�b_���
�L�����ຸT��`�7�a!��89�E�9O�
��bJ��	�=萤r��