��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u�7��K��M��E��j �M7@A��Y��L�!{��+u;-�5v�
L�(��bk;��=�	�j��T�ɢo�"*t�Pǩ��h!.���ale�Ѽ��&UI$���r�� �La�	ne90H�kP��˟��;ȅ%f����t�W�U�1���[4٣����d���������	(,ڮ,�6TN��UFQ�q�Y�D�S�1��5�����֋��aL����"�������~�eI�`�R��&���Rդ�sy~��b#��i�C2�������Z��h�J�ȿ�r��RZ��-����	AF������<�eùͺ�� ?�Wi���Y��wAj����@Lӎ���El}����V!9��ڴ�Z���'�2�L�w��N0��@�޶��?dF�g~+J�#�i��H�Ҙ�)���n5_x]�^W����@��g�4Y���C�'
M�tz���\�{���R���S�S���G�����
�)���_��E-J����l�t�;p��J�d� 
R��D"�ָ��tg_	��<�?#��E߿u�_�gv�o�� S�Q��TX�M��\���ͫAf6�>r]JȦ�)d����f�eΗ1��˳TFB\�n6��������.���j]pQ�D�*�����U�ʍf�_	��z����q�9�`����>�#.��	R]���ȉ��^���/��rS�%��f� �U��h�I���=��J��bt���8v2�D�M��:��SQ�煘��P�)"�+���Wׂ�d�f�N�h^ra5�W�x!�}�8�h�QB����A�ǈ���ϳpZ��HN���~L�b8b�L����
C0�9I���nG�F�gn�y�����a"l�o0Ƙ(
V"{��b���A�E�Ş���u`{�����3�u�}�Uk���!���	m�7l�HYI�mͨ��Ƴ����TT�jGXA��s�4i���b�̪�K%����q�_�q��ܚ���G�F�j��t��T��?���]� 9{ȋ�BͮbW@��]_�5�ӹ~cǊ��R<Ǐ�Hb���Y�|�{���ւ��t�Y���3@!G[���P/S��h�������z�+c�t��ޡ�}�	� `SjD�7T��Pn���Ĭ�;��%M����)w�e�B�y�y��$�Ɇ�j�_1����q�@�X�UCA  '�z)�\�(r�M�I��8}PJO�S��݊�x�$��l<�1���{�#��o��,��F��j�@�����1Xx8H�В�ԓ���=�k��/k�:?����YYh�
u�u�w5/#yJ�k:�������e��w��/ґܿK�J&��S����>�쨓���m�@�m�X���)��Z��=H�q�ߠ�L�*�U#�I�o���gu�G� �
�A��3cٷ%�=c�R����t�%�2C����[� *�I-��f���[������ez����%���	��7[�~J&Ry���^�Xchz��~����KY.�5���滯�ءݚ����T�/I>a���g��$nn_4�ԅ�}C)KTʒ��r�_[�<#��OQ����:�\�C��/�#8cN���b��P�H��((1qF������{�=�)���J�� tK|�@N[d��w�������f��#ҷ±w}^2;�f>���#���d���c� ��Kբ��×ݢڍ�����&�¼�^�b.�rHH��������N'��1��)�=����v��z�'���Ȣ�&L�	"�7On���d�������`�\ț�Jkpm���a0�dN/2y �*̺N�w��H{XML2�U4
m�)���Tg
�H���ͼ������N���i�ϊ�4�T}�{#:��`Jވv��q_��A:���
7�֨�*�v�ܦ��_�+(E͓��� �h>�2H�PQN�-i� � �BWu0 ��m%!��Z�^V�`�� g^IZ�V�̟��)�9�HdN��������9�^pXr�p��O�U��5��#���T7�ٜ�T��JM��^����)|xm��B��M��r]�p��,F|ygS�*�+\���5`�|%��;�[Mp1:W��%�O��xT�z+���Kuz*ˋ��'�œ.��Aa��;�#��L,sM�����l�AS�j���<-s�����6��,�Ɠ���򲵺a	��L�:u26�q���/�ԫ�סd+���+K܆��E)�̮����J��D�F\[��j�>�N��O
{J�������t�9��ܸ�~����*��x4J��JV2�������v׶���H�qӮ�(t?��>[��ʕi����%�3w����0΄�9�ޖ9���p]7�FBcC�̑D��--�4���^�;C�5�J�Hǐ�K%X
����]UW��F¢s���я�VC�:�^����^n��"�&���Z�~$���4R�QS@�n
>@l�e�=͂|�-�z����sw?N�j$�ڰ_�x0�w��Q�M�5�\Dޘ_	w+�i&6��&H�#��nJOj���!7�X��HL�F;*e]�jY⑕l�B�ʶ�!�Am,��Y�,J���V��u7�yR�s����#M�5�ބu,��
��:lŵ*���z��\j�,��-R�{\!���v�`d��	�q�K� $���\_�s�Q�Ե�'y�j�W!�E���`����/_A))n���h�����,���o�_8��P��y
oʄN���;a�S���*8̐U��(x�A�Y�u��̘>����[���ܙnn�,+�ˏ&ɉ�>�_��]t�]�q���{y�0f���M"�W���8zeL���8��uC>/�_��9��|����A�Vc��==���T)������T���b��!RO��~v2��r>'aZtF�?�:�Nj�f���*�Qe�]���] |�r2$�?�/ "Fzn�?�q��3��@�^#�T������bX��q�YSs�jO���&6����)qhFdj.Λ��l�W��t������M�Қc����������F�fY�\r���������T0%�$��P;F� }�Rtp������3�DHc�*ݹSq���0��덑F�=��������}��ѫw�O�3;ȩ,��ҍAKB���� �x+� ˰�g�C�t��z�MU��ۜ��BQ�BnV�?i�K^s*���f���1�NL��o��RcF�j�:� ����3����3R�>�J�=Y�s�H�|�]�u�������[;A��h��&��2��Y�`t��oy����*p�w�V[�P%~��6��I2�t�;�V\Nq���W�Qe���𩱦W6�������7= H�?BF��w�fG���?��?�Fl_�0��N)I�