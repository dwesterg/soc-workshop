��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>�3�x��=�����hR����Bj2���A��iV��|]��2La�MK�ߧ�~�'HT>~S��A��_�IB�����FU=��_=μ^l��8�޷N��V���n����/"��׬���%�1��d�m�T����'<�`���VWj��ǐQ��ط��D�q�)���J�Gp�oG׶�1:k�8�S�.-��(Xv�`���K��1�-ӏ������8���e��r �9;�!�Y��$�w�1	��k��v�W��,$�1<!�r�˥j�a�"98��-������^��Q0����5��F&n�\S0у�Z��8�XT�mOh,B��#Ջ���x�/�fo�7�y!��%��2�}�(��)L�vWB/̊���������:�����iT[(�T���.�����U\3O��3�ފ�K�?m���c�g��}8� �6pX�lnj�w�h��5E�sR t����Ċ�5�Ni/L�2oMcH�(P�6K/=�2�MnkY>��L�,���`D\��;��֖�Lޤ.e�^=i,�b�7�C�m��3B�1��b? +|��3,Ҏ�)�-OmY��2��T�޵����J����¤��a���(qQ�D�a[�����F�iF�N��2�.�N���n;�nΐ�B^4�6���aJR�-����0жi�m�2-��a�:ʧNK�
��7�ȡŰ�o�*�t6z���0%a2�q���{6���~Լ쐇�'�(P-�:�_Iމ�7nB�ʁ�2�i�f��3l�#�t7�������W��q�0��@���g������g����JY�=煁X$�7��U����+���`�	��	^��l�u̦ܪzu 2��,c	��8�S�.��V̻3s��5�T7�&{��-͸���1�nCqI^{<��lR�jLH��i��f
��}F9��#�QR���fH�T�B�27K8]���]��*�p���d��������zj1$ܤ^B3~XE|����>�%�iچ� �������7 ��m&��p��y�+u8d��"���8�A���9Rn�h_H-'1B������iޙ�P��a>��%����t����mC9"��T�T����pGeV�����>�wkڛ2` k[F[ �%0� ��)�a8i���z��G�B�8j���W߿"A�i��e3UQK��Cf	"��h����Pĉ>jBM��B"���=�mZ�9x��,^�ީ�N�*� hZ�(�Y�%xt��ݖ����bwD,��)���L˟?������E�|Ur��|�����K�s4w�������vO�f����9/;r(�A�3!վ�N����~�-&�v�ݲIko&�ĩ��RW肥y�>	̷M��9�dÝ�.���+��^R�ف�<T�X�R��wi9�!�CK���*N�p�o��9�s���ʪcLKC-��]�5'��|���P=)�
�t �'�5y��ز��կ��@�M�Uf�)��-�=$���X}�G�OE�Շ�z���������$�/oU�u?V�e���-�M��N0�"��:��s��?��5�; �A��I�O�)~Y0kh�T{��ð�`�S-܏��}�Qj�$��+q�ɕ�F����I�X�	Cre&W`�x��&r���LÚ#�<��I�r,z�yoC>N�(�lVDݻD̯��7kӲ�|����B��k�-~�c��|#N��� n�	���ĉ7�)5���)x���2����Ǯ�����=D	��9s#-v͒>���=@Hm�7u�hj�bs��̻�P�_q�V��J;��>��I˃;6���2���j,{�*�W�k�a5��cG'c�y%u]�{^`�OC�b�/��pa��Ϸrpd�Ű�Ɣ6�gjҢ6R�ş7���oϖ��(ZS$�*0�FeguYFM���>�ہ���)���5�[*\�χ�A��Q��K�a�7{�LZ����KT���i7��oƼ<kN<t��"�W��W��&J�WI�ɔn���n��I�*It�h�\3m��aS��6/G	l�QM�CZ ���n��������VB.����5~����s�)��YV{���ڲ�e��쵣C5EG���e�7��},:k��?4A�f��Ы<<�mP�� 1uŹk��y�ױ ���҂>�5ߪ����↖��E:��(<��Vɥd�wi������FaM���S��mč[-�n����[��54+b��,���Ij0��;�[�g����D�)�SOQ�P�S����P)/)f��{��OO��Wn���jݧ�"8.��|>���_Q��Yɝ��Wcy����%M�����a�蔷����#??�I���w������H�v̾0%�'��v�f6v�k������jZH7���t��ű�v!S��UtY���[uE��Q�er�m�/��S&ijp$R�]u��8��h��v�;�T�.�5+�lh�k��ت]�M�?�"B��.��C��}U�9��'ɞ��hӤ�X��f�}�T7)�9��׆y�/f1���I��s�AU��~�<�DW	����*Z-�����wӜ��
�i�,�劚�k1��� �s���-^x8�l~+����R��-\eЈr%���tA�2���Z�9�����ݏdW���E�!e˛A�gp���!S(���gx�)�T�F5�����:H�z�&��.�^*����x�-�n%������{�5@����������Ǒ;K!dg2-�t�ˊl֝���8<�h�/�
��M�p���e�������Ive~�_�O���wDr�l843W5�l�A�~C��\���1�\eە5�H��@�S