��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t�Ĕ��
K��|��US�LG�zJ��)�|P"�R��d�Z��{!>�*�gx�Z[y��<!2���5���>CmA(��ZWm��5�U\K���Y�ג.��,;;�\)��D�_��zgH�nyev�d[5l <A^�[�J�l����<��w|�S<�궈%�/�dק�+�(��hMF����-��#��4\Nn��_������r�S�o@�>��(Ox<��u>�Xb5���E�.�	�'_�����+K�E��8��IEݑ��M�<!���,V�ա��?�u=���@�-N)7�Xābecf�h�ةCw��a=�ݥ�H���G ��,�N�Yf�O� � B[9���HC���\~�b����¦�{���02~z���͋�S��.m�� G���������f�X�l�#Wd�ld5y�(fB��|ω!�	��XO�dʶ�<�+d�>G��ϐ9���Gb�ma�)(�]:&�ؒ	�W�PR�#`����z+�ESBU�V�/>aι���?�(�*����Sk���l��p8�l�^!yл9$g+B>�ʳ$� d�~+cz�*�`��I]m��=h(7f:��ǅ�d��$�e��٩�^o2	���ɱ���Ifx�Z���^zi�������!�K�p"0*#J>%��St��ܠ�e9GL�J���46�����0zt��b�9]L�{S� �����*#�Z�:�k\q˔E��^ c�%n]��0�<���߿�y/������K�}�/��>%�%���V�Mvx+mG�����8DdO���(�ֺ���vaq�������4e��{�Α�|� �ƻgo����_GK[�@�6�lԈ��&��P��Rdd�!�\f�qICN8f䇦<�뙏a�-��	�pVvU�#��0���|ms�� ��	�3,���B��d	x�qyF�:��2���k�Mp&E.�M���|�JM�"ޞxd�3�m��w�x��[P�+S�����GA���Z�!ҋ� �M��������p��cw��i��W�)�t{��{�q9�sR<Wps���&�`�I_�tfr-�
�=u8K/��@Q۲}B[%�brd����*��c]���3�i��T�
�G�8�7��{E�ͪ5��X2�B6�J�A���r�zФ��\OZ����*���ɝs��p��h*�;��-aõG�۵黕�Ф��T�V��{��Y� 9��H�/B�i�+��7�I6Q	ċ�V����8�#�����Q���f@���\��rb�s����T��sJ֥k%ERy$�e�xDtJ���W�b�=oگ�yv����Jt�Y/����bD_\Z �!K�0U�
_͖�%�	6-��O -�zn�Ӑ�.���H��!��]a� ��fq�Z� 
��dQ���D�p�����P��c��7p�T���[�� =&�%�z��K�KD1S�1z"���6�?)�[��0�D���ysQ��֥�#�;Z�C`Q��-{B8	��$�G:�N=���L:H����9re���C�dob��R�{P���]:�~vD8�p��L:�����q�l�@�o!�..��o ���̲��͚B@���n���JV,��[�X.�-���L ��L�\X����p�������6���<��|J� ��c�zG��{ֲ�B�����3P���j���f��@[V1��cc�����I�����K70-���b�Q���`s6����zU��a�1���.�:8&���"�^j��)B�� ����y���
9�i?HsKnIp\�Ѹ��1��Tv�<��H�����,�@%��+n��;QνC|ɇP'Z�ߨ����8Q]�����@��p=�d1��r,ǵ-�]O|h;t?���7CN{򣀦`ل �ʁ�<"�� ��?���ԜFJ_$���iK/s���mz-M���&�ك��\�Cs�2_2�F'_��ʦ���뇆��⾘RUՀmY�` \VP�P0Y�!�l�	/K$,P&= �Tʬ�PG�=��F3�o�!�dK؟QgU��Ж���)6��R�z���s�j2B�6WC�Iۡ�ߑ�j�B���U�~�E�V�I�r}����Dcm�^ T�,
�|X�F�K0J�H�L�6�OHT�j��7j�2���xM_���A���`�U
d��D�~܍�����V����U�p`�:b^�RoG��=�j�9������a�Ƈ�L�ar-Y�Y~���0�C�ҏ�����y:E��{�B~��TV�M���Ok�2*j���<`>��b�:��B��Z%j��IL���P��ק������t�Vz��ƣ���n/��g��i������c�i4)'<�#~�Xt�~��3z{��{�~ VM~F�q�s�t�����p�_so6�؅ �M����t>�t��w�h\�E���Z �2��CA�-^[�9�\~� +���Y�t�:���D�Q�6��uJr�/+,��2����!�hY��]+%|��֪���%�\2�q��s`� �v��R��m� ��r V�#��˄�-p�B=�%�[o�\>jk� ��p��S(�����>��N� �K�<�bi����X����Ş�߬~��_)#��$WYV�#�Q)Չ����Չ��"�P��o���B�B5bQ�t8=���;f|������u���Ԏ���մ|i3�:�px�_à52`�����@5����� 9O���eq�1,t(�Ci576%}�a��K��̈́���1(�m���_?�#X��Ss�6_
���j���r��)��q��/�{�"�X�x�I��;:ϋqNg��fK_4���9�46�}��S�H�{�hyBu�H�vv��n2�D@�e����A(���%��ע��t��<�X�!�2���F��Mc���e(��c�_�p��`�QC���7��YC��R��r�y�m Sڴ70���Ͳ�)�gţ�,�!6f?� ?u��2|ϕ#�;C��V�a���%�f(����7�%R��$Ȟ=���9l�e���2Q�&��0G
:�P�{�֋���΂�9G�@�%����b�	c:�>g�5��dqc:8&�ؔO�!�6G�y+���\.��4{�Q����`$I�T�BY�Fx����Z��D~�X��6�;��.S3^'�z�J�F�%�%uPm����Z�K�3�n`�r�2���g��Ϻ_m��� ��RFm(YTɫ�n��s��+�JNEn�_�R�Ly�C^l4`���N��g�x�qW��IO~�d��CTn7C^X�zbsoH@i��(I�^3�b�W���U����*�bF{�֊�.u��s�#�=��k�w4	z���Q�����(��`�B�[��=,r��;L��x��!�7�?%��/vo�5O����{5�Xn�a�;�V|�בts��f\�B7��V�A��~��>u����ȋ2"�jH�[K�b2�ŎCC([�M��E�"VQoDIU�/6QXd���D�_�(����J3������V��3�iF��J��{e+��h(%����j��M�]�e�|Z`�|@�V��Ma�Y`����1䉎fc�Љ�g��ƪ�V��}��k]|�o����s�Q�*�i+ܶ��[&��S�.tv�`w2r�+�2DeN�Ԏ���Vۍߡ�C���h6��վ@��6!� �������bK�@;�[(��Vp�����/�`��u��3fz��D��9�vQ^�=M9@[o�Faq�/t7�6H�� �\�Vx��3k���#dٕ>�m���p4n��n��C��:�����{@��������?K�$���V��c��� �h��S����mؿ��i����$0�.ֿ����F˙/'�M)E��hn4Ȅſv>����4��>���v%2b9<]_�ѾʱW�@%e{ev�b&���2�aU�ƌ�`�\��h�f�M
�D��7iM1>��l��՛a,X��VHR~�r�j�#>�Pq�J&+$%ÐC��HB�����k�*(�{ҟ�fWA�✣k�j*���.Jֹs�����+�4��)d;ـ��l����U�Тh���d�İ���X�~m�����:���a�9��HS!��L9�e�غbX��Л�����/��3�d�-v�'���X�!,^_�~g+BԵ��/��{zg�,���MT�����4���ݍ��om,�]�2��^a�#�&�Q��vX-3} �G��ҭ�q�]g��>�����p�`);K�ɔ'6DSo�
	�t�6L�#nzը�O>�p�4ԁ�˜\Gk� ����P^(lC�n�%وD��"#����n�$��0��d�Nk!Ű0 d{�^.$�&���`i���+Ș�1��>8a!ک�X�]�?�a�om��V9�d+���] Q�o����0��q�s��< \s���/K1V2w��{�U;�x �2�����]A����O����A�.��[�;E����|A�O�#��F )T_S�ɷ���iT�!�xԴaQaD�"k���d���V�t���l�q?��ۂ������M�?r. ���«���\jR5�}=����t�ĢmH e7��
źl�`���k�9�6��N0�KEq�ʂ��sS����!�Bꥵ�z��'��#e#j=6�r'���q�S�=�Ⱦm7DE�2,
������TF�g��j��/�~��{cWeq�}��S��8Xw�>PJ�_������ţ�������܈�+�H�^4���?/#@.B�.؎(b�* ����o��?ĝ-�w�i)��ln������]�:n�;-�W�9��H0˃b�;�|�GHj��5�C�%�y�p�|��h�$�YQ�,�z[���x
h�ʇ�E׾[�����w9�'7��u#�d7K
�^@C��1H��=�橨��:&E�
�ڜ�.��J�YRp�	��P���!�/̓!f,𮳗B��d��{���^U���6��/�O`�OӦƤ�
��6)Z���QX�������u��˖T�7?�?��c�n�ŹS"X����E�S�Q�����T���Zў�(����]�!�D���9?ۄ8�L�"���&/����F���|���W�B7��
q��}�3�˥*Vx���G��8��a;bdFyNU`�+����YC=���4��is�� ���0d^o|ws�X5<���Q����t+<U�F>�*��!���C��n|�0�ĺ�`�����zGS[7���J<���Q����_O��8�Q
)}�%��<p���B)��b�(���N6 TU	��E�7�.���Oo_ȏ+�Jh���h�H���C�י����O��J+��";���}������~ے���ȋ���iL����Ҍg�&��ճ#�f�������|a�mIX>�T_�e`�u�TT������{S� ����W��ꁉ���^�9���t�q�kMiHh>�����fz�һ^��gLU�aT�_ ��w�4����â[���):;�<�#�bT��ve\McO�}�z�^[�㭀�j@�~!�Y�Є�#�S"b'7�;��X�a+ǌ�u뒊�T�҇sz�fT��&�08�{���[��C����i,~4J����A�f>��Z�Υ���IxSg����eL��;��AF�USQ ��J������vp,a��O��"7_���槢�y��LWI�B9���=z��	:7K_F󦓖,��O�9<����ćkD�m��?�,)��D�Run��!q>�M�M�%L�~}��}�;İ��'bX�n�}�6a�o����ý?��"�	�z>/�Iܟw�;�r�����]I'�=�s3���f��JB�%uG_j��� @qW��Hj��c�É��z�z���{���T��r�N�� b���1�t|�͟W�ns���N��fi[p�Z�Um�3j}�9EyE�&��� m.7��o�5�R� �z�6`ga��m����Ò�mf�X)�2�j��XmP�I�w<^�;I�}�P��5�����*6&�pj�ϋ�ʺ�/�A��~t�n�ѱj�)1��X�xoL��å-��>׍RY�-fظ���rx�0��{�P>�����<�bV�Q5�Pvo7�y#�)�[	0l<����#�0@��',��ci���V{�W�.U���u��0��6�3C�	=�vk.qC��Y���Z�YZ`fY��^<����[H"�.�v���R���c���3f e�H�G�Mb�l��nE�y1�ǟ˒9����-c%U!��m�o;�<o�+H���刾$��]�ݻa0j٬�S�8p�u���JmL+�M��Wx�1�ߎ�O8{�0"��Ϳ�O�̚!�9�3PbhIC�'b�+�[�1��4T
��A�L�~�	����w���t��i'�1�#��:iV^�.om�s�����h{��^���S���/�G�8�Jy#	L�#U>.��� q1��CV���Y�ΰ�ƠP�'��F�
�����ҁB���j�޶VW_����]�E�ļ�=���9'�1��UL���(]kώ��B۳�)� !��³�aF��B�+#�G,�RkM����c��
���g!�t>0ڝ-�Q T�\�H���c�`석b�8�[a(���j::!$	��$��C.�L�B���9����wWD�F	I������mg�G�&���9��9wB�3nS5�C�f5ˇ�um�^�Ǭ���2.��{���.d�5Z.u<�����!�TZ�D�J�a �Z���c� �5i/�0V�0�p�a�&%�!��SH&�v��$��<n�f�T#V:������N�qꟼ�I�va�G#�� 	�H(u�@j���L�G�N�o���,H~�'A?�ఄJ���!�I�\�bM��*��?����l��s:׀��Ӡo�������j��ÚF9S�+)�Ok��au(`~��wM�$�_�텷2(�Ǔ�?Ѳ��X�`ѻ �b���*���"���<KL�$1ϕ��&�Q�u�F+��f�؞�P���?DZ��F�K�oTf`�\�M����U[�C�3}��)t���l!�7.h���T�p��w��$U#}���S��f�O�}�_%N�@�2�C�����v���M/pUG,�@Y����F\�� �Q����~��\}ݤO�:
�G�5̌���� �T�8��g6˟��&'*ڋ�.�fk�6���V-i��7#�#T����D�h�-ZZ^4N�f����䬙��e��vyR����$��Y.�>N��$yH�� l�S�-�e��%š�@�@CP����H��,# 2�!���� ��JX��� �e}�eA|���;���W��r���~�MB�};�$��M�XX*�ʴɞJ�������>���E�+�Sd�["�1�(�ދ��{��Ѷ�R�*�l�Ծ ΌVK�K���
�W�yc4���wܭ��8��B��:�ؓj�`m�nB�*r	K]/&d� ��g�=�7�Cr�իx#&��Hl.q��gu�84�c^a�I�Dl��;�b�����&r�	�-�Oj}�:�����^)uuVA�<���d*�Ρ�	�=�O\�o r��3�%5i�'P��{+	���֮�~h��f UMs_	�e[���z����~S~��yR�gi��&	�<S�S����Q�F�Ӵ�L;5b�jsj̲z�d1�@�n�&|��ä�.�q����*�25Xj9/�_rR�a{��AH�_����6b��#G02���9��˭/<����ͯ�Q��������ӞdD��v���B������5�BG�5
��B<Ggc��d�(���,� v<�����@C����<uB�E� V/\�#7�����D3���RIR�o�^���ڏY��?ӻ���9mA���A����CP���։B�~J4�a]��N��һ��b� ��q�GCQ�1����Vwe���#�T��g2-�~Z�B�(��R��gmH6|���Zh^�s�p'弍m"��>�ϷP�L��K��i���jv����n*1�"�<��PbHJ!9��B��:=���F é�ˢ�3R��f������d�3V-{&�f�V�p��!$~k4�L]N��= !uPa(���m� $��|j�ʠ�`��d���̀�1=l^�=u���gXH��y)�i��F��:�� |?a6�q)�x�wݏB��"x����M���Y����5�W�Ԛ��D��l�2)�J��6&y��7+vF�L��Pb�����: ����6��Ԕ	�f�3����[���k���T�߷��O�_�����Κ�aee���F*�f��tt�M�L���DRh���N���*�h�V��Ҍ8hq)���R`4�31l�C��JY� ?&�C�� �A�~�Z�6c^��)��^x��DF�n�t�ߎ=��T3v ���SS�$k�同�v��\m����<ŽK�gk)  '7���1YÅ���h��5��h��8D�1���s�5�RQ1��䧹'L�
<���V,쩅��:����������!'��r ?��"��"�͢kp�C�g��~�z�bb꺩�ǡ����+����knt\N�Χ�<�=,�+8;J������hjQf�z���G����ԩ���}7�LK�n��m��]��"N�2#��U�Fk0u�IT:��5MM`�cE����</K�nTآ�$2��q	�iSmj%9B�N}h{\ӝ���{Q05�s!�eX��&0��J�s�B�h/��4�L�X�����j��9�O[W���b6�>�XNg��4X�^�(�y=��q5`s�=�(=���<�����p8��n20�*�x
��[��Jܮ�2����xI���a� ��o��W�|"i�e5��p�����O_�됼W�]�	�K�>�L(mŹ�֫w�W��LbAD�]:�3�.���c�;Lw�! \� '۱�n9��	m�P��38�����k��}��f��U�D����c���,>�=�����S���KS#lFaH5���ƥ�"�IӾw�?��[Sj* �����=��O^~"����⇘/0$�Itr�$s��j4�A=�w<�)T�-ܚ����.�<�Ü� ������5�hV��4;]'8���|R��$����������L��1�Y�0`������	w,�ǒ���b~���ԚݪQB�~V�]1������&�+�BK�)�s�s�ٮE\į�y�#?��4��{ HT+&՗_H>��F�ȮD�xS��IGt��Ҏ�+��xJlY�v�v�;^�� :������%Q '���uo���F��3��} �h��V�L�վ���o�������p��8�
�-��=�1\ț���Lh�V�nY�8%F3�{ꔊPT�	��~�I�<�<�A��O��V���H��ٜ��l�bE��t�^�h��;�=��5nEi�n쒐�)�5S��&N�h�Z��������k������a���,aU�QX>�xI�@��B�\��g����S�|��J�](-�b���>+U[���L�p'��]��T;���@tY�"�Q��::�*�	�n8M��A|?����l�q��`��1��}:�@��Q~�Ka<�� �]]�@L{[}��=t����p��%�<��ϧ�W;zUEhf��w�עK7��.ϩB/N�},�|�hx08ȣ�- ���K�X(�K�L����L�Dԛ������P�M�j"K�̀K��,ea!t��
<&}3!L���,x�.���D}~&� K�Hfs��03���&��g4�l�kl�!�K �+�hǖ=�}�/�"qL�z�Nw��b�%d�����jQ��$a�ȣ ����]���OL�V!2���v�WF��g�+��9��_i��n�?�*����[��X�ԯ�f��������g�R�C��dk�;��%��wU�uJ��i�3�5�S�O4^�����+"��ٜ� ���!^7d�L�X����=�<�������ڷ���.,��a�,�����$y�hڭ��4p%E���ڸ�ǆ��bR��`o@�$�m*.�3�x0�ͮDV��>�o�k�"��N�d�����z�+-�Y���	d��y󤡳����Y�e��76t^��CR��\���`{?��Ss|v\�����❲��,�$:iZܯ�A���Lfm�l�7��,9恨.���i���ޥ� #@R���9,P�I�}���6G���.FG7�n��b�%J�-��iņ~���Z@�-�h壅�-
�m@ˡ���Z)<&LO̞8�X��e���+z�����L���7<�����*�����9s��2Z�3�%t��,|-��"V ��N�X�+�XCЇPg�eKQs������ b��Ja�,�|&F�������+C	;�%�L=�W8L��!�Fwٍj��tr�n^EA����S
9W����վ�CYP�� �P��|3 6k�`������Yt2)����������7���՟5v��D��v�
b
K}�J�W�����l$���a-�%f?J`�[SeA�lJz	���,�F̫[8�`ZW31`��5R�_i�s���M�A��?t��^������9H9��g��4*�p�m�.�2eӮ>)�^t�f�Av~� !ZŮn�t�v��F�~_��2�zG�lp�8�3j���sڟԵ�a&(A���3s�Et���A���CCŒ�%Fgɯ�^������<���թ~�B�[�)����.=.�I��kתc��	)�a���EN�j�ư�s��<�KMO�}��$���[��T��CGf�(��P�Q��佷��,#_7s9뵯���XX �G���~0����Yk����i�	_��X�b�"��j�d��u��Pz��Z�lƇ٨HR��H��.`	�����z]�J�%WaA��N&���%�5���L�j-�Lx�<O�q��3Hb���$�PO��ʴK�4+����ߗ�,�oOg�(��c����>J�׉M{�2�ށ�z�q���`���]�߃*���2�n-9a�q��(�:��	�Rn[th28?�P�ӁKjV�#�D�4PRW�����$�/�@\w�#k���'�YI��/H=�O
�G�n�2;*���!��\�4I�!�ve�{@�6ke��l4����M_�e3N�����6Q5�V���wF�.hr�_,�%0��>'��]�^���+.����N�1;W���t%)j��`��i���l��Vtk'#��ah4 ���#e]|��xy�q��9b��-񒀓�kxQ�X|mlM�,��E�2gl��\M��������-AS��#��p��^>�n�v0�ǁ�!��צɎ ��EC=|�fc'��!�k�j( ����:�4NK%��;=���c�mE�#�J\Y��㖻T椐�T�Q�fJ�����Iƽ�|O�X>	$���eָ������� Ʌ%�txj���G���=V[�$�o��Nm�:ڳ]I~�~��ʓ�I<��}n, �~D����\�ݱm�j.��Yg�h�m��;�l�F^�D�Uk���u`b�$i�<+��3��gs:���I=ԟ���M�=b��E�T3�m�]�Q�	�Uoa�GX���_4�Y�e��Q��/�`"�#?�u'�G.f=��,�JE�z�EQ�����.�:���k�Ïhie�������`䞦�~|3��s�z������8gڛ ��=�6��=�X��D�����'[���u�ŋ�Q]��LT,�[:�j�:��.�K6_X#A�P+Yg=���� �Ζ�G{�üH�ȋ�׌�tk!���Rv_��w�[�g�wZ~\��0�*:a������y&�<�s�����L�`|@�����k���%��ijb�l�.d��zaOMժLɞ�����Xab!��Y����VK�!�L�
R$�O�4
����ȿ��?\@��g�[ڻ-F
P2Y�V�� K�=-�1��;-d���E��hu���d�#�3���[Ri��t��:r�.�`|��cd�?ojN/]7@��G
�c����� }���P���w�Th��4�ūo�(垈����9�S�L������r�f��b��}��p�9��ӟ���Z��Fs�F�Rd% <�O��[��������$�#��4N�F�7������B{Z��8u#�w�ÈK`eq[?N��&5Nx������o@/��#S�����A6&7U���B��K7�+�;�Fx��N(�!~N�?�w�U?zs��Fn:Yf�×��cb�=�NUV�Ds��Y���5m'�|w\�*��]�q��#jA$�YFt���y���oA1?�h $D
�<-���
�C rOzr2��5=��y%��x&��k�X�j.1;y����X\}ҚJ>���;����l���0gpZ������	��X��n��` ���e����X	�r&�&9mg����O����Ί�5�{"ν���>�$�"��*k��l6N�ӳ?`#Ruo�%X�F 5��3>�wP�j��bn�=:T�BQT���1m0-�Mv%m��>$Z(� �DuG�5�N��?ӯqvcV��$��~_z�j��t�8Ce��+��_���;���Rp[0�r�j�1���/�h�7Z,jj�f�n�j%�^�|��ۇ]��|���.�P7���4���P�G	G��J�V#y���{d@?rN���&�Ŗ����Nqr		ep}E'ho�eC; H��wbQP(��n�~�&j���8���Zr��]�2C�M�n���P�s�=P�EL���Ep��C׵�[���FLt<��� �w��ēo�Yu��M�ة��Φ(�*�ZQrK&����5���x����:�l^S�ro��J��1��SF��D���S��N6'������Қ4?w0��$)����Q�T��K��Ć�����2QK�鼔��ρ��裇`����{�����i�_��k�c��~c�k%q)�\`.h�e#�*
%u�>�.?�W_T��8�Gs?����?b�̱�u����[� 9l�1W��Jii~è�E��u����%=�S�XҌf��tQ�������F�E])"����V�_Ht-�TEY#����� �Ux{x�K�Ц�#�W�C�rk3�vZ�C<�	�̼��'��)r�$v����#�^2�d�_9%A\ ���-�����a�3��꾂W�F�8�xP�)�A�>��۲�4��ʳB���)0D�I	���aI���Tw�B��6*�U۲�f�����5W[�m�r����̺��f&a	;i[����*ɻ]���b�j�y��=ϸr����,u���1���Y���vQ�}Bj�[o8�j��80��R{�حpD���X�Q��*�b�����Z@P��T�!6��q��E����BVD��*�	����H�˨Qԑʅ�#�1�)�ie>v8�|���e��e�熠��@m2'1 ��k��� �=���������4K�G�<X� ��|����^��wz O��. �Cx�y�.6
�N�dx�8*}��>iw/�Z�=����k�2ctx���n�v��$	q�R��\�}Ӿsv;%f�iT̌�I1f�
�G�e='��
?���b�[��X�W���C�f�
\ �
��-�Re<u���f�\��<�r����-2�����fyaw�����^�����n"���gӱ;����fy,}W�h���]��(G���b5���\�Rf�ߏ��
�B�Q���4Y��D=��j=n����fRER����T�M9Hs@R-�������w���w^=�̉xa��~�Q��r��Եr��W���BR8l��wf���Bx�����ڄz�,%�I-��F�U�Ѓ%�R��q�x��D�`�ֲ�#MX�X��`�����_����\�O�LtJ��y
�d$K����K9_~�X�\�Jr��{h��}�J�*\���)@:�5W9V��X�KBjc��7Id�?�`ڣʸR���;][�4'�I>n�����e�cz�t�`%,��+�J��?fsz;���?(�W���N�'�!{#��]w�t�gm�=b� H�� ����TjRk�~�L�n��,�`ef"�=	�Q�oL���ps�*�A�������|맇N��_\b�\s���4{�/j��i�m�o��zO<p��G|�f�$��I�-�3��I��~�����
�O�׈���#v$�f�r�h��`�'�����G�l�k� �?(!��r~)��:�D;��Jeh�����Vz�j!)�1(s������d���x�IM������.����8S����%NO�oR��Y� ^z���C����쨒cm?�dG����Bϲ�f9!0�B���l-XK��ا����燜��� L(9rh�B���A8��(�FMfBƎ$M���7��q�Q�ݧsD��$|.Z���@�׺�D<�^W��6��%���܆3�(�����8M�կ��J�x0��Nb>nǒ���T���΂����YxT�{h�47'o8I��Q"�|%���q*L�yf-B�g�S��tMA/�|MU�)S]��G�y�::.͑�������sV��护������6	=U��0�_}&�<]�ah�yFU !�-�������Q��2w���<�A�4tB1d#D��S��$Y�Q��Mp` ��xCפ���Y����-1�B`�i&M��taz��Ng�����Ѫ�m3���##r"rE��*���A�\�4�ohoT�7�+c\`G��?Y`-m��zS>�,'�C%ѳ��V���Q�ڨ���Q�՚�g`���Ʊ�a��)CRH��2���N��׀n�.*�I����܈N��t1�ĵ7|?Ϣ�Z*�v�-��a�>��lh���{#���A��2
��<�1?��]�?������OHN=�4��\1EҏJ�O����yR�V8n�p�[h 8�=ﭦ�s���9/����g�G�ZH���>��I�H�f-L.�ޕ�Q��o>�����!B�C�Zءl�PL���^���aI8=#��ܬ���J}�z�>9�J��1�	�L�%�ov���!^:�#�W���?�ה	����==�<Lvp�U����5�>s� ���l�@؏Cό$�)"�������L���Z�`���w�?�o=ʡ,{*��5����T��}���U]����}����i 3�Ϝ���?R��_%~!E#��,�W
�H��e�*'���\1I��K�o˛�4�tm�6R�Y��n���|q��svm�8%��JL��ۻM���%-�w�T��p�{�� ��|�M���>�I��Ƀ��y��\(U���I��J���pNy2�0#U<�4����+d�@|,�^��yD��BU�Ra�v�*S8O�u�ջ���4�D��#X��G��GF�����膑�R���B nBϷ��FV�p<^��H����Ӵ��A��v�+^Nn�ɰ�˟��1gM�׾�=i�/�Jn���O��6zש�����o���N� �&p�G]?j	�x���U�ч���}�ŊQ�A�
<68$�#^��XY�$>ܬ�b����ds
v�v�A-�\HP 3�R��H�_7��J�1,��8y���W[~���y ��gI�����W �-���BH����}�[�m��x>?-yi�%�P5i��`m�?]���%&u���Lx�d@�;"�b��1�T�C�I`
��2N�k+��eX��g�t:,��4N�"g�껶��"�������9��[��j:��
��L�d����?����v�ʀrm��lZ5����Y0���).�n��S5"�Q]�oQ�� ���-nv��� �(#��B��{Ŷ�귂��W���P+!����df����H8_���o��u��iV��� S:�j�0i�� �,�,�N�˾h�[��L��0$1Z�*2eFB���\��Ϧ���=4��
�he�I��
�K�yf4'}���������NAr���r�����BS��꽥����K\y���څx�?9wr5a�+��$*�c66���T��3Ҷ?�%@�#�
�ul�76�k��@��;�${�?�	u�� �|�#�2U�&`1�9by�U��E:��v�����!q��c�
��� ƈ��"�{��j�͓���2S�z-]�d]�����S�u��r�<���BT�����r9{�z1�MJb��ن-F�5E^̟�yn�Hy��s��Wyb�Þ����;��^�x��&� �9�+@:Fl���<Cz�t*�8 �F(3�7/b]I�[?ŷv���a��'��*���R|w�H�ů�.�=�'�G�CÑ ���ɍ��_��T����ð�n��w�$����O?_�(g{��pc���'�!I�lk�D�k(�I�%�l��R�V8�Hq�g�ȅ�zB(u�.�����10(��H��~�5ΚS���Кu�H�'�~���`(O�8R!5�E�� kk�^{#�SDT�A��a���oP�Ǉ[$�i�,-�G���e�.Kg���$�/�(�d�\���4mq�M�@� ���J�A������WD��������I\9R���[�x�4ր �rH�y���\���!_�O��9kdO)��=b���'��x�0�B#Ɛ��@4�(�%V��ܘbz�1=��U+v�	�m�_���H�1��b3�]�x�AD��;%/���͉V�>p��9�w��ؼ�i��-o$�U�'����^�X�>���%*�9��$t���+qR<=��H�=����.�[�U�Cc�L���)-ƭ��z�}�O�t_��mTP,Ո���-L��>q;ˇ��nr�C����:�L��?>@�<H�9���x��b���Jl�ךv��[̌��#@3lq���� ��Li�?��o¢�b�<�g*��7Ѹk}��y:�sS��"�
or�n»g*��>9u��/�+>N�ev1K�\���%^�ղ���t%]���$�r���ڵ��~��l��H(n�.�Ť0�rL�̿2VcސB��h�	|�A�0�гC&����r��P���J|�"K�|��)�?�F��a�.����C�6?��[��O �Y`�am(^��]�b���$����~��1�a��h\�o zk��)K�{l�9�� ��Sg�#�V����]�}f�	?��딒�G��dx+/.��D"D��� �=[F�,M��-�{Xz~�(��.����Z����n�ԍ��LaD�7�Qz6�[f���i��?�H@fi�n�����\�"��,�f@��śآ1����&�3u�����x����+��0e%�t F�&a@ꃵia��N�,F��4�������l.�U���]9_]Z�J9��>��40#�Qh�Ѡ���D�u���-�i���� ^�v�����rG6����rVh`b1��.�E}{�	%I��$axa���z|q���g���Fd�l����L�w�)ڏx/��,��;R���V>�;��)v|�w}��L=�h%��x�س9�d3_"����}Ih�j�e��+��t���F���6�u`��_8J�U���K99�.�0�'B#G`W�?������3�6�6N�"ד-����u�ݤ�xa�e�,�F�&�N����B^l�L@?�C��X$
n����ܦ���&Q�`�x[H���Kd�?���x_�>�)s<�i�S����A	3W7o����S-�71D�����әX���P�U�3�d�[�g�k�/�*Z�!ܖ��]�v����{�:k��^жdU$�{�,�Y3M�y��3o��u�����,��XZ�0�~T��"&����}IO��-�Qj8;h�s�p³ b)@��#Lx��,�s	��/L��'%`Tm��m�l��kւj�=r����AQgc�& ܏�Hc#��^�񪓫١���No �3��v׀��/�rk��R|R�ˬ����?i�D��Q���-L�)nrf����GQ=�;^S�T/�e>Ș�Ne��}�ܮڠ��a2j����e�Kޢ6�8��W ϴ�(�~R�ww���H����j	Km�5�ɪ˓�(^���y=����"�2���&�#J�*er.�ek���PiS�I;s`��7�â]}j�A�M)e�U�$��E��c��Q}�+��c4��b>a~���ԕw�Tl�̦��7�7}]H4�缝���_K3��+�Y-,yk ~��2���=T?$�U�N�%kv���p�H�x�/珸պ���ŝ�|$yx.�t|<����i��&�̠Gq����'�Mt��y|]!8�$l]緄��g���~����R�*�2���E8���B����oӔ?���t����p�M���{@��ȿl�k���v	��_�ͫ��DQ@@��������wU�۵����s�(*���_
��?F�>J1w�pIW	]��� a�}�E^<k�]a�=��OQX)�@���
�#LZ��ɬ�⇍�60]��� 5�#�Tz��B���_���΁�hS㙜m=GX1�,A����
'�a�j��]��n��b�@DW�]�O���r���gX� 5*���N���^}p�c������,hV������P�j�k�_���,Z&Ay3�4���ɪ>(�3�V����;����N����F��M�Ɍ{����uQ�����n%A
"��0�h��/e���.Zb2�-�\�S�^qKU�b�2R��B\�c�;y�������@����4��������V�}Cy�霽�zy���ǈ��uB��Q�CF��z�O�=hT׮�<���wg ��.��Lg2Ů;w��@���[�(�Gm_���[h�E-�� ���g��K��ǆʇ�=YD.���o,h-����ܖ��|�����.���Z�4t�->�
N������(��ڬ��ƥi��$��M�K+���Ug�A.�s?��������@�h~�b8!��Yb#���Z"R�n0��es�f1ב�!��.Q��m���C2�;�})�Uwjc�fy!���k�;>$�+O��G s��������9�h��Za"�0sS�i��p�� )q���co��{T�{��V��ϥe����ئ�*v\K�8A)9
�H�:����+�qJ5�z7Ϋ�r������ܩ�u(�(����ز�#e�����V�	��:�졘����_J��nM��Ǌ]�A3�����Dbw�i����t1W�b�L<�_��	�<Q��ͮ�|��$rDU7<=������M�B.M.��9��&�MY'��2.��$���!���œ	@�{EGm���j����ϻ���� �z�U ���:6��yB���6`�Č���t`Y���H��$�C�[�����]��[	��y1�*���s���; ���;��K����<3�q>���7R�o՗<菍�C����!<r{u�o�W�	���(8��H陼M?���(nI�g�Ievp���7bB�I�J�
4��L̥��Q�?���\�*3Ԙ���>9�v��$b^�m�}�c��ݥ�G,e,��N��2m��1޳��n�7�m �~iOC�������z/�3�J�A���I�k�~��Ѱs�]��}�.Ji�2�;]8j�GHh1�{f�>jʨP�A��l�}_�^�T�w�F�P@j��R{��ץ'��d���ɷW8b��~�(t("&A^�z�F�7�)հ�ְT����4=���(b0�bȳ�C�"씄�8��Z�5�2�on-���D��X��UɈ#֋\v�uoq���f��G���ի���w��� Vc�p�"j�v�R]�M���l���O����y2��P^���8��!��^�ot�K"z2�br�n���n_nn)Sw����Xe�N�����q8X�`��{���-y�qK��I�6��l����/�>P6�W�=�������	^�����n��Y � ����#���f�@��v	H#�M��Ԅ����F�^�1��H���)��Շ��td\x%�e{2-�1��Դ��Kʕ=�X`���y|��d[�'���]�+�Y�!n��-ܸX� XՓc�N/�b�$&��a�lbp�������,��q7q�@3�_Q���N�=)�6�x�2)BP���b��^E��PxQ[���졕K5j����D�N�͋薺���Sˉ$3GF����r����mFX�2�b�ō2���$^�7�)���JA<$W-�@�[�Ո�A�����6����*
@
a���?hb��OT����?�YU4/S�TS"|$��rG��^�W1 �I��w3���[W#�]Zl�T����9��_hH=;��6�<�Ɲd�оhA3&�i��pޣ�J'?����8���Rvc&��D�y�^�'��xv���P���߹��ݻd��	և<qX�J@X�Y?�Fqxr_��� �ܦ0�1'�����Kͭ�b�|I*��7B��Pʤ�H��A�̂���G��$e��\���֑�R�����h$B�cc�>b_�I��Z��0�r[0$�3��%Ay�$�痑�&
Sϭ��0��6��g\c�{��k�
W;Gk�ˈ����Y�㧓L�Ky�E���?|P��^��&�\�P"�bL�fφT�p�$�P�� 8~����LD��FK m:���a��S�����h;���*���=.7�-��3ؾA����,�MџSR��/B����I	7Ã	��?�X��Ֆq�:���>������պ��p?��$� Z�)@�4���T�� *SS���0SEK�ߘ���YO�U������b��U��rT;�.�ap4Jh9�[�;T�X�Ђ�X��k~ZIٗ
�]�爍�f>O�2�|�qW�x�c�bM��#oB��6�oqt���lڬ���cmt接*����y��k϶*��ҹ�
�cHgJ"�) p��P��p�CQ����0�(�#1u($*���yhL��;����(�f�����A��.�5u?�Lm�FnSvnC�+���7
�):Y�a��b��w�-��k<��F�u���E'�cIѸ�='l}�_ 'Lx��	��T-���nj�AB�P^7��˥���j��6=:\�)	4���At�K�+��W6%-Q��<�ۆ:��W�ҕ�|�N[4t��¾��z��v}Iem�K���/���E�WƵ�4ڕ����q�J�iI$�t���˨�k���𖿮XS~�x����2H��X����
�#T�㊶�9'S�@�HȖ'�!&���DWӫh�}W��b�����Ƙ������jz���X�s���@����-t�t%���@t��!`���0���c���
�UQ/�}� �bc�ɠ���5o������uo��BB�q�B�_�a*�3u����e:�?ծ	��v[�!�9�؀\���%G�0/k+����7����I���ܦl����!��������b�,��M�\�k\�p�3oP���E�h��KZ�};�P�����I}���g��S���,XS�K�#D�l?�S��.}�o��7�.�9T�yF� #霊�ټRR��fI��Qb�L���o�͌�z��^�P�����D�E9|=aNIz�j��(��
!N�A�Pe�y��}���/9wc�*yŎ�z�3ct�,A4TQ��҈0 zp^tQң3��܉�Vӂp�nXNi�~��,��A�P��� P��c�gx��fJC/�[&�w||B��_�.�,QD����.B*�s��h��gt�2@��q�������F��5-�[N;��Z`��XQ���pH�WEĩX x�9.C���2?%���1z����"pu7��,�J��g�'�%GQ�Sb�xo����Y9o(�RS��p.��nsi Xz'Ui�ɒ*y�XK�Q��ː�w�ʦr:l��{�c�)JAv���I^|�Va��S��'^vV ��HQ�AU�"�]z�l1�'��g����n�T}n����[\��	�7G㢧�C��#��x��q/���K�a��r�zj�WoL;7�渄)���rkL��!5(>�:	��M|F4;�a:����v#����bkk�UZȜ���X���.���8��#�K�C0�m8
S93�S��V�M�Ք���_�sz�ŋ�X=N��4���eЃ)��c{J$Z`�5܍��Ӓ>���^��NJ@�k�� ����n���<�P��u�F	�`q��"�U�AZ8�P:�dB5��Ku��J�")պ�s���4���u�H{�bo������|��̶h}Y���vRc�7�J&`�6���N�qi�'낧��q��2��O���ģ�J����脼�fD��lO�b��ڽA+R*6_�o>u����T�eGZr�05l��G��V��Z#i��Ov���H>���VR^�L�qV���+�@u��?aZ';C)�*� �q��{#�u{K�b�7�>�R�e؍��J�TP3��u�hJiPh�,B������4�Ia��{�BQ�+��~�P��Ν��}P|��2���Y��Q���å7Y��i�_Z�{���7�X� ,vfg�&Rye�V��i	R�?���ERR�d��1��KhV���w��Y�������ͼ�/�^p%6l6@K�|5~�/� !���g�`;{��Z��k�R�d��	J��l��kq�ǂ�����"<��mՙ5:��|�~�ѷ~,���Y[���{����`���<����T��]��QM���\�Mb��X�0�s0@c�Ty�9�J�1h:TIv�ݲ�S<=C�y����@�~�C>C��)���I�t���1�s�� z�f��q'O�ʡ�У�G�v��u�I2w�$�}��0��V٭c��W��ǐ��`@�F�e��}E�Th:H���%'PT�EJ���� �.������k3Q��Ϟ.�����b݈#�]�s�N9�+��ͫK;�[OeX�5R_�j�0��*[���xQ�c�f/J�7
r��i�E}�2�~���H6����߇^�}�[�⻨�+d����
4�n���˸Ahz�S��i(���_����l�Uȥ}y��c&�,ќ����_-cG,/�L�����.s����K��P�TD���*|	�\�Y+���^�B�c���ڪ�4#�a� q�0~�9;�4��{���ȥ����pW�"�Y:z�ͩJ�?Q�ö���l#^gg�B]DG�	mM�S7��ց��]4sޭQ��T���^��R��(-�;��2Pq�e-)n�{�J`=����=U��b{h"<�$�4�L��,8I����d<����\]�蚘�J�ʗp���	>	j�'Ӡ:*�9jAi,ҹ����(��qz��g����� gj���^��?p�_L���Zx~�4��GX���M�E�@�
�2�!��e�c8y
�Tڏo����wy �{�B�=w�?�V���4��û?��1��9�s����@a�B'/��(|;`SJ֢t�������a_���%��7��O�&�W[�:l���&��o�9��Пz¡��[�r V���Ȁ-4r�dC�� �4� ���=@��6Wi=��e�)4ֲ����2��TWo�5��Mǵ�ۢ�	W���3��1�q��y��������:w��i�Áڏ�;��s��{�z|+G.�n�缲4→kYΒ�M�"��-9����;��V�jW�B��T574R�Ì�b�SR�6y����)�ޙ�SU����F��t�xL��'�r���n���>�<�SrfÒ�4���:,�͈��>�`I���Ԫ�S:F�l?$�U!�=���������"c&=����P
�J��?��<̀��Х�dv���Mlg��=QJ���@}k�a��F���2=�©�4�8b�g���]���+���Mͣ�Z��23�o�}��>6�p�ӫ��x�젮�{��n\�cRѬI�WT$�]s�3P�-,O��㤈lQ��,�le�*$�m�1���׍-��gi _��̉uC�Ht�bx����\oAxxJhF�RH�Q��^1��:�X���ma9d����<��l��܏�;�."cD���)�Ck���]�t��hH���t��!�/�oƳze����)ɖ���U%��ߚ��5f٦�/"C����r4b��)�rK�I��?Y��Fkp���j$��i�v�n�O��q�p�/=o��;��w����Է����iM?ʼ"_0Ж�S��)_���<
��_Ye� ���FȳCRv���*�2d�0�c��."Rm�S"r��]	�
��}��,JX����sIl�x�O�M�Fi�i$��p�(�����Op�	I}��@�p�����B�U�s���G9F{췳hH�L�M[�d�+�4������S�52	�g�pZ;�oh���6.c�}���6�.�����7��O��hA�.�[��y�c�H�O�}�#Y'��{`/��zӽtO�Om�V{�H�7y�����P	|�c
��:��Qb	���ʵE��%|Hmz�%��܀��Vw>�,�Z,-��<ЖT1�ʔI؄W��B�����/�Z�����A����	�h97�Zĉ3�;��hR܌��v��t�Y�_�I���^�J���n���{ M�S���j��8#�k�ނ:,�$`���rCH��[��/,lO������f��;��n�gk>�a��j_��N����!폠��w�Eh.�Rm�)����B�����`�Яۅ�-�UP�`1}����.梼�����8N�H���@&8o�dG4k)c����#n9$�\j�?�Ш�%�R�`�j�XTYkx��]{U�.X��א��&�r�����±m4�Zү9���0���qP�ޢ@ fR��t�nܬr�L�4�mػ�yW)�?U�����3j�{=
#M�mqm0%]��]��{��k�A��]޲1�+���o��\)������CO���G� ��6(d�� @�Y��Y8}O_����O��m�F^�;������2l<���$��ߐSOh��Kx�*�	���gx�} A��?-X�2�g�.��N� �U�fX{� K�F���.��],`>!t��/;;C�6�'T��8e���B�-"�)�Ѝ"�t9��rk�n�5TqR�C�|��ʝ����{�K[��������й �����@M��Gk����kIX`����n/��lٴ~�	���{�g��v���Z��#:��P� K��H���v���\p�:�J00��^I�ճ��p��.�=XQ����})F��M�iA?�g	�LX2J��~ĝ��=WX�k_bK��ɰ��y�Ǟ�l�b�?�>�	�}=�-B�����Mq��bUo�;,q �w�XM�!�I&6��jf�W��;�梨��6�ɉ6�7�u��3����� X���	`��1��mq���
�. �=��1S��v��؊Th��5��<�"$��K�5�p��!�߱Nk6����`Df_l@�8�E�p*}���k�6�|~F��&[yMy��r��c�� -*!���7nM/��� Z��x�2���`$�T���c��#$�m��}���&�l�%��Ż�}o{�J0�����$��)� �37���AFS!��OO#��s�M͔HG�K�WAuI���B�&	2���h�����5dQ�����4�	�ׯ�t7/��B���{s����9����8d�53!
�4Kۡ��;O�щ
�`sT����E���iЉ�YM�Uj�%�6�E0��U�k�;���^ʖp\��	wFd�?p���x��� r�駾��q�<�Pe�G�D<�@7������X�)�����c���87Z���ʸ��%�1"vܚI��ൢY�;r�2���H�-i������W�7��H��t�L����"���_�Xc#�Th>�Ow�N���y}y�U4�8�5��f﫫%{��G>: x�Tq��Q�؆�}/��	wF��qo�.�(��Lb��&Q�
�g�U�2���!sw� �j�ޤ���������R�,ZT8���y�^[<i$u�@2銄"1��s[$�-�`��WaB찉�L���<�,�����{�8�����ӳ:��O��Ɩ%9����U�ch_� 6E�0��*JW�݌K��p(ݛ�"o�\)��2�%�1fyB��e�Z!Fn�e�����<��tD�ΰ_$����Y�.q��R�ag�HDl�C^�B@��C�-���[�U����i�C�R�1T�p�X�+޹�K������B�O9y4 ��B8tP0�e������֒�,N��sS���X C���2�lZ��]2�����m�u��Cܵ	�ԅ��:��x�n+ee����m�gZ#��2(����bД)7�_@1�e��Y^�����Q$����� 6Qw��]���&��c���E;�]^�
@$��3�G)f�2��g��g)�Z$�k�%�Fw<�v�Y%}�fi$h�ϣ.1;1̲߮h_������krpy\}U �E�&�΀�����m;�5����3��v �|�����1���1��\��Vי��޺��|S��@��+�a{!��MBv�Ҳ0���0�����
iV��r5X��{6�~���ڱs�OQ9M����l�8��I�͆ "��"̷|6'&
�ZO�`��+]%Vs���J��.�Ѧ�,����?���.�9A�ʆj.��O(G���K���a��4��st����g���\�bd���v��/�@��]&3o���t�����S �.�\��)>�fG��y��#x��od�tQ�l�W�|ʅD�
�$7B�Z1P�V���6�:j/�E�N�v+ꩲ��^�EK]�� Y� �������
���i�PR��+cN��z�x���� �'&�1�k߱^�V�ѐS��Q��Dr%�C3�	U�V!��դ��x�[�%q��f�4hF���B"t��t��?��S�d�K[�� $��_�?����G0X�4DCŚYt�f# DF�b���;����!U�Ԫػ�#{E�ȁ7����z���\����l	�i��~�Lu,�o��1Tv���B	��Q:��W�,wڜ��ޱ���k�51�8��t� �WV2�^�B��W�T�'� 0<ѻf���u^���!�g��c}�RO�,f����:��қA�Æ�e�s??C�`i���6(�DcY���ᒂ�Z�\�'y�;Ĝ�ۤԄsX\X'������p���@����>�׮���q���3Ç�~���^���ʁ��M��5Dq��Q�I�:Y� �ue=C�?p�t�3��i�j�ɽ*� ��K�-����'lϠ'�e�R�,�����Jo& �,����_J
��;���5�@6�-��w@d��k,�(��|��D0a�_�4Yw�[���{g'sq��*(��rÍz����_Uy���4��C��zt�e�����>����j>w�����A8�0%��̳{��8NI�}U2�R	��o���S�aJ�f���z��gM���3�P�����b�t2ؠ���ϗq$#@7���4�a�nd����T��wy?Q{%W[0
)�)6��� ��f����ŵ��MF�V\����Q ��VD݁I��y�KQ3�A�0UaS�z�}��#Cz���=�q�kpҼ0�qF~� y��*Y]<Ȣ�5@I\�w<l��5��R��+pڭL��Gi_���G,�)0�AI�߭3���-)��V�
��� ���^g��s{I�*�y9i%�f���e�m�0�Q�����Zq�9+J�Y�r�Kb"���N=�k�G�=Ж�	J3���-����;��&�5���a��Dؽo�&�����P]-�&U�p~w-��gbyH2�)ے?� �3������a�Z&�ǘX��U;�8�tۆe'��f��x�maf��V�dE���Ժ�P��Y�o���["�E�A!)������������ϟ��dM��ј�,��]��3��M�
�B�̼?��3�7d�
��[צ�6���(��>H�Y�#��(T`�n�_ң(�{'�{Ⱦ�7,2��;���塓U��5�k��M~�&���H�!,���𿶫���'bУ��G��KQ1�dj7Ƥ��μe`PE�l ƛ���[��2q�6��bgcaVTbG�?��[{�h(����*�HnNHf�����m��)��ٗ���2v1"���ml�B��tӮ=d ��kֆ񅸗��Ζ飚/,��]D�=�݊���*w�A�N����G4I�ۤ�$�D�U�ލ�\�Oi�Oo��j�����4hYl_���	O��m����2%�����# Ч]��,
f�H����N&��{���jV��ސ�/c�Ѳv.�+�@<*�¹U'��\�E[7�4^�,cA��b	]������7D,||A��~T��7]Bҭ��CCPU׹4#`k���Y�Ы(̟�N�ص��6��r#;g�p��s��d#�[�H��?T�M":7p��N%��E	��c�OG�pf�*�|�@�,c|��ս���,�ә8�#N�j������(�޳i��_��@T�Cb��d�-�@����a�Ky�MB���S�����9vB"�1��ҳ֦�^�po"��>C��N�ì������v<�4�:a�rNp/��ꝼ<�d�ڞ>�s3"8������;�4� -�w���/#Vފsf�����5lT����ڦ*YQ�wm0(Q>��Ѫl�,�*���~B�
6�(���u E�t6 S�ϳ�2���A��o��hb0���*��7�p���$���3i�Tb�>5yf�7�d��4���=�7�ܙ�4f���-���?e�)���۝~@|,���γ���į�]�@�: ����P!{�ʆ�4��S���8`��#'9�w� ��M�k��c&�jg�'��A����W���WX^t�����7�m~�Noi%���`��s���Q�ᓼ�D���:r;b���;���;u>,���M�N|�+�*V�����	R����DX��7C�ҝ�BBG���?�2�J�!�R���
`�lH��}f��TsAQ�rXUΛ�6Ýt�B.�����ӳއ��-��AhJ�^Xߵ����L�~.��(	J��T�ڴ��^X[ĉ�I�-i�o{��Te��V=  X�Ht��=6��d��p��2�O�.��i�&�|�kN/�%���F��--"m��po1�w#IĄ	[�u�\LE5Xw�G��JA�bF�u���ܶ���.�VS��E{ ���	@lEb�̹�$t�K���%.�����/�K�`\^���>�4�툙i�
��}�>�6o(��$�p4]��9~�#<�� ��\��)G�ϼ`��θR:'R�"�<�c�F?ӱ�C�I������`�K����b>�a:>��S�(�V����=v�2�P"��ev�ʯx�y��pz�8���M,�3�����������6;3ﶖ?�XX�x~�9�$V�� 6-U�^R�K=�0^�w�Z�t ����`G,oM����S�?��٫c
�
������hA�tc�W��Ez�h�������]
�Z�3�[+���d�*9��
��yɯ��U��7b{��B͞ �V�p��f�k6�Md��e�{3O��r��1@I�x�g7���ZXD�(^��ߞ֑ҞM�xi^| �M�HS���C;�oXoՕ4݈�N��2v�&����J,��-~'��}i�Ya��2
�e��	DQF��l[��0�P�\�1���&���T��P6�jX���@fBq4R`�٫L���WQ��fe<��#�������V���N@G'��{J%�%�	�jU�k����hn��[�I�/z|�;�F�VX5��s�1�"c��,���"�O8
��=�-|o�-�w]�m��,h����ݤ�y'�{{詨I��ᵮ��'��w �w���v��?z����M��c���D)�XCJTB0�:�;_��Z(��� �6ƉsA*�Ҳ�n?eZ���6��bSn,"�h��yz ��#���:�z	I��%��������Hn&�|z�Zڌ�#\,����Έ0)�騱����6ݿW*@8\�S])~����t��`�]7d�g���T5��m��3��xi)`p�1�(��-hOB���������g���0.���o�i/�޺~ht��4$S���y��"gcA�*��aQ���tG��`r��Ú�yA� ��M�	�1��-�5w�݋ٗ8��HT�'�ʄ�|K�T�� l	��ߢ>+��$¬��y�B�����p^R��x�����zA�k^Oլc�m�-xȹ@�XOQ6�������S�� 7��%�a�1�|;h�4�/���6��e��Z���˳���e~HF� �x�gO�-L�z0U�0��%|k�I�6��r	��6D��U��w�W{��9cL��v	܅���?��a|>���Zj�����Q?��G�~i��F��R���"���M@�>�Nk�|]����dg<��,������	�I�A֜��L�ۘ�k��v�˿��-�=�h�w:�$P����}Gљ�h�m����t-v{���w�3%�.:J�V7-���U�U�;�u-�ߎ�^\���,���x��N-�t0I�O�H}��	� pAvɟ�O�ԕ�5*��k�Z�󡯱�x=[�I��g�
��/�c���Y�q��s��=D=
�-�1d�hbR>t�BdM���%s�MN�Pا���z�B:�����(�5�ǣ��*���v�ڳ�y�o��yd?z?�_GXÔ�߰�fG�"��L�[�7��(t�A��7���+�e�Z�:�5�90v���B��Ն����e����n��?��CAbG�m�g ��u���X��t<�.2/ee	�z�|s}x~��?��L7�ƼEn�>�=e���>�3�=Ә	x����,,`E��Ȓ�sx�0)g�$y�����Tʌ��p�jC�ͥ��쑌-�U�Z;ѠjF��g�0_��vz��Z��?}ﱾ�m	���݊ ����)s~Qq��!�2�,"��{N]6b�<!�(a����ҋ��@<�N��K��U��퀛�ABXH/nbh�GhH������ft���wƎ-m'<:�D/��1	-��% `�3%� 'ћUY��J�+y��H��[-� $�X��M;� gM�-���8�����wP�}Q�����#�T^��`*���أ����a}�����{�������;�W���0�����F7W�qL48d����*g��T"�O��"$���y�N�x�ױ==Ȟ�����D�V�5��gwY�4��x���Gp�j��w�;:m)̗�8M'�L(5ꮼ�6aĪ�9#��YΖ�� g1�����7(ԲПJ�
\�����������ۈfΑ��%�Eɳ�X�������@���<ڨ��n�����<)Ek�W�dtӑ�I=��n����BEY��}���J��/��K���x@���b��0��KT�Z]\��֋��(������Ո�g/;�"�$�Kg fQ�s�#�$d|Cn� 졨њx	����D.8`C�E�	���b�����Z�jޫ�Ǽ�	]��0����(L��ֺk�>}R��p��Z�0g��ޥM.gL_��&ET���qѬ=�\�9sW&���3�|�$�ė�� 66���jq�28�	�L���i\::W}c����.����}�jW��� ���$���E��Ӽq�{�Oo���e���^�	Ћ�l!��,���UVm���w1}�l��CNvs��2����r�J(k'X�6��-L�r�G�T��oo���Nn+�0Q�����77�]����s"J!]���h
�waT�ҳ�y��3i�Cj�MA� U7"�J3���*D�z�VI(��\
�T���\k���їZ/� MZd ��Xl�$�YNK��l���%�PuO�4�β�n�N[��u��|��0*M{�V�@g�%���}*��*��tD�W�F�u�g9!W/���_�K����e�i�X��/�<Ě�H�ҕr8B���7�}a�}i����n���e��ci!#�O������z�&�� d���"]��j�U�;s7�F��;?��K����-ݛ'U�>�˒�q���R�'p#ׄj��Q��IMU){�C�7�)��$�g�,w̝����Gqr����Q��(Ӡ$!����@��w�Z����f�Կ�C�k(��]��l\
���,����g��:qu{iI��!M�_�]Ρ$��XIy�ۙ�����ߔ}�)�H��O�['��]qԧ%���$$�C��j]|7�4��҂��K��A��LOٸ�f3{��x0���n�o� �~{�N��[��J�I��1�Ƕ�b��R8�dE���4�fEˁ��x@�,�g8����f|-�$u���H�b��<)��b�QXt��z�2C
Z�I0�-�W���<�?�GeL�}�^��g����Q��=���e�;&"�}2��>�n�Sei�v��O��Լ��+�a���#*�z��Z8�|��$�_N���E�����J��*K��6��+ɘ�q������ˆ�)�������N���Ɗ1Bj�u9��#vk�M�*4SE;u�#��=� 0��j�K�S���Ό��V`��;�"������v׭b�W��	R�<!�,�=��V9����)�!��,�m��@�x���dಥ8��,���@�F�atrdp�����m�FRURj��I��b6*���ݹ�hT��zw��RŐ�H�/����#�+p՟�n&y��I0��ԕ��|�Keꟳ��G�F��� l�e'�H��P+�̊,J�m�f�qY+I��,�kt���%8G����X8^5umY�Qle�����8��۪�m�	�/ٿ��N�ʗiF��u4Kd��@W��:-JE̪_]��1�x�!y�G����C4��¢!��"�Y�?a)�2�8�a&�� �]��~�[
Y��Y�S)�+�����{Ī:H��4�g^ �È�ߥ9���}���y���%W��0f��Z��;��o/��x"e����������'�{^�)�%ş��;�.��TG�[�-�GTi��h��f��#�������_�B�)����/����ɫ���z�v�Z��Z�\#�.Jic�Ag0���q��Tw��b꾹������`re��`�/��HpL�A��t9Y�C�)��"�%�-�LZ�������H<E9�iܹx�*L�,�B�2�C�{�1�M[_��<�X� ٛ�_`0�r�g�e*�2t��e=���ȃ\�D�$#]"�u;�>�r g���:�E쬯��;nf��M�?x̱��拼&">�14J�A�U5��Y�8�翠�S���4���x痠���S���ʉ�͚/�1l�M���l#;��N_�it����>�R��p�=^�޽���<��+,��U?�����'j��н�ݨ��5�v㻲E���*�80�D�o�т���|��b��%x�sC˿�|��B��HCu��-.�q)�ɶ�8%W*��$o�{�QT�u!�b��0τ!�L�׍��g������[��?�S􎒧.�~as���q{�gOd�?�
@oRYb"3�B�0z�\h�m>�pi�ߊ�����Z���s��_tR�h�"ј���4/��esvz��n�}��JJ��1����,�u\'d�gw��Py#�f$��}tʖ���-��uտ�U�[�s?LƬ��TM][���ik
��s�#a��9��+�//ƋS=���t}�9T{9�[?N�B�� ^niB6�����~��ć�"��@��0i���*��/�lb��s��okmv��~�p���5yic�4��ۅ�59�j#�_1[1:�ɓ��w�=X���$���.��|�q��$m��:��G��*���|�턠�Q q�� �3�EO��,b��:���J�)]!�y�Y�w��pq��D���]�H<����Eɸ���X=ns��9�����F]���Iuz|: �����\����"D#q���1��n�0zqԕ�x��[9�$b�'	�$���1������)�/G���i�re-���0�f�&���4����c:���w���Ѥ�O�!��Q�$���I�j,�O��Z=���N�ᱱߨlȤ�n�����]A�f(.������y�1���4�L])���JZz"룻�\]�m��:$}�>�j�%���+Y,G�)�Z�ɑQT��l
�J�|咏��sxb���I
�\�\�v��_c�8W��:s�#�^�	bS^�Y���O�0���h��>�meªl����$��D6���Z>~���e3�q���@1�
�I:UmdY�n{:E�3�@�)s7P��yw^S��C-T��N�Y�ue�<
GyI���&�����ղIĜU��~�D��'�	��Uv
��J��Cr���f��Y��~�!���܃ԀL4C��RW��O��P��Mw{�#h�V^��$r�� �I{/�Y�@�l�+�U�bM*�*L���F�k�9,��Fll���
�8�z����^I����Rg�w�.c|�/�`�#�5��,�7�CGU:c.��o��#|/՛������8r,��}��f��k2�����m~r��Vh��`�#�;1&������%���f�EV5;��z)��JI����6����*%�U���/a��]���!蝢���2 X�d��#'�?*�4��4[JX9��gN��JY�B�N(J1�F��oqP�����_�Mh]�뛼%�]�����۬���)+]D��2�%(_JKȖ|����������		cd������Ao�۠���,PүbVq�4��V�2�����8��[�t�Yai���9��Ճ��\��G������al��z�0���C˭����<
ڿu<���O�}y%�K�c�o�i���<�y���g�;��p4�z�d��vǴĆ�}lS�̗�#� 7|�@��p��R�ۀPF�c	wg'}����;�X��+��G���2k�:o��H�]�.�N�_�MzH$��wU?r�Q�b��½	T�K�<�4�M#��
b�MܷK��Mƚ�:C=��������K�������uИ�?ǁF�$.��h7Q��ȌUeGW�z��k3e���ɸ��������B�8�a>`��kN���8ݷ��"�F�1�'*T��=�T����ɒ�S	{%v�T��P�b�ҳ`��Ʉ~,�a[5����ʱ½��R��)��k�y��B�M�$��=�e��q���ïxB"J�����,��{i���YqWt�9B���Ұ�=�9�	��M���l��_1�1�mr�|���T�3��m[c��\C�wN0�.�ۦ��?�)#P�e����/����T����6S��+�X�]e#=�6�UԴw����M��;H�7��q�3d��+�sgb�UÞ�Ku�%�c��Y�x�*0��E .N륣7�F���|��l�G{�� ��;�0�崮
�qy�}]D$�U��Z�~0SS"���D����P�D��c���޹!�Qy�����.�Ys֑}2�0�Ere� �-��V6}7�Qejfh�� �V$ȈU�_6j�YZ0�vS+)�PPr���j�z���HW����ĳ-�������?qހޛa��g:�Œ�}H��F&2ކK�C�xko��͢
���� ���% ��^Ƥ��L �6�>{ݥ���P�!Oޥ��a��2�g�ފ"�?��>�g���1�?��m�a`Ϥ�h�T�R���mI�?HjZE{���_Y�s:��8��+x\t�|�LmXTN	���\J{�J��$ �|�O�B�����-������]�b���5�w�_[ 6�. 9���]	�F`�lȧi5j�N�a�N�'%>ߙYn�t�VE�^��w�Jb��f��m� W6@Go4*Iҟ~O����2l�`t<g���'�[v�sO?X�k�����w4�W�$�h$�ub��Kؖ#��2��*���c��se���xb:��:�����}�5 ��b�~G��m�W^��F}�`;q����E2"̿��E�LG9n6T%�\(b�q�}�Co�٢䩑�`$nk�+�����¿�q�Kg��I�	+35���~&�ۥMo��ZBX��݋�R��%�0
���H�J�]�6|�ڡke%����iƦ�'�Js�:QPy��$Erw�Р�G���Y8��J��nJp�4ӑ�w��S/�H3�dI��9��Y
7�� 1��o���s�=�I��U=�(��p��ᓕ9���%�Z�
Ň��������(�z��Q�k�f�� %�
솷����m�S�}8�4&�O:'h%0�րY	O�s�	�A���?���@m��r�Q�/�a���j�d|NP��B���L>�/��kD��tޱ�W�yϱ���n��n'd������]����Q
$]��h�����>���.tg|iTr�{4ؘ��x��Hr�ߊ< ��Z�~�%_�u��Zq.�����J|L&���J��e.t9i�#A~��Uq.�MImM��IB}vqKCN|Q"������E�����2^p`
��{z[�>�~�dn��7��=��p �i�� �������3A
�7���;jP��8~�x�����<m��@G[�@XO�f��/c����ڀ�1�V���[\���:�	�0�RklP$il�@*h�bA����D@7J���7>#�$S���`���X��A�3�D����j���v��B� ����EUv��N�M�]�,�)	�I�L��曱�'�� wn��������M�|�-ۮM|�~��#9C�ƹ�(^m�kc3�.����`�������/s�n���ņ����z�eh@V��$��8r1�S$ܞQǴ�PI�whK��z�� E�����G�R�U!���tu�#�`�E��0��:�P�2P���
�(\��/�{�.�Σ�K������w�J��H��' O�]�s�����-.����J/�s:��@)���<���r��*W�y�r18��58r�
T�	�E�	-�;�.Ld4�g�/A�E%E� H7���j�a<s�U�`��Ē�T�m�÷�����}A�99[����(��c�+G��C�a<t��d4�;O'����쳰��I=�"�Ω��_��B���s\�(v�О�{���QB�9z9��k��eC��}2W~Mp�� �-ߘG ����U7Ja��r'Zkv���8�m�ҋ��y<�3���W\�1oa,�s-�_�_j�Օ4B�x��p�e� ��t�2Y�Y2�i7�f�̇g�:D������&k���)�����<���3H9�0rJ;յ�ݦJ�`�P/?2���W���֮=�EYm�}B���=�[�7x�Hmp���[�ef%�*\�]���3��X<wU��_���^0�>T�+S��X���&��
f� �ݧ�+� ����4�s�_���2����cSY��;�Ӹ��t[� y##���hWutҮ����X+o�o (?ᇳ��Y(J�VݹR�W�\Dp��`�7Iٟ0� �u �9��5�gH���%"����4���.�����Iޜ��="A+n�'�m36������aXHPЈ�G���e�x����^4�̦��oK��%�҆�)>>ì�A�$uj�E}{��]���<�؜��CB/����[�}pƲ�=upu�m~?�u�ω�A6wV� �ɚ�ڭ��uB��-��ƙ��d@�Dl,7(/x�u��`���;��G�f���4"/�1r�K��$j����|��尬�3����N��e<��t/�.��}��޾/2��2�J�����$���`k�\�������CXl9~z� J��i�y�a�Q :�߫�iӧ6S���K����o����8Τ j;���փa(~�QV��E%6"��<���7���w�q;P�.�S�
�pg�&ΎW��M���B���V�89���8��� p�pP�&N�*=@��i��: i������g�g�5pt��fѣ5��\J���>�]���{��Hn�g�|$ �H+��Wi�v����-";�~6z�j3��ꉌ���A���j�bs�x���^�^VnA����u�#�:������Gg�P:�͗-���fh/Y熦	V�� +��m�7�?�ΫS��5��>��hx,�bdE���2z��8AV��&@h�_�AO��fL��	��Mw��a��	^�^��.�Y"APת�p������������Izl>�"\D]�s��$�Ï����g��� f��aw�#�w�ϒ1lɄ�l�"����#��y�th{+3��+Sk�I���g��@��Y�W�G�ݸ�H]/`G�~��ޕ��i:��ʻ=��09��X	K|� 8I��14˜����"t�fe�5�څ�
��S�z����)'�t�6�g@VF�
h�����j�%�п]	A���l/��`�
���
�տ�$k�H*��a�c]9��f��P���}���G:�ʑ8�_���VvgXH�X�y.��p�]�r	}X�֊����ܮZk||��ь���5
CeA�}�^��`��m�~z����8�ʨ)#�'���#�w�=6�DX;�%���
#�6G�v+��W�j���=cJf��h_4c\3���HVf�q�fG��'&�p�D��P)?�T��>���b1�^��~�M r�n��#g#�[k�Q&�z�UV� ogKE'Il{�fc	x��\��b-z|ٚ�� ����_��:D��&��e�Pr*��z���'ƥ#�<�R~��&78Z������@X>~�	_��BN�3o	B�'zl�-����f��sYԡ���cȽf�?cش�[�����O?�v�׷/3����俋��ǣ������.���~d�C���z\1���a�q�FHx�Eӹڍ�mS2�V��[�<2)A�Ã~���f-ca2
��79;㌐ٰ� B"h��*���fN� ZV+{U��A4Q\�4����hx}ʉ/q�7��o�� ���r�({�Ʒi���8|& h\�4L���2� K�z#y}���g�f�E+:�1��E�5W}p�z�`a���B�T|��������!���~�6"�������Usg-�����ݧ���˜@?�N����H��"Έ�3�z��zp������[�me���3�1\
_N0[�rժ]R��N��,��8ǌ$���^�1=�ON�M.��6������{t��͡���F�����H�8���o��pT	.p�Αf@�a1l�Ã�-	Fg��u'x���y|L�x�w��N'5!��(��.�S��c�x��yc��u��x;G����q2 ��Bvw���(������b�W���Fch0�������D�a�dף����jK�/��Ѩ���Nw�j����P3z�� 
�+:��^I�('��y��F�ĥ�+I�5�S���n\��6�����^#�!W���ѧ*��u�!\K�*[�]@�O��]�1Ôc�qG4�AT�R�3�X+lZ<U�k4��'P����KPAG&�Gљ�-&�֊������rh/a�5�]Z^&(\#�Dj%�=���Z�^�Y#7��T̔�1Ϸ��
����m�,,Onu�3mx���=C-�����S�A��XR�g��m�+\����|ߪ�nt�e"�'F�阘�#^�&?L����[�Q�Ĵ�3
���%z�0G1?@�1��ȞM��VS��*�.��%���Lw�^�O�h�^�"&��������䓻����]���4J�.��ߞ��+���w-��H���"%UG&�	ա5�A1`��k��I��SJ�?@�Ӎ=��v�����g<^���3�����7�΁m�l����t��[��&�|][�&]�5Y��I����{?BI�ƒԧ��d�����&���gH-�ļ�$��8ՉOW���AK���ӌ�6�5��/�>�}�[�?��>�oɤH��Ĉ����_i�1` !���+�	~���W��8�!�
��b�����t'���oy�W��	���Q��Y�n0�Xd��J8�;:��b�?GW���D9�3e�������:�X�]��ˠ{�ӶR)ؐL�� QO1p��̋�e�H��%9""G�΂��Hzpjk�}v�� ��O�Ŷ����j����+W��N�%��~3J��Ɂ6��8�0K�*-��a0��V�Eڀ�ȴ��d�g C}�ѿ�7�� ����݀��U�#!��o�K7	\d�.+��zx�^�$��|^���A�Oše��M֥�EGv;����]�D]0�6��2}JQ�� sy�@H��W���/�S$�>c9똻�����uvS�g8����|E�����-Q#�@?�~Q�m���X�1]��-Vg�0^z��ao:�*6���VӮ3��w:FU/�;*U��&�3]/0�����#���QS9αQ#c���	8vԈi�Ě%����>Hz\��gX\�g��L���wW׺��E��5�F�քn�9؄�~y|�%C�3����6�ձ2"���O3n��ҊQ�u��U��I�9�\\N��I�؁��W*�+ }��Ι���{�e����u�^ $�0
��5�Z�j����Ό)�}JK�c%4d��,`g�6��cy6:�,9���As������?{��A)�?۪z �s���{�e�ƴ/� �q�:"�Bxwv).`������ق�Z�������b#�n���#�E �j�H,P�'N�Z$S�K?	t�����q.F�\�h$ ΁,�t��PRl0	l�J�t����+���[]�U�(�ac��y��7w[jň�~O��s��L nZ�|[Tv)��|���}�M���.S��IX}�8끁���r�J�0��X��,D�\5'ww��6X\=+���[��'�-)+ �!ɢg<�����RD���Ҟw�׉�P���!��y�h�^(�	`��=�/��6^�<��R&��>n֙�����-�����{i:z�eϨ\[���D�t��Ȳ�?"9!tT%{�b|�P�\$ڿKI�D�?)�:�ߤʛ|F����B���E�]|z�+�=Ys��nW�2W`�>�����P�zx��u3���qe%�2����b�⌿G�ͬ�&
IeMf'UC+�[_��f���$��N��F^_S�[�r���j1M����)�]޷�3q[Y$cN�?tH�4u�j����S��8�6�`��4�<\I)��MR�����r�����c���:�uH���$4�$�?��ؿt�������#��p1�qhq��zT�DU�iF~���+�4T̴񧣧]�Z>Dy/8�d%@%_C@;)��;�dolw�%aU0f�C]վv�b����a~�n$~|���i���6<�%��#�S8/WT��(����Ӻ���=l�/�۪|gAG�ls+��R�<� ��Hw�}P��k<��3�ɾ� �YW����8mP�]֧�˜�/Y+O�b��Y�{w�_l�I�'bwE��>.~1mEw�^������Am1?�M%v���y�|Z�����o�X�2:�� �\e$~*�Q�vۯQ���YF��k�(ڙS*����oAY�5
W�hZ`�9�z��u��s�&��j�upID�'����*y��-nq����9'��2r�m�v��K�������ӾM��T����X�r<�C���i85��>��>�0���[>r�QE���p$�f����­2'�d�daN����R�����*�%���9Ӂ�����!�\
CA�T�`�eX8��F���]4.&O��	��$�v���ޝ�
־1ipM��Mʈ���J�Z�΂�0��Q�M��Y��w����2��¨T�¦pfI����hIb��e��E`<�[m;1=�J�x�U��g3�Z=Oϐ�O�t�٠b\�;I�*Lc�N���:g{Zp�4��<�|p����k��w�M"܀>w�w*x�/����)� ōcZ�����g�5��6�pj�U]a��r:p��s�Z�w�w�2�y݀;�+`K-����j���S@5�e��S3O\O�mX?���HX�(�`�z5Ih��&�0����]F:�r궫4�z^���m_O1�Q�]Q�l�cL0NSދ)I��������U�V}3�����zNqb���Ձ<��"ڡKo��_���E���1#ybĈ�L�wQ�h�a�9G��f�Q��f���?�5�N��f���E��,=�4�<I�p�����=L=ߓ:�xQj�k	J�^bg툗{i�k�)f������R��u=Qf\��(��:�{&��$;�̥����y,��;G�p�'tg��@w��Oh0@���+��cB3]K��fB$q\)FޱrR0+���`"�=��~:�Ȫ�}{�3g�I[�*�kE@s)��٭���	ǯ�u�����A��)�?�#yH���i��S�{�+�l4�=@[�qU�c��A��MZ���Ҩ5�0�H�k��jvQy5x���x% �����G>�SY�b��ך��_������z���F�:��
�l�N -j~��#S����������i|��u��<]kA`9E3�[˚
?T������	�w�9�4�JF��|�8�%������&�^�<w��h`�e3{�ύ��T�^ӗ�r�A��۴L����Jgx�"co�|�u��[j+:��ߗ��Ǔ�a�t���m��4G����ᖫ��?�1ÇAp�3S\�LH����N�0g���
���F��l�qi1��)RW@����C@4���,�;�|�,�8�2GH��-y��v�x��=K�J)�o�]�묫e�`���[��`,��U�̚�1X�]z��-q]�W��I�E_$㘚O��3~oq
��{����@S�,�����S��*M����x�f�t5�7��y���}.�3���%W�����U���x(��o#8sht[���1��d9q=�<�՘ �|Ϛ&�!����SB�j��0Ӫ<�(��ބ��E_�� �&t��{5�W+%:&\3�n��~��9��w�4)+%��(��V�L�JP�t�*_���M�!����%�|a@V���?��W;��d$	%^GVq�s����=��m_#���y:�숊��$�3 �3:3i����B�l��}"�%�I!1q�6zl΄��T�1H�H~C�s��n)��R:�iW%]\=r�W����]!K�&Y��x�"}��Vn%���	�ag�'�p�<eB]�\s-����{e�R$�6�����]��?�i/o?#��kw���	��6���	,�y#��P8w,��iZ7��
�4�k�������K·1"����G湾n���ZD�,L&��e*���?�u�z����t�@��˰}cE�B�s0]�����ƍ���Q ���8�?d�#��j?���<���92����|�T`�}kjns1�ރ�I���)��\g��QQ��	|��[��h|�l��KU+�iw���o߮~W�f!߽�|�DOV ��{�iR�����2��.M�<)E~����$e�|��{���\�,}WϚO��<�z���Wjc���w�N��7��U�����*����7x�6m�WnС1��B��d͊���.S��,Y��~����Q q']��	�웲!�^ae��ӎb�zY&n�� �J3P'a�E��!�Q����/��K�X�����e�~R�3�w�B����%"� �D<��2w��N��᲍�&��
3�/�&.W+�h��#���o�2况��(+�LG^��� �r�Scd���|-��.�*��D�A��:�
�=H�V�3O����6uK�����M&0����7�*�͙sIll��po�I]�}Sb���I���xT��a�:���O��o{�&�t+���cI掕�*Ž	�<w�E�e9�F�`�ː�nrb��?���g�H%U��ڲ����L�S���k�i�u��8./��`�u��X��J���1.��G��	-]΃(铳�0�z�8�?�a��sV"zd��,�&_��Ϲ	��4�+��.��������R=��cY��m2�p�<HI�zd�?@�8��F/��RMo۱�?��G~�����2Rȭ���ʮ�)U;���`�L(�?s�I0;���lS��Xk��4�-tQ��T�w�e�̍KPr�Vb�����`������ON�e?��͟5��AY�{A���Wg}R �&�S������&G���Sy�0�����G�s�}�:��B�Q`I���"��ʒ��o�W�Cg�(�,X��mY�7@���#�O��l�R[VYɾ�a��xPW��AM�/C֠*t��}��K�I���9&v,�\K!:��h�
 s�B���0���ғD/�J�Q�{)�� '>i��~-�b4)�`�>N� ��@^�GPM"��L��,�Ju�V�n�R�А1{���q�"�N'2�+��;[;�P�D�{�kS%�u�9�o�$�H���~d��q��a}�Pf����-A']��������F������Y"�_�_�4/�t�b�#|P��j�=�OR�M��
e��/ƃ���kKJ8�d��j�����}�Y݀g^u`^��;6��w��RV�����OG�PY"0�ƏV��9�s�{$�<�Lfr�9;�%���fp���D�̀�����~���a��?V�[#���*�{u֗�'���C�_ķ�,U??��L�a��~o�<� S��[�1c�	4����@G��)�Nq�ʰ���_�!�%�~!m���K�(���7��4#��r3����E�VȐx߰-cD'\(������*P(Z�Z�a��]��W�1u���zM��s�:7F��VY|�>9KK��ڻ�c0��ђZ���昕Ĕ��>^Z�D��$����Xtt�\\�XgT�r����)z����ߋ<T������2�� �f���ؾsO$�V�G�b�;����ay���z��l��lD���5�rj[�(�V�J�@�OF��g}ʪm����QǙ��)�5d?=4g�ۢ���y�U���P�Qq��sZ��Z�{��n���Ț�+"��B9� ��IsT�C�Al:��7_�!G=���lo���=:�$QG?dT!�OZ>������P8�m�����pO��L�~9�s�9?z���W��V?��LC���ev�[8�93��~��]6Z�#/箉����ᙧ�prj��q T���ئ��x*������sp�B�����hXF\Qykǳ&�:���'���㔡u�C���c&/J�{ѫC��N񊱑M��ݞ-.���$�fCt7?`��m��AU�Is�^?LN�����}}\/mC|ؖ�p�jO ys�
�ѪT ����h�6�n�O���?�P������}Zysml1��4���4*-����r���D���_#�ܖ����/��a�u�Q%�3J �ӣ7�SJ<�@p�B	��~ k�[��Y������K;���f��s��DF��_�b��T�?���~7�@��͂�@�������Ȭ'3
nƭ��Tj�	Q��g��$��ʾ1�c�xu�݉o_T!�?ā�G=)IZ<���J���b��՞\4N�u`��q���W:��N't8�p�=���zm��SM�v��j��`��O�	��t�k��4y���u�O�Q�i@(� C�WO ��4���~p�Gk|e���]���8��2':~���S�)����1*�o�ļ?B�4��e��S�=M����p��\��"�)�:��,=Ɓ�$X��ô�X�+)�Ҷ�-�h���04�ｏ�
/{�Gh�'G�,���̿�Q 9�U���A�O�����M����)גO�JqP�X�/%xYɷ9mE��Eh����m���%U�|o'�ZcT�XP����~>jX�k��m\���1���J�?x|B��a	��ٗyRD��K��Hn{���S�_&��q+��G|�U���D�� g����ZM�yC��	C_�?Ȫ9�џ��z��Tb�:~ql��Õ���#Sϼ��k�gcY��zց���|ψ}�!�B��_H�77<=��(��;&�@��#X'ٍ�Rj0R@b嘡�T�M_�(	��ٖ	A�=��8�:n5�H�w����d}���X��>��������-�.�����,�rE�
 �#b��2���l3 En��s3oq��~��6�M;�,�0J�M%�b3���,/y;W�
A��yr�	D����8-nH�2����UG�CԐH��j�4�.���,�D~��[��V�� ��W#��p�ѻ)�d��r.�t��K<NU-\�M�sPb"g�#\�qYew��3[�Z���p���b���M,��>^Nk��\((TH��u��HS0M�N#ߐV��BR T��S,Tv� 2�?V8��[��m !�1��!���}sUU�Q5���	�~�J����y0lb_��J��,|���ek�2�,�iy}ȷ�fb���
�D!΂J8-E��t��0�j�i��/˗NFF���]���7�
(X^1��&�W����"a{�?{���m�1�EcA=�|e.x8��.!ω�V��>�u��@�˴!7ckݛ}��#�`�E^X9�T�>)�)�:�Z�$��������1W�VRCO٧��F�ʷ���G���_�=L@K��u��	���"���ET���j0��pߨ٨��cBbR�//�����tƗ��;�7��lA!\��*�Y�fD m�7�25���Y��R������*;��Ma6�q}��QE�c��\�,� ��3X�iن%�-z�H�u6�ǕD%�D�I�V�<����,}���+��$m�d�^	j�	����v	�f`�T����r���[Z�kc�н��X���+$=��S�&��-�v���~�/�]����=_H�(�xp�e���V�c���W�O�&q��᪥B��ԧ]-��$H`���o������g�_8"���8u�oP+<� �� �Щ}I�7Q�N�rj�
Ws��Ŋ(����f=B(1�&�V������/$�s��,�6�0p�쑺�xb����=7�l���|�H�Q�C�Ռ���[��D���Y�Uz��T^Q�k��#�_:�-o��Y΄���y U��_���h�����Ͻ>�_ V1CX�`qfn��gL�C��`���e���p�OP�W�����e����n�x�b��;�RZ��e�7.�\ݬ����3D�[X�TzI��&�23�"��H�y�w�)F�Ḹ��vO��L#;�q��l�)a��:�M�'d�Mw����d�䀸5�H����/��?]�5?`T��!ԃu�"�M�?�0	���� ����H��f���s�����`\���p�N��qf`�B���4��gB��FXAD�����UA�v��8�=1z�֛�LL����.�����S�ߜ�����h� ��Yˣ6K�{]>^�^�� �M6@)�x�`�}-?`��d���s�O��6����XԪC4�c�-�l����
m����t�HZ|s�� �Q�˜î��|��2U��{�ܰ[)`Re��cy^�](��c�Z`�-0���]�
�SM��kDD�l���i|�[y�
5��{Y��Zs���V������i���йc�k�'Y>7H[��.��K��H:K$f(w��aM<2̥�ц���	�4T�&�.��ە�SM�wU�?+�-	9�ڟiE6Z���\��x����P懖��8�?Y����=7g?!��Ȉ�c�9v��5��ҵ�)�Jy8�:�D�.a\��5���r��,�њŭe@�K�U�e�����;'M
{d��n ���T�O�V��A������p�_��5����o M2�����L5���F�;'Ȏ.�%d�(:�>^l��K��n�� �(����rl��' �pΏk���=[C��\y��Ft����=���p���b�\�SR_�%29���mP�2n��"*,{{�N��$�*V���B�"P��.DoH��r��?ffft������_{P�m+|Z;�ƆoWv'8g-@�378��;�61%$���\��uF�ښM�$i��hw|#'����~�P��֌4zBû�v����Y��.sݰ��3%t�|j]~����$��7���Ϯ��@|���Ў�V¦��.�N�ʙ��W͒,Ʈ�-ΒmP���u��d��q��9�&�:� }D�uuwlqVK(I��`ň]�f�CL�MwL�=�%_����J��j�-�����fl>wvgw	a
��Ozxw1dO��G��CQ�/�� �#3�ρy4�ϊ��"+v��7�v�z:j��KMRF&:�_2�ڴ�����YL�%����^
��Ro��B.� _*
.ZJ
�/� Jz4Zlf�`i���[�M�DS�a�T10W"	\"4�%��8����2ՍN�r_a��7�x/د�C
E'��'�*ם,���m�M֕p_r�?��?a�LB���ѾOh� ��d��<����3ؼ�>t#����~2��z�����СNh��NE
����}��) 7�����aߑJ�l�c�ϧ=I�[ZN�ĝ8�dlHI����ų�53t���������%
v�/|̤�j��^�>���lQ$BW/���Z����첍D�f����˕K����|];^�=zh!�}	t�H����II�G%����ݗ����X��%��9%��?-F~�xڷ5��|y��;�z�U8E����JV����إ;��{J�|o�sa1�^ � ���R�O{���(�ƥ�D��>:�������M�[;�~�u��xuԑ�JЂ4�$G#� �@h�zI��2�ұ�RN�Z�./^�	ˉ��]��XPJiQ�j���Lk.��k%�~�[�(E[�qC��J�~0�+q&=m����W���0��h����V:w�������Zp�7(}y�͈��ݪ\���G~����L���W��t�����?W;��Q	�=�>���������%�5{/e�	�!�HhЌq��h�~ض�s���Ҝ���K��Cb<5��
5�O��� ��f��GhFE��&��Ow#��̺���a
4�J#�Ƣ�غ��f�g:�B�����w�7�9�Jh��� ��d����-����T�HK���P��g�{81`�/�T���g�1Rb�:�G�1�ܻ�n2�:�`�B�G�z3+�8>��e�0+`B�1��ۘ;���Q<�ﱇ^��YD��X�'��o����5���R�W������H@lj̓$+�
ƽ,�[ށ�fh�&��"�������Aw+'��B&���U�#L)�7d�����!�~e�>� I��~9'��ⴍ��8"�֕��?5ý���"�G�����k�%D�i��;(Ϳ��#T?�v�1���I��{�s��z>vC��[Q��z�CZ$͙����:��QD�z�KQϠ~�).,��3A�:�l�N�3Z!���P���?��Vo��:�̯�'3�p�Yg���!��"�f��K���]^�k�
1J�����Q��S!���X��zj'Ŕ���5>}�U?��}7Yb�F{�IO_�[�;B�!��3D"�o7 �nU/sD�t;�@��&�� �u��u���I)�8� �-��D����PZ̼9�!��0(�)�^�?HKkk�/���"��Zo�E 
;�4F
a�t����t�F��C��Q>�	���t�[���	�ʚ������T��h{a�0&8�45V7Gk1�q�5l���������M��dj������і�r_A� �_��ؖ���OЕ��2e&��
GDlg�Oy�/�r�}��'֨��|->]9�Z0�C�yG�/��_�?�?��w�G3%1n􈲌ɬ<�)7�Ɓ�1�'˾8	A����XV����mi��gIf(%�_M��Iiq����l,��W����i%�O��`���SP�Ǭ)�s��{k,J^@=�n����5+lc��~4�t�1���+S�Q��([�s;�j���h�z|-�ǜ�w/F��[��_��J�����h+V������满�����O�Jx�_��K�+[�۠��|~��N���;v�J4��l;����,d�a�|��b�+N������$2D��&o?{2±����4�w����A�i�#�F�f��d}��	�'�(���Ũz�3K&"��KMs�]yM$�א,_=���R1�Aި�r��Z2_rj��rL��O����{QMт��zA�-.=�`Y�zvjnx��&ܫ>�7/o�LԹ�*��!t��/��a�:T]Aq�=�}���$�[���)�F��r�e�� X�����,��l��\kN�� 0���s��N���w�M�N�]6�(k�z�m�^���1�D�B��L,�Q�1�I@E༼A�N@��7�'�鶄�^ꪴ�i����Ǖ]���s�W�'��N�$7tF@6���0K5�l,�7?�o؀�sX�^"G%D��w��K��������sV-�������3�J�m�y�q�뀮c���9�F:�!��C´
�6<7Xa�)zp!S+�?0d�8��j�e�ҬF�s��ZVr�A���հ_��*���F7*����t˵��㼎Q���\��2(��2Fq�.j��n�|2)"��*2�m����a��!��]-N�m��\�ם�b]M�Ml&=`�LX�7������/��ΰ�'���$�RVF	�v\�R0�YI�:�L֫Z@�>6X����d(+Q��ߙ�#޷"�9�E7�W���E�22�L�t�1�(3�
#;�W��H~vQ��m�t��J��U���Ֆѱ�ف3����	B� ��U�1�v���������	G�W�68b��u[
hD�'��2O֨�j
�&��f���5��P��]5ɱ,�,NA���2E�X���mb��me��)^t��������)� ����]k�+S-�Oe.����,�A��#E9�H�w��/a*����p��*�?^�k���EY���B�D�53�dK��[��0r�m7oX�	en=2�/Y�t�$�?b�[��t�r��ȣ�O�ݱ��h��S�챡�6�\�EY$�&��pc�h�����X�����\��I�yX���M]Gc���x���$?�I0Za].qÆ\������Yϐ�΄h�C���ǲ)�V�8?�~�������=6�	�c�0���rԺ�;X5(}:`a�L��%V�Cʺf������~`���9@G6��# �S ˁ� 3��F��#�����U����i�����Q������t˚M�R�(��i�{ڃ ={�ϕ��?��v���Q܃n��?��xA�DM �	(�7c�Y@�z�)A#6�����y�?J� ���"Ud5ܸ������_]pX1:Je��]Ca�y���\������ɥg�v�'6����-&6ާk�sS5�&��kV���<��hGU#'I���
@�1]�I�(�6��´��J����7���咏�٢/��B��,�i�����hf��a������ҿ^�!�ن��������v���7p`��.R�J[���1�>υ��?o���܁{��@���z�-�)�OR�f���:�oǸb���bN͋��5��5Z�L��;���j�[o�����V���]���E�~�Ϲ����2(AQƉ��B���p����M�6��H�?�a,�`�i]��Nx¢�36Q�f�?H�O��d��������vWT���k�rq��vO�,ʉ��,O.���-�����3��G&]ZY�r�K4�Ao����,\)GQ�ok_����T��05}R��ҫT�G����M"J&+��~I�[�Փ����dc��Wo��uV���ʓ/Vn��������z�r��_�}��4�Es���X�&�C��o�n���#�Z�����'��3�B�nR^�{�ld3���ZN{�C@>xi@�� �t��GW�w�k=�P�[A��UvYi�S���n8�)24^�:S��j�=X�μ��9q�SS�pN"���cƀ���Bt���r�50
 EGU��F��9iϖ2MZJ�w&��|��+s��r�i��>�}�Q�~���|��So}>a�Ѳ�f�[�V��d
}������2Ym��I���u��@�c�U��OVP�6q������T}���c�U�����S�#	��x��!A݂$�B1��eդV��xJ6McRQt%�sקx�Q��<q��|�I��n߶�|�^-�<� c���!ف��?!�|�h0B]�����wu�	K�]'�����b�e�Ӈ�����rG�	��5:�=Ol�l��eV<���L=H�Y.��'9�dD�U?3����E=k�C�1h�/���㪐�"��)i����+c�.�E��2=\�`�<:����{�`8⠸C��v��������B�y�a���l�v\��d��.��t9��5&D�B�wqٌ"�K"Dw�Wq2�t��xqW��v���w�O�jA��Q�s��@�P�!#`;Hݓ���5@����X� �n�M���W��M���aNۈ�b_� $9�7��(����IKvm�n1G�E�Ƴ�_�!�ء�T^��ު����J9��iJ�ۋ������Xԃ�0 z�EZ�S�c�GĞV�`��e�	)�* "ƄN�� �������a�nKG'(8i��J֮��7Oui7~0ͣ��`0z�7�:��
 	[HWX=�9���b��A�� �B�|�3N�ӣ|e����K�F�����a+נ��n:��x������9��<�*4ڊ�AP�ǧL���J^(����{�m��#��1��	�0ٌ�s��;�'�3v�TQxt�o�q�a>�t��ՙ��P6q�E%�]�>�����;	Akex��` � )ܕ�\D�å�
��j}�	eE��ļ���p�����u��ˬ���&=�}\��fO�#� -bک���1m|a�h�Ǟ.ha�`�5�蓃�p��{[96w���6 ��� ��̢�_nk.�ܺ���$�����*�/C�)���0ls2��f:�H��p�_��68�ь-��Qu�����qL�h�:���ڀ�cB؎�Qf��~W6�qu��0��РIܿ�9�iз|e�A9LP~�-.	��sz���������T��*�w��1q�U�Ǆ�-_!L��;��̀��[�=q�����%&+Z�^�e�E�^���<D�嚷�4��5����n�q=|��4ɢ���` ���XChQ5��8{�����\[���&h
0��U���T� ��EO��ʟF��c�Qp1ˊ+���MO�A����P9���gBԷ�λ'z$]E'D�֮mb�ج��ױ%xF�=��Ł0~.e�Mr+�[6ApRG7p���a"*�.����%%�LW� ��������U2�ݒ֕�yŁOD�"��fµZ�h 'a��~[�5�� Aы�a�R����(4Q���C}�U̡Gm/�� @MS��f�z���k����	�+�Z�T���5s���+���{<��=g �E�j�5B���#y6�����01<�g98yԚ\���%����RK�̆��C�g/�Ə��cD�m�x7E,�D�*�1_ ����T��Z���� �|8�n�³�v���8�����@;��
;c�^��~�T<G�� ��]"D�=�i-��۪��[է��N` F�Vf�`�_��� C�QZ'��a��Fu�n~������6�,=<Z�R���s�%@6��'�Tb�͡�p�z?�f�"���9���r�KEQnW
y�7�J�4��5��1��%��0��c��H ��V���Y'̆յ(+@�m�kB�\7֢*�;��#9���aQy���4;\�.��lZ��t�%�V�2�u��Q�B��!��z-,�v3���ٽ��f�>
�ŌA�m�	��K3NRQy��	�ģp�Z@�i������
x��!W�T ,f!�qv²�!#���=F��-izw�/a���X��&��<���}�`���ۚj�F�s(^�N����+x��ʪ��6(ȇQ����}%$���.P�e��~��"�t&,q�&m��9�����Ց�G��s�t����s칐6Q���G�Ѽ^���Β���w�.Nt+�@*W	 � �owP�{��1!����߬F�Ĩ43)T���ӑ��������*(�+�����,>7�g w%T���}��j�vgl@�1ͦ��5�sM���ͪ���CS��x���a��g`�1�7�*��Y|&xe"*��P���j�^x�
�:.e]ل0�0����e���Z����$wy� ��}�֖���j{��'0�`R�����*h��v�3��z��\j�*S]���'R�9�^�>�<U�Fe)&�ݢa��O����ۭE��E����z��}_~��Y�_����WT­�b�	�_�����7rx�!�X"	LT��8�pjn��}��2M��S/�<FU'�r��D��J}0��w�.��4�#Ǘ�����s�E�\�`d�����{L��RҚL�Y���ȴ3�-��rpffzP�);l}�������K㼟��^=�ס��U<��h��7,D��|r^�ٍ��_Q�#�k�e=�h���u,8���ީ_&_S���32C\~�6�����T#I�Y��6�o��������77�a�m��uWH�S��KV��[�XI!g�ϕg��x��r�Ԯr�:��s���*3�_�����T�@��c���{���3���(�8!jH䑳f��!���[�b��K���I�b�%1r��;��2ڍ�*����i��N��`!��JIMќH)�^׆�_����TJu�o��m�;f��s��]�*�� `j=����)�rA�`=�&='z��b��<�_r�(
TB�%a��K�V���3��w�C��L�Y0�Ցb��;�	!<u]��Z�rI,s낲���|��ͯ�F�\= ���.R�A���磬�֔���-��v�)��
f9�|��$�6�/Ş6|ځ���:iY�rR�	��A��4����&�cW���Z����4`]i��[�{~h��ɱ���S2�R�rg�D$��g���Djɖ��L�&�J�����W�B��µhڂ���Ǧ�W��_��܆*�Ѯ{�F@81\n:�r˜W�o���C>.��������Nt�95�r�����d&�2y��_HVV��ު�)'���w��:�Xu�����-�����:��[%�߽�x�Ӹ�(m���m�p�i+y��o�ue�b��2^u{�$��/F�.��?!7_��֗���*.%�ֱ�×�#y^���X��T��{|����tncO�j3wR�Gȵ���Ur���g�ndѱ�fc��RL!�RX�C�ZQ��a+��4�Tj�����P�/����$q��k���u-]�a,�H�{Q�
Ð�DY�&L��Wu$���m���i��ʡ&i���$�E�$�(*I;��N��ێE" ��T�>�d�}���,��:���dRG�C����"��3{P<.~�2̛�<0qC�p����An����Gh�C[#���>���葞�w�f����C4%�R[+B���`G�.X�f�L�}JS�\����x���Z_�Nr����S��\����C@捞���#5'@���Q��l�$�+]皳e�Sϭ<d����!~ G��Dh��|ϴ\g���O�2��Qj�`jUObhA�W�Ɨ��:��k	=�(*@��á~��y$�7H��E�[>A�����5�1�MX�vF�[�9b��:,��x4�aVC�Ih����@G:)�Mt��>���'>�������q� 0F{���n�5�~�w�[$�d�`GoU(ggt��8�����B�\��^��%K�R�>����|��\P�{.y���1���,*����#Pnp��6�`k� $��~�Z���ůo�܅|�
�8��_^#�����x6e3�<!nu[��9˱�m
�m#��ᨼ�1]����MK���a��6����/��[�B�����)r�Ԟ�;|�0N!L���qW|.4�'�?tG�K�I�{����o�s/::#�(Թ�\��y���.��v^�y�M��P#���1��Y]9`�#�&_����X��xD7U����h����n���I)|�Q��k������%sYMٓ�c�`i
���jcN�����@SU��<2�Y�8�X����8U��XC'A���u��f.�8��Hܧ}�+�(h��-�9����+��]~00I��s=�_�����UF�+ Qa	=���Z���CJv��MO��6F�<�(\��岎	\�di�'�c�=��Of��>��@H��o�@&����0�y�as^����\/r/q�b���>!������VDH�$Q�@�HUK-���C;�,B�_J�D��<�;�`@$ 7�f�v�y����j�]-�gfn��Mᒯ��� �S�����U!����߮�(cJ.�}�3�uUfG���QӤG���%�Hv�����X�-���D������dk�܉T1H=�k��tTL-�T�V���_�6J�g1�#�q!B�Vr��]J#���86c��J]5��R�>�䨳 _���T� {وL��H���7���
�{> x�(�'������ڍWg���f��#B���E��~|lHD7e=���_�� Q��ϖ��Jn�i*�܈��5B<�� �g6Y#�Y��J4Yd�=]���~�TC*�ºk��'|���.��'MH�RY���4w�	gk�?l�mB���A�@TTg����W^9Ke�ҵ2�~j~!��? �?H��i)��a.����y�V��TUU�Ԝ��/u�Udp��<�9��>V�ߒP�5>J���߰ʚ��Ԍk��)�_w�k�5��Y*���Px]�?��k��pC೜�+��d$�;�<!{�f� 4o\��w˰�Y`NXP�ZG�m�ٿ_�#B]��  �M�N������-/)�Z�Ǆdg�9
�b�D�4;c@�>���_��'�;�9���7��F�ͩ��YD�s��B�a]�Q�إ�U�A���Τ`P��
X8B��D�ƖQ����v��C�6�T�T��ՠ>hg'�KМ�\�q��a�B�`?nY������~O���	ڲt?#8/�A����<b7&�!����5����ͣ�_���%�y�ϥ�b�2Y��lamr=I	��续ע��'�����H� �$~��`��m��l��������6��7����`�)-�$&���f��X-]�%�1�	�G�c�qn2�y�ϫ��v_7>��8{����B����SPN�K(oL����{F�2m�b�3��x�cE��I��/��1��C����a��m�V��7�>-��Q�R�,s_�d̴�6�")�ZsA���!oJӇ.��鿧���^O��̈ v�D������3l;��>݂���v_V
�TrXC�m4�ni2������h69�I�֛ݘF�c��>�� h�1-������*�I�}��0���7��p	��(�I��3�0��X)^�=PJ�o<��D�
�_gLD"��I[��Q3!�[PHJ=ٗ����7�͟��mb�/C��ZRX���l��@�-�$��2C��f��fZ4&-�!d���X����?�f����R�����b��O�L�TE?d:�� 4���|�߽V]L��ć�j&����\rs%	��:'D�Ya�6��W������˘������%"YR�`G���N����^��9XT�%k�� 3���\ L-�X2����$��t�ګ�����`Sջ���VLIn	A	I�ld
�x?CpG��2#�Բ��6� R,��(ߕLTek#7[�Iq�L�yKHMF8�#:4
���7��m�I��5�w �S����Ʉ��/O�ڷ�ist�X����рX��f˜Z�+<#��>sA�Z��ʂ�n2Y&�Z�$�Fq�yh���ƒ��b̧X�+��~�Z��	�*����-�:+�\Ҫ���R��-��^0�@�m�q���q�y_�]/�'Ϊ��*qI���Yl :m�����[0�{�]�A�6H��XX�f/M(���Q�.��Qb�L�4�ޠ?y�A/Z��^�5���GG��k�j�$Λ�*���?���qt��/�������SPe�������sR%�. wu��t<z� �a���U&�꽍��v}�ޢ�n�J~i�i�ݥ�#�3�w�P2 =��2�X��H���
pg�v�5x_����ZQ 0�%�4ztyD9|m��EvJa/�/S��.�q(P��R w2N'@�6�n��^�%������}�YXqf���ڽ�-y�I�R��9kXf��)�v�,�qñ\�0��*�!�D��\�� ]�"$������a�O�u����!��&�N��y}�/�T#�5���=��,�^�t�Lg�j�s�,�OFh����7�N92�K���u����c��3���A�_�j�I���p�b-���l.S8����ë 7�q�%���۩�<Ū�i0-��
�`L^
��~3��fKvqP�{t���<�mv�;a'����Kˡ]V��{�M�>�L��'�V�p�a�sٌ����`���IF�_�����Fo.�X�	��{iA�@`2h��T�
�5n	�hw��k�l�A�ޢt(<��f� �5c�1P�3�}r	��8��o`�z&qP�0�
�[���*�-���^N�J����R�D��gH������=�G��)�ItF[��K��xR�e�u
˭�9��L��:P<::p��y;0��Ն_ˡX[�5#[��pJ#�9��}�B%�1] �C��ħ���7zT?�]B�vD���(������k�����3�/P�WjO�����=�>e��`4���X:��J�G��B�9���k��}�2}�њY�P��U�/�%���jC��5�z���yvI��A�]��E��gp9l�f�X��q@���VՍ>��;$�F૿a.��f��D\H�3&{���i`0�&�;^����[1��#� $�2�gK�f|Q���� [�[>y�q�#>3W���L����*\.�9qk��aǇۊ_x��S�I���V�V�ff�$4Tfop�0�0Rj�N �$X.���N���ϝżxe2���:F����Jh_O�?�^v)�+����^4�0>	N����T!�G����rp5
o$⹭�G�� �}?X���NK��e�<���CӘE����TVf�6/L�M�9L��W�����x��_t����z�߹��O&ߵp}YE���4�w��5�ߍ�o�,��H�3Qw���,pnO�=a�51O!���q�L�V�@�H�Ol��э�a����&�A���;ٞ�6���A����-`&��,�0`���M�L��0-�I�)㏻��B��P����iv�#�]˙�8���KƬ�k�y�Tȇ�S*�k����y�ғ�9>0�S���~^s���<}�6UK�Z�ݰeP�
�m�i3x��/2�aښ�Ԍu�4(u^�c)��!�6jU��Sqo�|n�WK�x��J�󮽥���Q�*TÙKiɲzJ�u�B�B��J�r������g��Y�uq���'P�o^���+Z�z���J�	Cy�j�HD۠����q^�o�+�#��e��rdL�̯o	��O=*�Sd^�M"Y�8�&Q<."�Ѡ�� 	��)Ҟ<��gҘ�����+�~$��A�x�e�;�&�Q�Ak/v�w��:��-/5w��N�z��@���3#)D��^hf���\3?�� ���ZG��ǎ�pV�fe�P�P��Ys��u*�r���d��V	� 5uo����u�����喾H��nAA����qJ��� ��c��o�,�5�)9D��}¯��a*CͶ ��WL qq�b�-���x�6��@��������i��Oc�y$/L�y�b��{Au;�y5P��:��\�O9 �-��^|��9�V'����e�4�oL",�T���ֹquk�<=E<c�ȇ�N�n07���M)�M��ݷ�LS����*��VO���<�֢�i>�v�q2B�R�)����:����4/�	��	<ȷ��g�]��)�7�a�wE�k���B	2��][-=�뾟�k�8a�4��ɵ�>�4hNm�������9��̞B�F��[,��ݖ���宱D�lgK�E�nd#�*tyTo�f�@��\��Y������,~�IM)PҜ�'v0.� �ĉ�� ����Z/���e�����(��ⱒ�$�?�ھ��/x��sP�^�(�Z�I�ٓ�w���T���~�p����z���m�:IKm���b��E�)7��tN�Jf�ZD���)�w��	���¼ n)��.�B]��%!��۽G�J�����{Te j���׬�p�4�Sb��;��m:O{�b�v����k�u�������	B��|�_vT􈎂����P��
�	����ޒ?Nc <�f����{�R�+(���hm�ۼ·�ٟ0�b? ��}G�,\��Z=L�eVq���'z(Y�U9�6i-�j6?uas@�8����d�$�-���D1Gsmݓx�:P��/�������9}~}�q��~�����`.�6�wu$2R^�@�lH=���B�Y�i���Z�o���|�c��NɁ��؝�����H�'Bu�$螉��E�����~���حc�&����qj�;b?Y8��v "=��J��2�pe��T*�U�"��dT�[ul��tUж�PbO��u����.��D��3Wkb�ї�{�m8�����K�g�3<���7N�J�����?M/�w�I�s��N�Y|�!�Af��{f`h>�Q�(ٗ�0���Hv�O�+��%եuZ kk�?�;�#���j�m��������\�}�O��m��CE.y��:A3������XK�+C��/��Y`p��Y���/��WR_��ٻ~
�1�5\�(���)�Uɓ�I�����U�SZ�� ,#���N��-���fN��Q +��e�̮���0�<]@�#�c.9@/i����]O�F�p��и���"��痡�&�_znx]v>��l��Q����Ѷ'��Rrdz��@�(��}�<�$ǖFO��7����8�	0�2�����Zn���D���=�uՐpp����8.�q�>0�N�U5<��ǩ��L�P�
epEm�vJ+(V �W�H,��*4!�
�iĵ�����=�+��W	��J�bP1{;D=�ct��~j�����d�ӄ|�ǯ��\7+Cz,ɕm	-Yd�<^*��w�����h��>4:Tq��i��"�"�����F��$��a܊f_r�1� M�ۘB��Ц��/h�~���:R��l[�:m����<V�oH;o� �P�FRU _��G�#�
�Eg��f�8_�x�n� �F����_�����H�)�[��ᒔD@��>|�S��kD(D�Po�d'��c-y��$�^�8>U�$��v����O4��6���㊗n�ܜ���0�\$�Kmw��h�)RM��� b����g�L|O57���ޖ��j�~�q_����+0K��e���>�B��+��a��uH��	�V�������R�ýX����>{������G�p��	�2�g)�n���#{x,*��B�����IW��A���sΔ-�r����'���P������
�ڡ����v��x\}�q]�MV�y�y�#�ћ���'>���晄�k�h+EǷ�q�m`:qR��r<�{+z��(��I)��:���H����io��������I��uC*b�d�li��g��ćKho��yp�ut�G,�h5�ɷot�����&��$T���
�,a��)�����|3��?[�-���f�n2�y�]������y�@z�U>���Z�Z&.)D��e��vP~�яq��<��u��3&F��?t�D��Oh��V�:���>�!��?Wޛ����D_�]�M���2�qݟJ��U����Q0�T7{�IF��N�ue�Me�^fGO��D�"EKб���fY�F�0k��QwF�(���mɦ90��Y1�y� �z[�,������Ѣw��l��
���?K�j�E�q��E!4�ϸ��52d�h�00B���UNħ�rXl�o/B[�t1�����%�?S��C�У=�	7��S7�S�0�^c���x9̷�2DE��5t��;�˪>�����Oԭ[�wT�5�j�j�����+9�n�#�j����{XS���aU*��:8����"X���#y��he7�,��$�E�Ք��	)� �"�A�ڗ��)8LtB��*[0� &NAm=���!�"7��_4B���-��-m�����Se����n��9�Y�X%r��;L�7;�x�	� b��I�i�?RO�^�Ǝ�
��n��&#_�7��ia޶܅�3_�X��]n�m�I�c��]��B��)]~Rj��]��T<��RnE�cw��k� Ub����l[����#t�Q"D*00��W=F�+��XM�a8���1��N�!$x�1��]k�_oj�x����Z\���[>�`0;&RDEĢ���ݖ������\�D�V(��;��]���Smͮ�T�~S�+�i_�<��,���cjM4��$ 6�0���sd�_��z��O}*���%ڸ��>|�<����bsh�*M���G�"��X������e�]�֤���b��[�bAz��Y7��b9�P�'F.�����w}������}�|����K� ��_ر�!�=�f��%Eo_E���,�n�~��)i��޲�J����Db_��&��s3�@����<2u%�P�3�0x��{�PZ�Ɡi�K<2/1���-� s�����z�p�T)��РdWR�RRo,���p�������_ߌo�g�jN\��1��C��+����d2)���hWۂ����y��9�yXeH�=6"����Y���cß"���M�bd>�
�[&j��nN�����9Z6&0��� �Fjk�f���a?(���t[�@c�s]CHa�'���C�FIf�
^���C��u���zW�0>#�f�W�;��;d����Sr�hÊ�,��fY�E��.o:�M��UGW?N�L�L��>�:��i>�j�q 6Y��e�'\���3�[(7�e����zd�a��v�2L�e��~D֌lZω|�n������7/9w�|�g���ی	&��^F��]���`>׈狭J3���/2Ap��g?=��0'�Ԇ<��J�O��fC������o��T�l�	�1$���銷S��A`�aSyX�J%��1%Ȥ�������}�X��o
����31^:�=�t��#�������!q�4۰�2_/���C���f�6l7�TZ�27�ܖ���I�-0�v0�Y#���&���u���Q�[���ڦK�F ٢\>��4	���# XÆ`�u�=���S��XSO�<�t���P1U��	��
��-�|i�3���Q���M�;,�	�����p��*��������,��z��4���pf��!��=�A�(���GVFQ�q?�ު�)]��v.�#3���4���s�{[9V�-5ys���y�=c0�\�tX���Y�x�S�N?�CU�>r R:�3�ŀ�}0C�t�b���f�-��JR\��F��1���B1��+S..K%��ٖ�Āʼ�Cc���tb�cu\b�3�v��c|��G��/�C"��+���8�,˃�$�ϭ"t_�����>v4�������J�������a�$o����@~�$c�����̈́�^B�7φz�̥��P2�P��) ,��R�5�!�Ջ����C���j����ҔeK����]H��]f�^ݧ*Y�PDԐ�
�Fb:���Py�e�Ϡ(��!������x����W*���(��S|�X��T��*���,��{jʝ�a�B,�.pq'�!��m}�<�V���~��2�qC)R�v߆��@3o�R��\��gF��S�z��١I��@�X|UI�Y��<5���G"��]$g���"3Х�  ��z��N��	��	�����)!�V�"�w�Hר�~-k�M���F(p�<�y��;I��m>�O-��mc4�,:7�_ȬA	^+yb�,�K�{��2[�L�^�{��K��'R�"�ijֱ\��$���,G���[�V��m�����J���0qX�ח鏣����o��'*���S�f𜰊�N�SK������˗ ���Z׎<���E(/[�s���Ω��Ca*��ɡ�F��z������d)Y�
N:�ч���x8�B'���"oVz^�$��ຬi�Z���xf�I�­����YB�<��{F�{�J&��d�yv������8IK�D��i=��BC:Q�[4@�.����}Q�%c�ձ��VQ��M��Ų˂;V_��j1P�["ew4'�6�� nA��Z��!<%r�\ˇ�he. &	��2��M��fj�����
��r���^�1$��gMe�@��6�/b�<!j1X#�P>.x��p��׸�	AGN�"�XǶ��1� �A<w�5:�R���ia@b�<���lX�L�$={�zCsK�0-}v�;�,4�y��+r�h��֑/-�7�v�M'��#���0oP�3�%:�+��>m�B+IY�wh�p�Q�u�J^~_\��s��ui!в�K�n��M/�[Ƿ��j�ċ��[�yg(i6�S�72۵�ΰ�v�n���MŹ�/�%k�3.1b������/V��g�Ʀ�^�i;sj"`p�3��A�������b�!~K��?#{�`�	I}�S�A�I�#��E���h:O/ˬ��*jBv�@��^��o�.	����;�kx���k~G����)Ƽ���9�M�'$"��z��K�t�C���]|=&�h�A�ޙ$��ݛ�L��C:��U}:$*���B�j���F��u��&���ZU�1�1�]�"�(&\c���&��s�S�|����6�g��#�\��ݕ���@Q�:fa�Z����lV���A-�Ô�`R�=��l�����k�d�}>aFu���$` �"=$:���};�9LǺ�x�0��w5�`��	�B�8I-��D��@��\����t����{����U�C������t��7�]���� [X�1��{��	pE�W�q& �/˝����#�'H��eJV���A�EC/�զ�]�4�o���� �SB�zj���I��`��q��j�� �J�4?��IDC[� Ϧ�n��k$.W��69f)��v�����61Uk�dS���5��]J��9�ޫ�!O[ެ[W�f(}}
� \v۴�X��@`kmm0��e��a+�}�x"N�_S/����DSuq�?��=���oM�L	�c��5�X+�Xך'�yQy�s����S`������Lj�ĩi�oIt�G6iyQ�7�8Yn�J17�����=}�M�n����e3��X�l���XCW��s�ؿ�4��ka���3t�ܕ�[@�%`��OΪ�{��Nߣ�_!#sa 8Q�s�$��9"<��~P��Y��3�M���~e��T��le���]�$������!P9�S�]�M��q��9�'X�R*#m~��+O�6dx���d��#�M4�����!��\�ͥ�@8�A�I�؃������zS?<�-0���l��_�9�~��c3M���K|+:�� sc�Hz]��}q3�N�V�4W"�c���(	x�_@>���04\�}����J�F��^��j��Sٍ��N��_OХ4�.���e�CN��� ���k���Uj.�����g -��n�둆u�oX�5��Lt��/i�D��O%'�Ȑ�y�@C+�<8_O:ν���6��%����Iw�'a�*о�������1��ro����(w�iٻ�M��S�Vq��B1F0�~q��a�����9�w9�<���2��ITc\�_2ӂWr湙n�[`���h��Dr$�9��
�)�W�A��Qbj�P)���k$�JQ���K��R��P���r=��N�t�%�o~��c�pBf'C�ݖw-��A-�F(����}��z�P��z�\�s�- 4�2�rB�� ௤T�%�	�?aS�O�\�<$eT�ϵq��`������u�4�d��u!�]ͨ��>�T����"�������B���
?h���]0v3��<@T�đˌ���Z�a����^�ǌB�]�XcB��+.>���y7������I��r�����ad����Oh���uj_!��_�'	��5!�8��Q�q��Z�?38��eTP7�Ŵ���G���Ԟ�n���"m"1���G�!����	�YdL�y���W̿��{4L����f�g>��l�m�����{�R�#'��~��ub�uݲ?RɳE�%C�E��o4z)��8�V#`�&ɺҘq�	�i��~��u��4�m��ۯ�%ec���9n�j=j�B�$�Τ�g��Qì$����t�7^�<A���-%=�����~n:/��S���r�~���R�n`$��k�-�@b���$j��[gF�R���x~o�S!�\6g��������C�)5��݉�]�n��F�(�2Dfcr��n&)6+�Z`��6O�(�����b<N��F�k#�x#+h#��_�L��������T���n}djUٔ.��쟸ωyM_��W=�>�}��X� H[ŝ�A�>G�v��SH''`v�q!�9����U���bL�):pz�X�v5��W�d��')Q�g����^�\��+ ˊ�nf5R��|��:���Ŭ���0��L�\����K�p�Q�'������l�mx�	�(5�I������/�[^C��S+S����0���ª�
�]A�,F�m���5�K��jX�u\-���V���d�����C��Q�avkO,X5'�Kd�A_���AN��#���7�N�K���b�kÈ���4�w�����P8�Eٟ��g;��µ�E}�ǖ�N����%_ބ�g8��1��|)=�>�p�լ��q���q��r�Ġɗ'p�Hl��.����E�<K��c�}��%Q���J�f���~aO�� �j�tRRF,�ѿz,-=��0��;�]P!�5q��]�E(���Wc޳_���Ҥ�kg~�+�n���hE��IN�T��O�j��!�H`Tv�C��7�y�����t6}�>��y Uy��X.�>�`�ʹ�����wy����ސ�w|X_(�Vd��1_?WԲ=9�ΚԘ}�R�OH��t �/gҗ-C�Og�9	,&P��1��[o��;����h��#�$y0��4;�"V�r��Z���+Y�B�B��s�>�� �U�'1'�~>��q"{@~*�6��+?y����1K)��c�5a�GN����&ɫ;v�Ѻ4q K��l�]L�+�c
^���=
��O�8g��[�~Q��v3��L�OGP9P�-;�z����+0�X?��@aK.��P�����U����4�>����p�/�����e\����F��8�x7�%uE����k������KdU�z��s�O�eX)\ik��;�������_�M�h��T
�	{��ݛ]�&p�U�rj�$&;��2�: |���y����u)F��T<@ՏW�T|�祸Mw����k�B�ό%������5��ճ����j=CD�(��YPU����I��_����a�ǘ^hy����H�{���P �$ZT�qb�.l���[��5�4q`]ni0��42�$�Gt
�WS,-uB:/)<�!>�����-����a�I�A6r��ʫ��L�nq&@�����<���Z��=`�-n1�-��9E"n&iH�]љ $`���$�|���A8�)��8��h=p��{�CI��7|	~�U�.FC�Ag(w��D���`\wr	�^u �#�QJ���jʳ�RBGU�2厈U���#�m���#�$R��2�z*�I��M��A�_|2*e�;؄T�ǭ"@6['�4N��Eiؾ팷v�����-���7���|eYb��[��-M��&
&�F�z	��0JNI�!�����[AXs��Cõ#��v~�������R<`��ki2k�"xp[?lC��O�/z�C� ���Ѐ�����w}o���v`���D��YB�B�e�iL!G(E6_Y�7�ܰ�[Q
��Ե�/^�����R��&;_K�Ժ�}H��I����Q(�g��-�t�G���>�τ .�W��e�^�C�6���=�|���~�������ωE�'�A�c�^�O�G}l����N/
H����3�jsd˿B?�?��n �����)Z`���Q���l
��+��V7!�q-�j Y�j�i�3�����u7�R�4&l�;��I��6jBޣl��S��2�B��Z�k����zY�0�����>1��S�8��]�g+�ƥt�꽢��&L�AEk��)���0J}����+5��@�ǡ�=�wV�~N��gv	Q~����Sf3k!\B8W�bIP��eM�M��T8_�;�m���Z=B�G��V5����'��k��l\i��vC��v񟱘&CD�Ĺ�H�J��g���N�2���`��ʧ�,į��}lbЁh��$?kJ3 �t�,���/�7 i�-	�������U���nB��܍�V��:��yN�3z������b� ��X9��D��4q�� S&�Q������\Z�c#���h<�������A�ҥ\c�c$�� r���b�K�v�b�|n�( ��;�y�3���M.<��$N�Ӗ��N�dyB��4���.�r����Ի����`��	�qt\�]�N���P]h�W�P�c��nz{�40�dάq2ۃXD0�p��eǅ$"w<& ��D7�#���he��qȴ0���iM�o�N�EH�?�F��z��2�(�L
����5�^�>S�C��s��}��H7�G՗Brm�Q�ۛ��<�Hj��37#�����s�o�� �M���-<^ԙ�B�(i��2Q!�n��m���V�I���}�=��A��Ie_I��A@}_��@��|���z.���S� �3#"��ܐ4�S�]l/�� q��M��@���$>i�.P$�.TC��Ȱ�ҥ?X�G�big���,� vY����a�26+S���E]��ܗ@D���9f�i��).�su��8X�S�|3۬��8�ק���t��G�Oc4����n���X��u�4gF5u�p� �d����d��do	%EKO�b/�xR����}'�y����7��{�n���ǣ��Ă���S@��/�)���=|�������@��T�4���bnJǌ�����
-�,Ǫ�뒠���/4ּ��D�Ə�!�D3hC�M�� [�߫Ψ��`~��"rZSbE�C�|3�Iq�}'�z�SzH��).�;��3��Ts`�b9��� �.<�x���#d���fd�r%Oڅ��Bκq�L��1��;d60z�D��}��8�a�I�7�Y5�9���d��B�����B~F�nqI.+��<@�l�Mц�L���i-�(�+���D0����k��1�XDyS������u�%J�ӫ��p�op�^��t2.:�∼Ǜ� ��`�[����1��zpH�������"���㼱���M?B!?#���P�T	1|��%"kU%��Tדt��e�J���-	�Q䍒p�Gʺ$����E2���7*[�+NP��9Kh�A��09\Y���� ��j���K2H��r �f�;�!����KR8��@a
b<��9�+���=�o��&���pU��c���abeE+=�����;t�+G6Ӓ�ڮ���n̬��^���l�N�;Q�{�����4�DJhM� y�s�������B�V�p��0���f�d��� �;��4?S�씻����'����Sa������J T�߿H-+��ӅZe4�Rl��	��R�� �[�x;р�x/�i�ZY�&Vl验Kt~/hآ�z��N�B)p!%�>0?M���_�핡�1�(l�z	V���Z�N�%X�H0�|Y��{`b��}g`�c��'�Qh��[���.��ZV��l���jҌ�P��3�Fl��Mڈ [���Ca��`1X�+���:�Z�r>��φ(�/%*Ҽ$�^0��������`��z^�	³���j���2��P-̱�)S��N���#�qn"BՂߠ�
mB���U�'�՛-!���0���r�Q�N�᠉�W�	dJ8�ɲ5�nLdJ�������8��v�$�Y�"�kр��gw�:�C��$V��mJU�����MKo�	]�e^��o�g�t_�����=T�ފ�vW\ֶɎ9hi��,dŹ���o��'���n�t���&���΀�G�.tͦ��g�z+|��y$(E�s�9Տ�JXɔ<V�!Z��r��]s�f���{�(�"C�kt��s+������{m,7�p�uB~��i�qU]n�'�����:��s,���/��¨���l�\ �q6	amH�W�G��`B�ۈ�r +��ȋڽ�C�R��U^�1��?i,�uj��aZ�D@ab��rz���9QW�K��h1��y�\�"`��4*�n�#J���Ǩ�F�rGm&�?�˴Ǻ���w.�|�Ť���ʍ&��ÕB�a�d�t2����?�*��$V���D�����;O�x@���D/�^M3��R����v�h�T1�鑪���* ^��.n�5@�M�� �L�d����T��\�W^%˱�4��:��/�8�F��V��U�˚��+�v�Y��0�$���,��ree�0g�}��/"�
�Lۄ�5r�A=GV�?�տm�9[ͨ�[�Mو)�KW�n�Y�OO�z�Ɏ��>	@�T%�A��W���5��	w��.�@y�=�t�C��T_��}*��a�Z��F�9�p��M%Q�H�mIV�~6�����h�a&l��8l��䳊8Ib*�c�0��K7u�-W�����7Sۮߐ�n�@�.��BGjQF�]�B�����d	��i��R�xB��w�`��W2s��]��U	Jj��RMÿq˼���l�V�����S9&̷M��[@�S](h�M�U��&i�4��ikY�a��S���2A�OA��@��Ʉ�8�f-����d'������2�`ʁN�p��$=��ӂxs;���-���
(�9�L��OxB_���
��4Tt�3�,<��v@l'�F

��Ɨ���
��d	%��!�m�,�e����V:�Ѱ�ۯ[`�����"%��������$�j��)����D����X(�S�&!C�B�H_�&:���Ў��.�h/��a��⏼of���OT��Hd�"y!�m9vU� ��I�L��ۮ˵˪�\
a�]�S<� �P ����/�Y��{�ْR��v|^^%����B�b��Y%~�'�/�͠��0J��A��b˽��+XX�BE�3/�L@෫^�r����t�@V�uMx=�U"�,�N	�w���'���D9���TC����W�Ț�|׷g���,�}�U��#<ه!����)h��F.4����\��uM�3���U-�АH>�9`��I�<O΁,_fH���פ���p|
Nf�eN<�"�=��n�J�`�8�,j�j�^@���b���p!�6��ⷿW��kT�U�P���'?����	~�UKj�\�Ҹ�!R���8pl���~ �R��E�LƛS'y�#1ʞB�Ha4�7��p�@��$�	B3	=LY��2J��U�FQu����.k3o��se߃A)���5��V���g��&�~��LQ�����!xX��o��O�w�=m!�F<�~�A?��G��X@��l�5VA4w���Ա��#��gS�Ea�oo�J�-���i\]�F�uرz?c|�>6Zr�>�T8��r+ڛ�U�POė�|�]�����YGh��~���Т�;/��:�C�"�� �"6@Cz�� Ώ��4���ߊ��>�n�˅X�^�#5t�}�dg"QR�;.���n�6�>]Ӆ2��1���w�����y��0����֊�v�oc=�ɿ� �����Z�G��K%�OH<b������i)�7Gl�ƍ�NصW�%l,�K)IN�(��bN�-�ۇ�=�8��i����	4���e]�p6萊4v _��B��$x�����?���Wa��0r��7��.h����xM�Csg��h��A�|�7��t?N�ㄞ:�p���9eX��QVv~��(R��T f-�������hdK�|?ߊ��E ��vRL����M�>�/,�=��@L�|�82$J&/�������7�hP�EPZ5���آS��r\�Ȑ#�ݏ]�b���I���&��
V�]҄�����1K�SV��/�_���[x�O� �݂ X�n�c)7.�M���Ru���'��q�], ܮ,
�R����ѓ��^-���=I��G��o=�����wD1>Gs�Y����З�����}��}���HX�1T�M�%?$}o3G�dĢ��\��cR�̖-,�Ր���j�F3`!��G�;�c��	4t� g% �^c��%bԔ�S�\e��W�r����9Y~\yHN��.����8���-.��wA���9�\�Zޣ[R����V�J���WE ���q��n1�<��QS���+I>��]�r��u�ݾ�;��s�
"$`^t��p�� 1�Бº�� }Fi��Z�����f�����޵(��/[Y�����6Z�O`�æ�Y:�VF��}����&_E��F
N���a�/�r+��Hi�fD��\~Xy+�kWI��k.��o��8��J:���[>6�RMG1h@	�����s�����N���~��|q�ɜ
�ރwPS�4���:#a�NЈ�d?%�eZ��t+'�H#�ю43R��n��I�,`�Yr�{E����	�Q�U���y�	
l�o)�d���x� V,�̳\�'�a���9�w@�����Wb̏���Mr��ʹ8�h��}�=���U�F0R�6H親�-B�8je�n��ӨhIpr@?ϏEV?"d�˵/雂1���ky�HǆE�q	@�@';����p�L�������2����5Cz�pz�˝���X�4]�j�-{h��	7h�i�^>�QY��P��lLs.����ϫ���J}ڞY�����u0�bF4>��n~�k��λ-��f�������0q����0���j�8�v����:��6��{������n���a�v�qn���~(ʹ�~%}�B][OW'����[��j��=��g��͘9�̈́%�V�L��^)+��;�������#�.O����~k���tTף@�=�#�����5���r0�(�W�G�n0Q�9V����T�|f�-ڛ����Ղ�z���ia���X�CFo$a��y�s�Mǁ)�س�������=m��N�@�Wf��G@ݿ2���tB�L{��;B�A{��9(*&4��vi*O�?����	�~�	�����7f%R*H\kd�*�u@�
�wgO���o�r���ђmٖ��,�NI�q���vg4�fu(��AdR�Ct���9��f{�'��w���o��W��"��͙D���G�>���	|@a!�����փ���ܮk0�_��b��hc�\hĚ�9^�9m]��C�7BY��8�i蒘��zP�h�,'���q��7������vT���r�z�}���t�hM�L�y{i`@I��=�3���>�F�&�	��v�4R�w�˂�q�;O��96ת� ���L��>�+�5Z'|��MaI�0���q_�xڡ.�n�]@Z������6��'��p �hdf[Lk�>��7̋��gs1пp�M[oڀ�/J��r] >ڪ�f'z�*��d]�H����ѝttdĖysIO&6��4�4Bf�Ik�_�Me"P���R�ˤ�;��^DT�a�7�!��8�xY;T��jw**����I�g!4��x|�q(��<��1ه�nUe�Ԣ�Mĥ�K{l`DE @����*^��F���5 K�=�
�#��4i���I<({6���\I쫳X�����%`���Q�5�0��������6��j��.%�8v�y�b��ƚ\��r�U|,ƙ��#m� �{���b�G��I������z���g�F�t��)&bd΅�m���q�7Α�s��T�	By���W�A�W��ʆ�"�0ۢ��E�6�YAv��ܪ�QKrE�sb��JY`����_Wzcn�l�nP?�v�����}%�l3��������x
�L
^QN{$LKbsP�Ia淚�Tv��4���c�[�K��v���أ�?��CK|ڠ���� ��{�� �oh���.n���ƒ���(�]G�6�xѹ�[΋�Cn��`�s + \?$�Ecc��f�_+^����p�hj�~��S,�i�h����<:~�>W�m��@	C�z 5c���>�xtf��մ��C�,�4����+	H�����+���(�t�b���=�U�eI��t��5��������P�\[6G1��i\��%8���?+�7)����{������C�.[*�^>.�Ӛ��jLp��Gm�.�!�s���2,��Da��dS��ϭR��#���jE��N\�����̇k`�k
 3
S$p�ݖ��`�C������P�49�>Q��+����M�
�ty�H�����sE�QAY��uv.���Ć����_f�<%�`4B4O�g"î�kU*�Op:<��X��延c-�>��{�)H�:���
��0�vN���3Wr�)B����8Pb��o�7���{l��x��]���(gbʁ��/"��󌜔3p#A�K`�4�3��]5��`���ұE�r������Ԩ�
`��䗿�ә���7������D����f>�I+�k�k�&���Cr)q�!��ٛ�/ϸ��vV����g?el��'W�e�2��0'>d.#� �3���L�<�4p�]�+~�A��q�A�*]!]T�t��m����lNZ��x��\ٗZU6E�\�l�����l�"p�L|L;�A�*��ٰ�N�:��Pµ	qt;���������ɝ��R.q�k�
��N2ò*�_0T�Tl�L@�a�U&-�z.L�19�����s{T�B�G��+�(�0�5�g�P�>�쨡�W��*A� ���0M��M̵���ڶ|��i�V0����#�P��*V�}�;&]�"wN _��mUS�,�	I�p�����h4�O#ρȖpvW&kJ#M�@Q�.�񷳺��g���o�b��!�`(wa.�M�I_&�1֚jx���&Ř�Ǽm]��1����B��P�`2�y �ώw@�y�rxE��w�U�Lw�i(����6��Y��7ނ3�Dm��?��ڶf��H~���"�ݑܭt	��ID�]��A��Z�7�1�J�s�����Ҝ�O���I���wݴ�=�r�t��qI���0�'v�����UY�7;��Y�/�+%
��oa��`:���G�]�N��"T�p�i�%�����1�<u~O�$<yȸ\���aœ�3󲰲C+*L����1�⢕�?��%�X��bP�����g)�&��8�$Sw6s^H@�~���3b5���O�Ek@��Ux���ڤ��&;�N{×�{N�٬���eg���, )�o @|=Qܭ��J���6�4�5!EQ���_u�{6�x9��.dqr!���7 ��]"��N���y�}$�Sm{�@P���m��+�P}Trc��ٍv�M��lpӓT��}���ݗ9�ߢ��% ����JH:�^-��������o�˰OXo&��[R}��d�
s��A"�+.&��y��P��#O�as�Ǫ�/�ӄ�z�=gN-ڜ5�����imD��*>���ԩф����ޟjf0����������LK!OI��ņ�ϕUM��Ǐ�R��3{y2#I �r*kZ���>�K~.���	�%�k�_�������᝘�#�X��>���#�,�:�/��-���W���f*�a꡼��+�c7�SB/������4�v}y���|�����w��\H꺉�]�@�*���0�V�ޗ�� �kv��O:cS�E.�K��c�#zIt'^�}'6����aH0�#f;6p���:��
@u��$�T�����
gei�B��OOn���8���+�c�@��*�iI��q����7�t6e�T�W�A�/���;y�G��8����ǚo�������j���*='s�k7�
�G�{p��-��$y	�"x<�#D]{7����:���C�r9�u�"�^�5��37z5�G��eTy���(����Nͼ�e� ��i����oN�t+$�xIѶ�����oT���Q�[��y4}�(PG-�H7��>{���42h(���lPޜ7F4Rԯ�W�������yL}M_���� wX%�wV��60\�%YE4h˪��`��Z����r�BӕF�#8�P Z�o�b��	PP(��Gx�����r��:,�l�2M_��R��F�FC��(�hn|	�|��˴e�jOD��8����eܥ�ꑇ�k`]|z���E��=y{9��G��w�/n� 6PY黨�?7�����]��Ë�FL|tJ�8����GT����3G��Lk�*X�Wc�"�%^��b��n�@L_2+p�!���]2lw��Wy�|�΀K}����J'v_
G�-O�~~������(du�:�be\�6���_�Jd�H�v�оhYX��܀r"g֊,Xs�B�'�S-����I�l�~m�xN���*4���'����e_3�ks�Ѽ�*H6)���&^�%6~i��l��i:�I6��%0dV�i쑉�˯�?����#&���޺���3���9��G@Z�2G���/Q�|B��0���5����A�]o^�3�O�O���p	��]B��l�[��CeNx%�Yq11�28�";P	�f�[�V�:R�qy���B{�ţ���)��U�9׹���%�|C��$���]����^=xD���=m��ABd�8Ɔ�M"���\Z�&{�ˣs)^�]�Q7��wn�9�G������
D�0�|!�@^1�q��W�X������F+�組��Q܀�������K���?џu��c����\=<>�G� q��r\�>�Sai���9�.���'������׷��$E� �� j�A����+�[��n�>�j-��,��u;E�f<Ar}�B&r�P�!67�KY�:�Rkn�w?&�=݃�		�����"]X�?$�pM.��φYz�\� ��瓀g�%|�Ƈ=R���e�h\@D.L�+,sY�NH�����W�ӝ��ތ����T�O)3*[�qc|��Z��CSV�x�X#>�+�I �z��^�R|�0�ᗘS�*�u�������]�2�g�Ʊ|�������=M ��]���/6pj�Jk��[0p�j��jlN�$c �J��4X�C*�q	C¶���0|��#����K�ǌ��1���vl��頯��dC���u-Ď�M��4=�%�� z���ԿW���<g�� =:(�\�>�}��םc���չ��hO���o��@�Rp�Qwԗ�/��[1r�ɓi���x2��9���?�����%��ճ�T�[u� �MS�@�f۴�{��/)�)k%�ӊ
��7��(g���J�gר�/�W��D��P�S��)=�=�_�?�ۊ����E~@9*���_f��$�{���'UHAGAǋ_��)7�.V�bH���#(SD_'�G�g�J��ѓ;t�z
BL�m2��!�A!�"�����uXo}+K��D�4��x���`�׆�5�g�.x(�lэ_�r0��X�늪�(�B��H���o�V�*at��y�qQVr�}�`��o��g��_�8������+�
F�I+@t�5&��`�q��j?����Hj�~��XY�[�*D�M�`��l����Ό����ں��n��4�W�}n��b�n�;
��� 1�B�r�w�S�����R����"^�o�ְ&Ky(C(�O5��s�'넖��-�0�<�:bR�{��e�j���u��ҷ:�>�%���p�Xچ�S���s��H_G������8}N�= S�� ��gJj_9�sI��!C��NĠ̿��L���z��!w�-�Q���qT4J�+�H�4*� �:Ձ�� 9J��v���Q��Y��� u5�T0z_�8�!�
h,h�����Q~쾶�S�κ��I�!_�N�oTCix�\N��.��Ήp`�<��5sfC�w�S�D�u0�T���i q_4�D^�b0�9K��Sfy��f���f���ɇHG�b4f�W�x��8N��`�+�{�OW���kب(�J1����6���$�\{b��<����0���Qn12��� G�_�vFe��Ҫ��f����6���w�躀7�|s�՘�s���FV$�jLԾAX�5u�~��I�ɱ����݌,���~������B��)��E5���Y�-��3��<0��ӻ��wt�i��ѤXVW���G�/'	��m�R�n:h���z|;���v�t~��ћ�$'��ɏ4�e��5I�Ro���Fw�Y��}^�t~�H)zӝ�F��f4�X8�W��T��E�$vغ�4���9L�,��)�*�h��ŀ��K�G����[&����)��ʹYY�=���s.�0e2��9�p�^�j����%)�҅�[���U��A���?V����<u���	ώ�x�:��V����"��hNI�͊���w����~���6���D X�7|�(�3Ҡ�sS��=3R���{���&�>Aj`�ׯo�b��8��`�T�+�*���"%���?$���>�r_TUx���j��yь+0#z�K���cԊ�)���Rs�K��y���N�)7S�!�B��:�V����	2q�e�¬��| U�`�s���b��5��y�c#���l�>U�EK��H��|� �*�W|�׭��)���VRD	���rK����sx;(�f\�&�
��k��
A�̽@�����E ��w5��8���7�����δ޾PE��3V��������b���K��y�a���p�Ѥ�Fϣ�A#�ѺNk��4
U;��Z���!�O��,�p�D�� �_oOD�����ܽ�F,J���l��^$}��7FîuΥ[����vE+�����k�m�T����u攋��G!- �9���(x��V��ƹ��j1k����jO@�+66���+_��y�>�����C)U�9�]=�,~����P���$�������!m�lք��Z����#f�Y�ނ;�`�ȆҜ8�	�ǯ�22l>7�U~���9%׳#�;�Z�mj5�2c�NX^"��ݟ6;�r���c�h�ۭ]9�4���<&�V����.#I��mk�g��Ӷ���!����0F��);�x��΍�h�8�I_�X��"��Db�B�%����▂E5�!Ľ��B�q.X�+���N��}���/������٭,�b�F����'��Ez��\��{u s� �Mo���#�6,pJ�3
*b�d�����$��ܠ�I�`���''ݐ֥�k�D�1/�'������U�+�u��Ԝ���w+��y�}�wf�)-�&�6g���!���@����i�c����=4�vr`�ē��cJ9s1�L��)$د�Z��BC�c��q�r��?���>�L�t���q�N�� �7�����Vb\岮��r)�!��eK�I�<����_�?g��G�~�� $kd��y�,�|�AS��� z�C��`D2 �ԇ��="T��Q�jŊD�Z?=jwur~ ��^i�mu�z�-�PA���نe���<��+O�"��wb�� ���<���7���$&*�oA�������s{S�<���;������e��Y�[�W�4�%�dZK?X�' ���xmyT�:��xo\$4C���>S�U�;=�vz��<5�*lah%S��&e���l��Ƌ�jaH��V[2�j?�8���{nPhO�}��2�^��2"c�G";U��6���ܷ�;��Zh֫/���n�r��
�:�k.�_ զ���X�\��?o�."�ɵ�S�y��{��I��#�7��F�n�u���]A
�����e_�z`r�d.���� �{�����t�M� ��ZW�9�&�&k�sN
֖dA���=����c�,�9]��M�^���|��\P�9����F(	-٢��/V�u�>�t���T�E�S�?�ד�@L��]|��3R�[>�ʂ�W|�q�,0H�Ȍ_0�}�W3	Ƣ��p5p�\����ڸ�3%�~���1m������5�9�g�IiZsW��QΈ1�ό?Z�p��#E�x?�(c)ӊSj-P 2z�=��GAϳIԼo�ö�4���t�(��r0����6ӯU[��.�!�'D&��]'�+�ë��pmg�a-P]��rN܀�I���� jSQ5�9ww�8��>�On��x�3�N�@�C��Iv���K,���V�Tp�8tP�g�h�ꑐ>�K8M��G��R�#C{�4}Œ	�V��b�DdXG	d�7	� �ι���r`��9'֏O���d˜��-�Qn���ep��oW�(͞Gc��"�$ =>����J�	}�F>E��g8&�s��T�r�/&r��a�s�.��V
`�{ng��:�Ð�g�>��>tw����w[�(y[�tZ��הZ^�[ەW7C�+���3�2w})n���d����^�<폛U��%��x\��IH���~G��j��RQ0<$w��.�2�d�ř��� 4*ل�p[��rXW"ۺH&Ja張�0�l�~#���yB���f��x�Q�3�l?�J��ȩP/f����^��)��F�B�#�a���q3�v,�SV�{H"y�>w�Ewa)�yW���q�B��hSt3�&A�[96*v�=h=$�a����+y�X?���:8����7Y�R�	�LS�~$�8�= �	�/��~/Z�e��j�C�]���<FP��_������;ՓJҼ����'�ܯ 5T�`�e�K�z ����^���6��M���x�NA� D�]���Xd��TtC�F9�t��ݯ"��h����w���o-��`�Ls63��<a7+��ԳUV�� Vt���Ϥ��ܳ��v��������Vh����oa�����(��RK(5-�	{ۄEr�I��Ԩ�x����z|�zŴ��6��H���]���Aby0����bX�J�p[Z	��"���A��{�r���7�T�'f���i$'nܲ��U����{� n�� u�h�j-����zߎ�&8��X)��=�+`h\��-���@13��=�S�>�5�G�m2��X����.�}�����y[;�{"
��{F�6�Ѕ�B<9'���./ �*���v�k#�{���X�R�B���u����x� ,N͎gK�j��WNr)����2��@�mL�5��B�u�_d�ɕi�����#K;4�r����OS���ð��7Q�O����D���n��\��zp�s�dEwx'�����Df�Դ����:4���8��4�x��6��3?��g�ɟ��Y���a*��T�S+`�h���H/�������z_�.���6�6�2��[n;�w��$��S)Z+%�2J��ON��p��a'm�� �i��y=\�����|����-�ɕ�mZ&�A���#�����J�K�AÆ���1_sA �D]�q��fYS�b��DA��@��IyXS��`ޫ�f�w�	#	�@ /�
�m���3�6��FptM9�;mrlRJ�}����04*�%
��3�4T�	�c!�GG�'J$K0҈@1:�����*��oCՍ1��u�"+��1~I�~x�}[/�/�z��<��O#饕��n10t�{-��(ε���	ǡ�I��P�����t�[p�
#[�u���񈏙gXAj��@DnE����3@6��>�u��
�X����IG]�ހ���u�lyu(.���JQ�k'�{b����i��d��i@"�p=��_:u L��Ƴ��������}��OVU�����h������0�A�;��ۊ�������������c �Q){{�u�G�?���DߗE<��Ü�T��+/J��fq����nKX\I����C]��Xe��	��Z�����r}���j�y[�X���Ʉ7}�Le�����y�\m�.�ٵ9����@��������rv�����Ui��>�f/(���7i$|��!J4y�`�j�nY�c�h��<�Dw1k\�� ��4�b0��C�?�V�s���v��I�L}�IXx�r�9,�/
f��qF����6��E�	VH����A�?׻���d���K�ɶ6�j0�J���js�#���2Z�b�BZ�����PbjL����e��\A�w铬	�U~��0f	�
˃�ײTi@ ���¾"�h�r�s�u(&�q�`+�3d�6�E#۱|����$�b(���C<@�8hh���y���]5����C�&(��ܾf���[���-Ml�
(�j�cC���<g�����WRr鿪�+M}'�uP�2h��B݂*��G�a��o(z�7hj�r��ݠR�{	�N^�r��x����)�z�b��t{Zxt����}��U��������ot��@�]A����Q�=z�?}G��`$0�$,�����\_�Q�&��n��M����6���ζ7������&�����`����/��*P[9��W|,Ψ+�{��*`s���"�v֛��omȗ˝��F����T�zwh\3�qK,,�r��r���ȳJ�t�6����ĝ9A�?��z8�g�ĭ/ܿ��aqʠd�Ό���LO���;�	i�����`��,.֟#YM����{�9W�Ñi\3j>{ �x�����������$	+�o�NBݔ��9uY�(U��N�!e����a����x
J=`�r�؆��/�S�~�����mJ�fyD�7��]lJ�diLCdVAcN�����7;�Dd�v�ԃ��	N�tBʘrL�}p���<:��g��FpE]�q+�-�z%���4��<_��Z*ٹ�r$# �Z����g׃߰"�Z���tʯ��0]�t�#��!�!+�^H>2oNo3�������긘_�B"Q-K"��ct�
(A�.��*��,\s�\�{�k�
3g5���h�{2{'J��$���Ә��/�g��<>3�C���j�&���Y�j%V}V��cJ�~�B���J�N��u�h��6NQ�#�}�I25���#�~U��6�mδ1_�����B��0X�{�pⅮu�����(%W��o�^�L��Ke�|A\�>�̋X�2?����܈R��׈?���'�Z�X��t�+�1��i9/~��t.�ޙ*Ƨd�j��=Vs�D+�̦�'�W�*�<&I�
ŵ��ڬH������d,�뗟�w��6�z=X�sI�7���;��m~�Ή�ε���d%+q��%>��w�B�)���.E`��*:�ģ��Z��80_}�,�(�-�y|[Y�4����C�v2:�:��%���%x6�!���`�أ�."F����H�L�M�-'��gWt$���͝iI]F�'b�i��>@9xuPk�OQ�њ_�BA�{�{�O���	MN�p��%��ﺥ�ޅ�?uX������eH�� �}vМ�/1Ն�*m)=��e���_(����I)�pӯ�1B�Q�H�4w|�]nZ�Nx5�w-��(����Y�ϓ��4��޾

ޫ2������Dd�M�7\��o"� �������r�G>n`��ד�JT�.o�l�jR!��-�fY��_J���*���L���8)����Rm�K�TYͅd�H��>|�j���
�(tU��"�w\g G�]m����K��h��e5n/�s�b-�,k�S�N�Gk�er� ޱ�.IktA�[��4*!}C\�s� Dd�65/g�q����F�Փ@��.�>j��̻}y�rzU�;��G�J;Q;4�α��TT��E���g�|��*����^ �)�|$�ˤ\�d5�ynS<��@�߰Y�Mo�7��š��ϲ<���r�*��n�b�>v��!>�	؆�C�2Z�c���l�`����<��_�.z0h/��2.W���Z)
�"�rS�ŦD�^���%��+1œG��:WU'`jNǞ��bw��HhďЫ-5�}�������$����e`{1X�'6l�?6Dw��f��DTsi�D�T�r���]{�ϭ_��+Cg�W��4IC$CQt�������}Ճcf��zV+M+|i�~e�3~1�PzO��v���ң�FR��5C{-�� y�Zނ� $2��8���gd�H�8N,��b�XmCq�j�q�y��[�BGEiaL��F�cT�Vf�%`㽥YOR��\�oo׿��lk����w�X�Z6������}�(D
�:�N���L8�!,�Z���$5�h�)��B��R⊃
r�t͘QS��A4�ɭ�[+ż�.�����r�a���F�MS�y����h���A�H���ӂ#g�]ny~#�,5jV���9��K���D����)ɥ��q���Ԝ�IN�"� �x"�"��"�J4����kTD�~D�VSZ�;��6".[���VZ�ѿ���	���H����:J
����b�
����;��'��+�Q��Z��J���		�J����GU��L�uq�Ί.A��:*�q��i�wu���~���Vj�jlL���@Ͷ)%�_�h�乡��ݯ�^	�%��?J���򘖔ux-����%po���;�5�>�<͸�9M��/���4�Y�O�w���m)w���.!G���]�)��4Yb����`��b+��6�!,�g+�b�EL7�p&Dxr��RAM]����#,��2\9Ӧ��8�����p׈|i��"c��(��&{:nx��G������h~�l�ZYXx���'�ñ�'3|��@�:�Xl|���v�۲�YԨA�mq��Ws�
X
!_y=��
��c�mh��CaP��D(�t6z�&T���9D� 5�m��j�~^0��~@݆Ͳ�� ��D�G�FN���J�����e#��-K�!<��:]-����-��#� d�h#���1�JG�ixk��e�E�Zh�#Aê?��~�0�[�mnc�@��l�����4�;h�R�:H�֌R��� �k�t��[�ɭ�{����TلZ��3?��\b��'7~���/�DfY�,ng�x�����܂* �+�s���I���46D�ѓy�"3��NY�������qt�(�{g�zu?�/�f��ʍ��u�F������]�HQB'[������~��W��v��1Z�@a�_�ڙ��c����(����s�W�FE�5iՑ�ҫa�S�/S���	��ؓ-ZR�� ��Q.���,I��Z(�7���o���d�Ө�ʒsm��wsg�'��{I�L��e�)`���}}���@�Z2�(�$/�΢	�����>�_��f/�N��.}LA�.K�N�J�Qv_�]�@��$�b��c���(����0�A��+I�m6�[��)LE|V����L��Gz��:���֩��G�b}jq�m(T��TH��ͰE)�	��1��|[��S��!VT�C�Nk��3p}�>s�^�q1��D"��ȕ}�H3,2�Մ!�i��Ff�)�nqƀk\V`B5��.��~#���>�B�i�"��F��S��A���MdX���j�n��r[����k��[�I��^x4n���Z	�g�mOu`J�R�Jޜ���Nic/`P�v�X�C����J�<
<l����f|_��5�(�(�^����C턖��6;L\��vޞ�A(�$u,͍���8
Pӧ��|���y.�e ��Ś2#�H�[���~p�l8���`�U�rQ&%�bk|ˇ�r٩�z��䵉�1���!ץ�ē{*酾G��Ї~�_9?'B����&0�0�"��"��e�0�Hfc����ƄEE������FP�xG�y`J���ф?6w
�r�I6A��
@�tE�m��>�B� <\�7B�3�o��|Z�����T���d0�\��Y��ۚ��<|��z�0�[GF?�#S�H�@�6�!q�j5�-����V�?�N����|�<�r������Dh`wR��)����o07�QZ,���-�A���j��f�������~d$�|^=�]G��:Ө�3{u&fHe~ܶ���>�������j�P6��5"�:Z�4���
��2�K_����d_����t� ��	����Q�?䮊:�ѐ����S'Lٽ� .m������Dm�L�&1��=��q�N��O�.�ig����H�E��$lCy �L�W�t��A�Q�ņ�q U���1Tv��3�U⚋"Ȱ���eհ@8j����v,�ct.Xħ��b�B��^��TZ�`0q5�K%�ȏ��JmQ}bJ�o;����<��PkYX\���R.��ɱ�D�`�|̳"��]|{章�˧��3)n�.�NF:-9�� ������`�ʌt ^XH���W_ھ�K������ߒT�%R߈B�Ķ�:�WL�=�28tr�Ì��(��|�b�ˀ����EܩaV��h ?n^5�B=��V��(,|p�D��־���g���l#+���ӂ�˫%���M�=�5찄���v�q����+�1$3��;7cZ=[u�B��7��&9j=w��Pʟ~�k�,J	ZA��a��ۍD>��s��F��������m˗>�Y�X�����eF�q=na���u9h�p�s�*Z��X� ;O���j���~΅�|������K��6rXQ�є��.�t#���粪�K!��(/|4����d|���M����<�k��.�]�ȯ�M����	&TxR2�D@�Yȑ'@)~��4�`+<g�#��\�tKK��cqK�*�콟Nʕ���${��a({I��K��7�͊�!�'Oh�Ъ��x��Q���J��O�W.��7@g��9g�^�ٲ:��q�O��K���r��?(G��W��Y��c4�:�w��2x��\�j�:�a��O���g�,��F@_P24)H$�`��� 7���w��@�	�(�L�3]�g��}�KC�0��#F5����h��5�(Ama#��� �蟗�:�L|]�!�`2!���~c�M���D��VM��~�b��qr]3`o�m�ǕF�5b+�C��?��ڈ��l��� }��o;�ЋjߙƨJ�,H�;hCY�x˽ԑ�H�n
Nc�a��ĩ.aЩ&+||�$ Q�����A��Q&�g'8�>�Z��xb�N��3�yߝksw(��[���m���!E���[���8M�X�wL�GO�s��_�3u�q"�W�b,@Ouc����z h{T��؏��-����O�V`���/#Z��"�l�1kB~t�͜���9#r�N<�mΫ���q��V�3�)�
A]�����RS]BG&/d���OY�,���9�߸C�
bO&DX8�ʱ���Z�*Z�P���� D�����c��?�����Q�H�@g�u���p��l�h�uN����A�B�|P@��n�|m�菳'��؅B8P���e��ڋO4޷���[��_�%s�P�S�
C�G~�Z�%_��@��J��`"�&!�#���_��^�mue��`qT����F�O,� �(�1�!���0����#�_���@�C�b Qc5���"FE�5Ecq�X��UtIzt�s�������oٝd"���5�RH�������Dڛ-V� ǁ���-#�xT6[�	V(�;ɷ��kA��̭��g���ᩯ���\��ҥ��P^�V��W��\1r���[Fj�j�1B@u�e�}�7NSz���"R@y��{��^�P�?ܾho#�qF�hI��{�|�+����o��(�]�,�ⲵ}�JP�Y�uQ�	�R�M�:jvZ�&�@Vna��	 *���S��?�K��=ʝxϸ:�f耱��g��fx]�0�k|�N}��k��P"��·!w�m
�l5����A��Y첧OY��YGVu��\�Po���u�4P��j-�o�d�&�J�� �!�rᓩ8o��T�X5��/�A2~J�!|>k����6Ԗ�ï��ނ���x�@+@q?�/WZ��zJZ3'�ŵ����_�_�]��S%G�6��#ο<��Br$�4\a?鸼>w
B'���a�д9�"p���r�+THv	yZWHG�T)i��e>���>�R��۷�?����"z�����Ơ��1�վ��{��d��^֎��(�G�պ��uOx��k#;�ŵ|��.���Re<ޱ6���h��DW1��P����w��е֏�B�f��eb�7���;�A$�|.���S���V�!8�2Ɵ٘!�A���A�	�]_U;_��:}�i6L�W����Q�Y��� �g )�N����1ڸC���F�tA!P9�<=�����eDV�~�+���Vc���b��:�u�&�+셮��ʡH&���4�g�+��#r��Eꫡ�&��2�FAg��Q���m�/��=s��8j��7����!�+��B'!��]�A���4��m^bv����Q�]Ʌ�������"�pb��j�����Xa��Y���Q���WTj�X�Q�^f+n��[�ImU~�ؒ�f�l������=��Gz��9�}�fC��p	h���@��镛��V�x/�qg��L�gB�"���\M�� �E-Rh!v���S����L�cD����R�B��LpoX��r�X�C��i[��rcx�wweݸ�z����<@�Ȟ�|-��8߁� m��,�R�ʤ ��f��t�.'ݠ����|�a&3����h����2��6��d 4�R�ǖշ�,'�7�YzU�}',�-~�&�7#Q@C��a)yH)+Q���!��몂R!R&�� �"��b�"Ѐ��}�?�1rVd���/���G�)�]�D��uk~�?��АrrEW��7���P�A���1pV�菈���+����Rr���~��]��X����d��̼����W�z�M����o1�9?H,�L�ɠ T v%8�[kN�����_!��E͕�#ȴ6𑯝�˜�h���nD���;��ǃ��� �7^��j���%V�j38��=Z�`_X���tD0f���v1�{dm�6�
4���L�uP��:Um���Ym,R~m=
�X�����G���'����0���֖�l��x&ΚB�!�0�"�O��\��S�����jevyM�i�M��*|t�A�{SU}�����KfI9�B�Q<]����hDzu�F�tf��φ6�{�F^��7�����떼�̳p<D�]�w�ȷ���J1�`�vWU��Z{-��
}{��Y	�R:۰f��K,|R��WXW�5y�oɪpu�s�>7�sUś�O>���U�[{�ֶ�x�ĶpJ=�a8�Vͳ]n'��b{�3���7X��]�Yl���6�߭�#�x�����30��Q�mZ�a�+�>L!����y,ګ��P�|��F��N5�r��1g=��ن~����A����o+6��^l��Dm���)�ʜ�WR��/ =g[S��7i1 j\0Cܥd�i�E05�ͣ�Hz�/K������k�����O2��c�yD�*sHv�6^֧�iz�
g$v�ބ���3 A�5h��g'?�F�\�6-��y����������iC�N���z8���Y�
�/����h��ӆ����g����Ѿ����7��?=�
��/$Pn}�R������X*��M�q�J��܀���0��A2�B��S�i_e2S��J�9�S�˞z���!٣;sQ������>��`5s5Ri-M��&��e\�˜����g�֯oޱ�4���xq�w���HP�g	Z��K��2�=U}�v������MM����맸;��ȸI���1N
���j�-ឥ"���ݢ���<4n �.վ�g꺅�m�鿯�i�r|�(�些zX;�,%v�"���`�:��V�0��w^�Nt�3#�����w�^� ǛU�1���tQ����ˏ0h��D���`�g ?��_��DxC�P�8}"�C%USXDd�q�,�r"ss�`���LK����s4����By]�=b9 Z�!3/Z�CO�ߛf	輴?k`���C͎t����&����Ƭ��'. ��
���S�������U��\i8�?]r����#��'�^�X� �p�����G�L����!�M�9N�H���TztĽ��� �/[u�yS�E�(cy�V�o�Q�,&�?;��ߘ�xH3��}n~eR��z<1٭�,{���9��\�P�r<�0�vb��)��Z����|�+H��r�߀O���=C���F�5n:?ؤ*����N�/�]�U&F���J�(c�P+3˴F�V
/�y��t +]�����s���V�_ ]W@m
)M��?�&���s��!ATD�@N�k�P��7 �R=�R��'�Ó�/	0_�m��9�����"r�hX E�S��AV>��p��4�d��%���$���o���0I��2sY�y4a��:���P���gl��4��&��*w�wK�.Q�p������A�3}�6:�%G�Z�F񦷘a�Sp�מdDF�U�cE`�#�)��`"��.RD�l{���;z7�n;]���K�J��,��*A ����7LwJ�A�4<+>�c���H�v���H�9 ���H-M��J=��d���������@}�þ�w���'������3���d ����	�ô�=Gj�gk���6Y=^�\��6�	&���m��Ye��U�{�Z�B��p��^��^.s؃�Z'I�*���?ZyY[��;���~���E�a��{M�đ[�*�,����̷��rs��)ag��mʨ�޹v�ㄶ�m��� oڳ���[��V�M8f���.D;�hN�މꬶ������r�*��K��ڶ�c�D�xۺ�?*�5dS�	�c\�n���W����LC�����K���:T��x���P:��e(X�|te|�i}l��������_�2�b�2��tv\ ���2�6-n�y��liJ�fv&T(��9%X�,���9�K$�>�7H���b��OB�Gg
j6�U�Qi:Z������?G�
x���i2��r�
P�W��M���(EbZ��L~�����8SW.�SAS�Ϻ�j�m��xN��I
��5��Y�5*�`��xά��(����Ą@�©��ꢑ&7�j���_sv�mf�iz_R�;f�����N�9V����`m�4��-�;i��{�=�q���~4d��V��*��C�CW�C�Dz@LħpC{�/44𝝂��i������x��v~�5��蓷8���㈕�ϋ�Mfo��>���_m�;�˜��c~��p���T��R����M�NA���s��Z��|��H�s�_��Ybb���,�ld����9�`�ƒW*�/�񴰽���yn�X�y�K͋j�lt��bL+C���p��*-���T;�g1 d��A� @�H�&6m&(���k]L��Y!&R:w��T�;�p�Z��5^����-�
��Y���Mֵ�q�B*�W9��G�����oΪ�������L���D�=�H_�M���'7��l�x���$Z�r��o��!�6>}>ɐ*�tz�y���"n����S��<��W���e#a=Hk[��3|S���A�^��&����ZJ�[%��'���y�}���=���@?�H�^Pa��Q4Qz 97�Fmf���ıj�/)_�|�ju�3ͲS�i�d��96�f��+*�#8�"�&�m��Δ���sƭ���+x���f�4� &�h�u���kc�u������l!�d�X|X/�\���=���P�����L2̎�T-�\!��U]���)�ر�x߿K�"3��ъm���sH.]�%�*�u	�����,0��fҹ�!b��� v�5ε'�	�'[ﾚ�[��+��2e�C>�1�K��4ܯcp�Q����#��ӭ�k0x���\����G6�[�$�p�%2B2�-��ueq#lYÇ�¹���J�sN�F�g_�������� MY[*-?�Jw?������}���eј�z+��fr�(���x9�#�kb��NG��e��\g�ujV��ʓ���4�𯮱F�`4>���5�{<��W����*���v�Mm@�/?/����~��uςP#c����p4�jB6�-����%*���oo�\�mq
!�!ۦ�ڿ׌��d~J1$��|i��w��lj���R��V���o�mN��C�ot�ğ�)��/z)`�ǌ�T+_O�N����h�5�ҮEJ-���|
���&?'?-��u3�D���	�]�-��Iq9}����C��ќG]!�p��ޞo�줔��U
b�}�-�X�d} =�a���k'2��˚�RS�����v~�R�R��-Y<�A�7�-Q�6SϚW�3=�^�PO@�+��1g�O���_�[�b4@s���.�7{X]Gr��u�=���f���Ǽ�� YJ�Ɋ6G��x\
��^��1��i����')�n���f�XFv��W05-��DP�wd�4�2�8�~L�oT�OҘ���h����j���� �*�>�@g.�0E��ҾI8��+��Dl�T�У��'+Գ�$>�<��I�c�ـD��l��TՊ(��f�_C��#4�qpm|�P��$��W�|b6N�WJ�ƙ��xKוu kB0��1�d�(�V�:�7̘E.�Y����sb� ���ɣk��#*d��@�?˲�/�����F���0�2�|�Ág�1����{=����D�g\CL�v�]g�7�c&�x�g� �$��������_j^�*��U"4��X ;���Q��SRG�C�$��\)���?���I'�~�V�J���8�E�b*E������.nF��1,ż�2��ų�a?�|"=�-���5l3<+��W���Π�-��6g���9���gNPޛgsd�%g���c��Ǉ�[���U<�*˲:�����H��K(Y����h�5/��ƌǑ�6�G(�QlV�#ʄ�x�=0V׾L=E���>��y�j)�p���9�d��F��X���;!C�<K��{�;c?��u��kFק��\aR!1�mrNeA���in�G	!2�UGI�Q;�I����쬯��?~�����GA���,�ƌ�T��a�r�{Ѻ��cÇ! ^�=[wA�x��bl�5��p�Ha�"\k�T�;g�2	��,Z����yK<���3��_*إRۘ��mj�_z�������p	��.ddw�Q���1�L���Xr�6�:�üm�K�b��bW˙2/6%���[�~����u��R$ݡ�񿵉�>J������x�\�����SV�(��?���Υğ��Dlc�������h�]����$v������C��F����k�*٫�Xv���Ux�l{�����pA:.��ѹ�L�7�������ts(&Kk@M��'I�����dJM��/}����H����y�Z���uO�J�>֗ݪY���L3.�5D�ɖ�-��-7�l32���|f�QV�#�/L6��eD@��\	��=~�hdoE�?Y�.��p3��o�_I�)�}�a|�}�307f+����\`��3C?�|2�^���}��^l(>Q�'&H�������J���g�.N��³��*LHd`$-�4�J��~�y9�k�%��(�=1��ݩ�ܨ�	�e5������^��[$�9��)��#��,v
b�d��g$�<庻9Z�U�`&�Jq����p5�T�!�蓒p�܊M�y��n�I�GN�JZt	�Oa�%%�\��4I
�v��-7-5:t�S��ݱ¸��j�!��a����u�
�xx�Lq0�m5���gz����cQ@���0�'���~(���祘����t�r�<��,m�|�b1�.����$#k�oP���k3�=-mٺ�"�3W��|�����<8ʃxU�x�C�3��.c)�I���78n�����_I��R6�_j�RЪE|!���Z�i��r|4
����=o���0���-!�1G���-�
����`l�""T0��ua��^t�ll ��{z4=!�x]M�	Q�ҋ�%���됚K{)�k����=1�K���6%��y�.���$���d�ьPC�Օ�[@�����,�?`���"�(r~�����4}�-�A������[#͉i�A�����!۟�U�0�!x���#�àЖ7�<~B8���L>эZ� B��&2LcL�9zQ�t�B��>%#hA1q�e+����a$�=�x%�\�A�k8��l>:�x7��B ��?�|�~���G�r>5�$l��nWf���IBl�B�
�Y�ʽgf���.�0�S�y�[�>j�R��@m��~@�'�B%��h�9����"��_Qhљ��G~�!iNIP�7@<N��K8Z<~+����eE��"�yky�o�4�m�Q��21�����Iv up�����°i�E��(��΃w�\��͓<<_�H�<v#�kU�dE+X��zVN��|ŕ����(�*R��B�\�Ω�a +l�.
^�L�AY��?�`�o��3�^60��(�(yԉ���r�q�`�y����Nt�As
�g4fM�}>\����1� }�u^G�R��LoUH�4��#�`2�[�;�v�cƯ��������af�7y��?�N�&����Q�ZVo���缓6��4����Թ�<��Ҿ�����[A������ʮr�'MXn�b�����k�� ��[?}*j���<��Y�������i�tg��n�d1C�yX�bc�2��G�{�h=���Q���;��v�8���EH�[���[�'crY��!MSi�"�0�*�z�crMK�.�����_mN+.�"8�a�g ��� qE��9���p^k��E��,K����baf�ʐ��tz���fY���B�ԬaZ���«��ڑ�����(SmR�M���z�0`?���Ud���X?�*Ċ���m!��v4k>��=��FZ�$:Rv`}�u�<�\?�[\$�ʶ����@�`7�j���n����<���o��3�����`�]N������R��0���ǃ]��&��Ù�!���M�:�tDb[�&�� B���/���u���h��e8变~���� j]�y�/*z�/N��Bgm����8��)f�͟��@�@�Z�0%�tέ{!��V4��x?Y�%��_>�.����ң
���1�}c'��,'�a���4Q�S\�u%��wܿC�I�+�:�$�[����v�'i�B֧��7o"��_*ꟕ79\r������V����<��xQ�Ip:����k8���~�Dۻ�_֪p �P�q
ɀ��������o���?+�J�����n��̺�5� ���^�	�ժ����('�2 �4g(���p
+�N�?�Ӛ3�R[P��D�[�S�@<�2�G;F�-��3��>1��\�w�GQ�(_D�͡���Ȯ�g��3ʈ�, Y7n�ai�o
�}6��*��e�yʁG�oo/���3A45Yi#`)�&��S�i�����Dѷ�������C����������w)O�2lȣ�����_�s�K�L�|�&16n��C�ӹ)$櫥�$��X��[z#������`�&()�|�@�q|خ$�\D�{m��i�����៫?Ӹ���;��[LwS�i[�-�B��Ս�61���Bܑ�4���ź;B�55����az�=�:��eǆ!%иN�]ވ�P�=�ҸzF�����Ck�:^�p;�w��UW�V��ީ�ox�����Y��:`w���8@\�u���<��E�F��\NiM���p"w!X"��m\�
^�-��^`&�A+IB���I{��*VZoU��'��O�MPC��fFO'�_")g�\<Ŕ���a �M-�Dp�z�Nd�K��� ss�4u��5����n6��
c�*�IkF��C�ȴ�!��jS�
#}���P��?V ��04ݺ�g׎^n����׉KJn�qB:�v��(��7�7"!~�uŘų�>�]03g�}�g�#�Ӛ�2��Ӱϓ��:�;T�g���p�ǖO�m&�b�Q�7���%,w����`��v�0�r5��Ƞk�\y�L�rC�B�D ��&���qp�~F�p@T�n�����%�/�Æ�x��E����Xb|hP�5��8� �F.c�E�I�`��C7&����y���\t)4�`�$����J���m$\/�]�+O�x"���|���嗰O���\qJ��̾A��4�d,���@pU^�a���B��@p�W�I,k����ť.�+�oZb3SlV!i�g��������la����6��sd�s壻����W��䰛ޑJI,�qBEь?)���a� �Wb7�yڟ��j�BC*��
�Bfi�=P� �Y
��ft�V�X5�r���0(�ţ=�Ⱦxζ�I	T���ǌ� �����O�.��y�_���w���^��მ2f��@]��Ⱦ��C��b���3D&��"n[��d��R b�����_T�~�!�6��װ�����b��@�Y��h����pɪ�y�z%7�d_?M��娏qny��r%Xk��}���
�5����m^���lN��ꒁa���`���|�j�UlX��8��b�`A�B }�!ܮ�ؼ�;�Ima�(U������aj�܏��JӮ�#eQ���;�} ��&�1i���ld�Z7��b�P�<IRX���u~��?�����m�Cz'���ת�I���G��1\�����7�?����Z*�xyF�H�u�o�j4��0E���쁷H�N���:���汵0+�HO'�L�6�ZxѱI@1�h�$g�լ]qW���n֡��9��>�z]E�Ώ�&���3w;�Sui��l���V��!�)o��oÌ���A�U���)S���6���71��q�)G�-Q�4��I��q�-��dt�ch�#�Ɓ$!=��ʣ�䚈3��s�Y��|P�zRtBŠ��G`�z�,
��9��xd
̢��c�y8�uq�����|H��\<J�I�^�����D~	x/��q�VİK�B�a��s�7�܊�G �7C�\�$��jے�-�>�Ds߾9j6��V���l�F���b�� ���K���ꐻX
ʥp?`��p�{m6T�b.ɓAF��rw$�s��%�`Y�Ƈ�6j#K(C���}b�G=U9��z5T�Xʲ��} �Ax�ĸ#��G��X��W�b�4��V�	��i<�b��j�v�>�@�	��Ts���g���z&���8����!Sg8uS�2��>2F�V=e�6�!c����B���2l�*������Μ�$ �a��C�T_G�5�,gR\(���h�������N��H���ư_߹{:�En|�!�=CG����Uh����Nk��͐�TP�H����)U����DHb���:����
k����5�N�$�Y�|���M��<'��'�}�챊$��99#f��[r~ć�����J��Z�q�Xѷ���'���K���F��72+B��w��I]�ϊ�����|���=��Z���Q�D�U2�Ͳ<��4,_�6��`f�D�!��l}io��e0{���'0Xm�h	t������e	oZ��̺&0ʞ�86�4wZR�U��)윸�րb�n���Q�Y����HbX�JySo7��s�`:����|���$�\>}���c�|G"�	����P<C����ϜQ\h���c�E�i�
bt���Ǯq�Y�G��,��,�'�=7��>�e孼fDVlT{�
�R뉉�����GӪ��
z�ZQ*����/����#- +;ٺn�ż�\<z��#L%d6#��fj�+�A�dٷ�Q wI�ŗkw�Ʋz'�iM���F���E���?� ����C&d��>͞,�0��Т��8��f�a-K��S��RX��u�NQ�?^M�h��k�2e�e��q�ψR�Q�n���g_F:�8�����n+k��焔��<,'��ΚB'�"�z�\WJ��"ZuMP4� IhI��	�)9i�O?�?ꈨ
���D!T#':�o�^���'BKF���t�8���=��p0��>x��>��t�|�;�1`�kc�G�3Ӳ��A���Lz���i��:�s������߆}���2�IeC��<�� U����éD��l���P��~�#V3�	7��a�>@zSsx��=P�;��l�x�3Fd����	h:�j[!s���_���,Iܕ9z޲~i���lSj�;<E��RY�K����@ .��Lc�/23�Ci�逻�̇���+�>~Y�WrF�J����&Z�Jنx�)[[eG]�v�e)4W��<<#:�eQ<+�?�ս8^�x^W�$�oƫd���cz�=R{���+ܛR�Rps4<R��"eG�4�"ZG;����#���5�����/�"��[�W|��іP{d.`�K�L���<�u��5)���V�S�[�	���ٓ��qn��:��^���K ���fO]��T�vSړ�V���L��U�O܂|����բp����ҿPʷ�:��?�ԑ��aA�
~�8�(A��~��+-
V��;,���O`��� ���i'N�h�?�9="�|.����.�o�UK��:���l��\YG ��H��ۖ�5f��}��_�,�?S���sy���[��z>_�rD�(�p�~,�(��i,7 ���8&��~hD�!u��͝�7�4�o4	U��������0ѡ�X�o엾w�2��L{�'��w���&8h�ۜ�9�A�=lP��C��WT3�6�<��Ll�:�r��	��-s�K��@�ou2�2	�A3���R	�Ϟz��	Ι�[n�m���J{�/u�,�k|ĩa�������o�ǩ����w�笺��B�QIϮ���Aˊtk08�R
9$�y�ᝁ��Ćm��D2A�9y6���k�{��c�B3��)\��֎��L"3�K5ƣ
M	N����օjl����r��-=���W���v ���	�4IrQ{ϓ��%dX#CF�*6�y�þg#��α6
2M� bՙ/B���J���6N�%�
"����Lk�ŷ-C���B�,2����ؤ2������P�;+$��\�=�>d�^H�Y�/oЦ$��]����yi��L�]���=Y4��
���.�=�muPhQ6���[9ޠm9M�ļ=����/�fU�4����Ћ ٹG␿���3�s��`PA����vD�Ax���>?zA7�JH:�J��Vᮽ��'o�i��H$��jf��^���w8Z~3@R�0x�B�mŕ���6�)�]�dJ� �g��u2��(�����9�T�)�Ϋ�������x�et�e���I�ή�m\��n��X%duZ=,��V�A�t&��8�h�(7S�"�cbI9���-#��᲌s����WF2/l8��BRc��@u��&۲�V���R[��}�u($=aW������F�2�w�K*^#�n�j���l�}[9���Y[Z<j?����@c��gV�qɀ.�M�7K��c��`&�0��YT��T�i|�]-|�&�*=�() x쐗��b�l�T������ܻ�Ͳ_x�^�]�H��,t����^}�"�x���;�������0���Gښ�*H�ɦ���W�����3H*�Z��p�a�Щx6hO��<
�w͍S_�)	�s��^���[�<�h�M:679 ���� §+���ȧx�����x����������^*�t=��IԒ����F�oj����T!#
ruv��!��B�'��Jo�Â).)���	�����4��c����C2O����ÂK�iP�l��?Q!|��#��
j����%��)t�I���S��LS�a-����ve�G:��U�e5���B}u{Zn�Ԣ1���ʻ�{�3Wҹ���*j�#�.$�.�1��l�J��܋~M����ҟaMUأ5�9�G���If�`+�S��4��JC;b(�w�L7f�����k����.m���ئh��!:{��p�j=����jT5k�"�g��CSzj7����@�G�9wC従����Rs��� ���;c�B������*�E�O��Ǒ��紀�N�H�;��Y���lM	R?/�����0�cd�_.N��J]�SV�g�ʓ}����wJ���o�<��^�R���M}�|�P&p"�Q΁�����c��}���Ec�n�!�/o�����x�X4�������:ܳ�g�Srn���]\��t�h	-������i8�Y��+q�r�둈?\��м�x'��������EZ�[LTI�5x杏��te�R�y��h��%ZKldb���OKL��	��Ԫ�`Ć�
!��R��=|��*���Ɏ����7{�K�Q8��dVy�� ��nG�:�� �e������H�����PVWl�X��Z~o����ໜ(��I�W@rqR���q�W��[_iߛ��7'�L��m��C��@�f�^8�k.h_"��$v(��Ѷ���7p���_j����*���޵C'���~)���_��ka.�*)���m�w�BEBvYdD?NҀmt�E�:7���1T^�a-�X�y����,N����&I[m��s>���
�V�PI���GG��ݾ�Lз'7��c8,�#jߒ��&�C��
n�U�{C_ ��e�v�g;iZ��gȐ-�_���i�!��)A+r��b�6�����s��2QM��37��g��$���e*��e�T��;��8��B�Ҋ��ϣ!�£L4P��h��'�
����	����&A4a}a��8�`s�-�}��9t�R�a��$��@P���������- �=u4)˛�1��E�I������ �R�[_�:6�Z�v_ݯ�ay����I�%9Xt�p��D:�w�4�ƍ�L$jm��Ն��fv�w��Ҹ|�W��+Ru������>C��`g���Ջ�,�m@	��j��_�4���N�t�X��&Y����&���u�1ƛ>,>��'&�)�
-UĚKֶ��]����A�쑤�>�[6��#��:�&�b���_N0���k|�>OY���/p�l0@l�0���=\ô�rqNS�m��N��>Gu+���އ!�m�`�%���
���}�¸���Dc)d��5��ۚ[Ü����䢓��9�?��,�MS�6>G�G��"����)0�Hâ�&�mT=�Av�}�,��i!ܟ?(�(d����,�|�OI�R�5�3x�Y��ʞz�R�:F�����7x�q�-$՝�j�yx)n���������Ә[�Ģ]�H��Dn���u���u��e�m�=������ؿ��ȶ#���1<�k6��0�j�P���Yi�o�� e��c�y�/Dϩ��*�ޱ�ym������U��ܐm%������y�_�: �0����)�r=���a��#p^WK�G����l13]���~���D�3�G*y�?o���7<�"��
&��L�8�3Є='��ŽaΥ%f	��-;r��]U����d�"j�Uۍ�$�J2E���:r���9��GS���H���K�y�L����A@�a�x;4��d��܂���5:�a�װC�L9Ծ��G�&�B���K�e��7��Gk���b���!�s��0�Y��Q�ǡ�E$��3y�F}�|~z�j����_=�R�k�b�mט��3 3Oz���Wr������uׯT��� �l���H�ܕ0L�G�A*��C�8�o\-A\��PRM4�55���g�V�z�t�'=��>Eg���2
.[,���\'�����,���M�ȗ ?�)�5A��#�-��!��f�4����t�֜^��I�>��i��}����	_om�J��V��v�#���g�:"����}�6��oEb����-Wuc�Fe�I���=�8���ڊ=$t���r�l�~̴��A��A׵��'|ô����Z�rȆ���*◛��+y��*����N-jS*~H���d�U��/��6�gR�?����w�.��c7�ez�re�\�2�6��Mg|_�I�NI!z���2O@�_%�pfh�%�n�*o���U�l896xH��y�@�=�:��4�Ֆq#��1��&��Q�r�ê��j�t�.B̷A�׍&�Mq��@wW1VY�9���8��P	�����jW��핶�ѡ<C�]��` T�5��i`�+��XE5H�uC�QZ����eaYS��܆�����B����i+݃I��I�/ۅƣ=�E�>A-� =��R2�gtꗣr��a����s*4���@}�(�o�oGA����(I\���ϋ?i"����;����K�&
�[�w�P$�B�����Ҕ�PM�����]T��$R��J�Ap�3ʄZ8[+х;Q�:�p�Б�?��"���Ů�`=�C�*���n��N��(�O�ϺB.�]%Ֆ�~�y �r&2���MX��n{��!gb�*�x��Pk�z�[V	/�{G�p�#!*�?x;��G��@|�[�<N����k<׫��8�o��L֭t�y_�*�n��_��Τ�0�|��7���?K5�#Q�̥�eã�
mt�7l�V��%�)	�R�B`X�����k�j��2�ĉk�P�ێ��31aA�V�J�v�����0�D]v6�n����t�r����7v>�Edga~lv�n���.it��o���)�JPM�+YF?��C��N�ˈhp���u��� �0�ve��:s	@`��h��p�?�頔�6s4z|���KX�&%+ɰ��K�t�y���>�B��y7z�����/Q�xB�S�_�*T�F!R`��	hu�P	��i*�IL��G\2Ճ�����	�!���cnh�N�9��/xO5�68RiŞ��)�G�5:=%-��d:��8F;��F��~qC��FV������!R�8ZI�7ޕbU;�b,s!,��k0�1s��� �)Cm}KC9��OQ5��ߒ���d��������<���n�P��)�g�~����ɥ,[�]|6G��(A����*z�ߍ��!��#�)��
�}��6���r؃<����|
+����J̠)7�L�Quy�ٕ���3V�Ѩ�!�f��=f�R�O�:>u	��2l�D���jM�b�w82����g�	�s��%kV���7�����q�Jf��>M";V�Mk[/F嫢}W�-&"�Jе�5J�K�=�]���&U�/מ�yhnY6���cmy���ʂ����~.B��!s��3�%�2s#�h&Ρ����Y��"�v�`���|�e��z���� �_��`ݡU�i�2�!�&QWc�'�������&mGn���ѣ�����K������X��_�o:	�o(ܐ��wb���x Z���B�}QP*Q������u41(��*,fb�L�w�пnM��TZ�]]rĠ��U�U��G�?ֲͻ�w��,i�_�L6�ڌQa���X�l6�eRA��s4\0��mcv���Ie�� ��ҩ.ɍz���#h�v�"<1�a��2̈l�m�� ۡRmK [+�z��dz65v�+W,#�A���f0�k�qs�,�p6�e�2�4��fJM@J��_��m�V4���g���U;�F:���3f�
Zd��a]�&/��
@fι�/*�H�J=�d��_A]J>I�q3:rπ
�:�ȓ�a@k�\��pr6be�b�xuaMvh�er.��,��.m\`P��4Jαv��Z��R@v���6��pnoߩ�����.)ܫ��� ��`��KS���Te��EX�[Y��d����(�{7�[�3��.�,Nӽ�����nЗ^$���<3�t�cĪ��8*T{��Xw�����X���j�m� Uӈz�{�oq�'�hA*�ˊ�V�HŃ�>6�tV��Ĺ��u0T�t|��;JӮ��d[B�� "k�>����q��=�?�������ݵ�a�/�m���5�+w����KIy��܉�Nq�h�#v�HM������\�kӢF�v~f\�n�y�#��Pj�'��u66k/���{�1,N��}��f����N�^O����w/��?6<m�7��oR�\��tU���v��#zf~I/��S3jJ���^�b:-�_�	��j��{�B��uF���>����lw�[/"\���I=>s�>���TK��Y˂RQH��ؿo�{I�&|��R�ge"���iΌ^}���o�+T�r�Ғf��'� ��6����)��N��㋏��5mAN�ئK�i��������>��uqT�-s��ozY[캬}��	�z6-�����	�5��#7���lC��*5nx�3�qKP"��@�7�æ�?%�ĠnfVy}�Y��>(c���0d�����q7^|x4�9�"B����
i�}
�3s��O`��bⲥxv��w�ISK��l����UoNb��?Q�����+w���)IB�Y5�.E�{�$�����8�ZE�Ũ�3 ���Y@Q��Q6R��B����o���+~�kG*�;�[�I!�u�qr��ͫ=[JB/5qWA6�3��M�ϗ�1��/9Q�����$�v�?�H���?�7�򋲽�&!c��_�l��0hQ�Ԗ$e���
9T'��_���إu`�t?cig����^�Iҭ_ڊ�^}EQ�[��V�-؃]P|�d�[ׁT�sM��. �X陮�(\��#ˑ� �+��'3��4�ȯśG�J�GڬB�6�Q��F�91�N�(���bcq~0�6i�uƶM`���<��H|p0��޶ض�3�蔴�0Zަ�uW�A||���t� �A�*Z�/�r�x
3�FC|c���v�|\V���i����9To�����X�#��H&�ޞ����YW�<��Զ��Jm��ac(����^.8MF�Vz��`3,�q9��������`QH�	;%U�բ���7����y�IT(��mW�&J����BC��,��ՎAU���ҼF�#韨�˝���ϰ��Z��a�����S?{(K��GĮo³��{VS����z���v0a�k)rt��F���?&˺?t�$���n������Е����S,ެ��T�r��we�Ol��j�#ko��_П����$�X�Ә�6G�����1�q/�I=���\����Y����S���v/�r��SW�O��ɫִ��PB�>D/W�c�`��45�_L�G~�џ�v9��q�8�C�\� 9���i��N�y.�#+��� ڰ�K^�p[(�֛;����h�B��v�+�/>��9�3O������\�w�J���k��MxAW�"�.t0��ޝ	�}W}��t�7�2@&�rx�Pίi9�n�jVfw�HK��!t�	��A��#0����e��i^���%�����S�('�*�T�m����Ll�I�JZ����=�f�����K��]��Ҡb���jz�,5���MS�US��8yߜ��V� �a&HI�b�d������e�2��!!�V7��c�)�����|�}� <�W�[�]*aÔ�5�2�`���ig:�?q	×�vm���1�-�/À���N��Ԍʬ|~��zQa�w��;sa�E�Õ9�c�|�,-*�'��KO-l��>�P�3.���-�i *�(��s��'b��HvZ���U=w���R�A�s��	Ȑ�4/��(rIT-�}�P٭�7���B ƣ}>�� �VBX��wd�eOD�|$(� �]E@��	��6#��Ҳ�*��3�ڝ��C�v6��T�ܗ��1�\=��+<pY��+�h������oQ�#?ͮ��\K��*�ޘs:��L��Is������Y����*&�2\?�3�d�x�YW��d{w@u�Cs9��h��r���=��!j�ԏ_�Ve�.�=9��K"�Y�~>�I�G�E�����&��o������,y�v�;9]XWo{'dUR��L?m�1þ��f`6���%8��{=с'�z��� ϰ�>�&���J��(�gg�.R�a5P͚��b�Џ�} �H|5��AW������\�'�l��љ(�U��X�s�(�"�Sl�i�jQ+���U���G�V�_`YDY&�?%��f �w+0��q��8#w2#f�7I٣=��]���)Ju��}���^�@�C����k^�e��s2���� S�q��s7(�äᜐ��Ŵ�pa5ơ ]���a��Z� ��)���eh=�>��2.�y]�[ïp�T�l�V��)�)������X���'�%-Z�N)1�+�܈uj���.�(^���$(�oťm�y|�p9�=*!%���-���V�̶�pp��xj��C7Ua[�$^pR�1~��ld1��u\��浈-dQ*Z���"��"�r]�i�RE�y"��T7��+8S8C*����p�TC��a:�{� oq�Bj�y��/��@|f�'���ɛ�]�*k����_�~�LӉ9^�qBkɰ���o�\��w�9׈��-��-&��0���i�O��c�T������(���G�w[p����+���_Sm�T��A����]�jR�pwqO=���?/�d��`��<k��F��b��n��|�	:�8f>���j�ea���)�Q��B��.q��ɓz�!��W�'��D�|v�]bg0��ƣ�ջt0u��)�h�~�{.1φ�rǋC�W	����
Q@?�9IY�3 �;��n�)�Pֽq.��Sn,�S'��J��2g<�R��~�<��ŋ����o���F�(Ó�w���r���*;�+��Хs�|����
vW���eb�a�����0���2��\T�g�vi��0�O9�q<�I��e�����Zz���u�^X�R�l�s}�J��D<Oy�m������5�֮�����]w.q�����|�C��s�Dbȶ�����0d��K�ئ�b��8֙9zO����W_w����	�<U��Aڱ[���Fa�X�x�M���mm�)�B�����/{������{��PZEe��;bn඲=e�U�Nq��pT�k�����[T@c�4�z�r�z�ѹ&u����T�֨Pn"�]�|j�F�z�.Y<ә|d���@�]��J�k�f/RH�J~0FLEf]l�I[w�v���)�x����:T�����%��4R��1�|�����fr���>^��7R���3���]�5c:��7g���k�6�NϜ{�8�AOE�/��[��L���T�\�J�Q6��̘c�*�(��E��C$���(- Y�"���� 38Y�	��o	�%W��[�;�>t��E�AUb��f����6�AEhl<XS$��o�42Tb�tyc���^J�]�L�`}h����U��[S�L�F�5L�$��e?�XVվtC�P:����Z�P�Vl1�vكt������7�r%��������l�z�8��F��R��J\�,�ս��u����@�hH
����'C壔?}́�)h��� ����z�
��,�'O$a�QGu�^�͵���RN�1�܂���0�6�lG'�댛���YB�	23��Ik��c�@�!�β-#���c>�ǃ<ef�d{��6����n������˫X�8��n�ڬH=A�^���ޤ#�����ʹKһZ�?8C4�M�o���6*��Z��lgm�2�z;�i8��0��R�V:/���*���$d
ĠO���]��F�l%B�z�)C"�˱�3� )d��w�0H��!�Ҵ-��R�eƚ�G%� }����+^�0�5Ư���J��(�W�XA���mI���C�u���J�y���
��sz�@� ���[7�y%)���y�3 n�n�Q��h_b��g.0��`�WB�#EH�q�fa%z.��(Z��>v4�8�>�
�#]!	��Z�2�#�Px�W�]��>�9��hż�-O$�P7��=�@��Eɜ�f�A:
�͠!�r�H�u/�q�W�mGC�u���_A�H�l\D�'���������fn	�Ɨۿ�'�z���ٷ%q����X��� �;^�.�9�UɌ�� �B��,WV
�Ts��7ܦ_� ��.Rb��xx����? ly~��*6��#�������Z�;q�$�52�<;h�7h��P���]RAhQM
t�z�Z�5ƥ�^���0�mc;���O���}R��hH�`0�V�����#�%�	�S52�#U[h��7�PF��;��&a�*��?Bw�D�	HqiH�ٚv��9.�r/S�U#]z�Ri�~�c�u��D����%�������H��OD��-6�d���R�GRd�%�2W}+�l�ߓ�#@Q<r��C��oi�4�٨	��;oÊ����zޙ��������<jyOX_�i��[�p絡ߙ����_&7�*�_�
�S���*�G�^IA���9�2�N�0s3hM�%�a��%X�<7<?YQ��$�H�5���Oa����b'�<��Znd$�'�vQ:z9���ncߩ!~�(y�Ζ��,���3���~��<z�!	~@�L˫�7�]�Y3ӛ�	
uw���Z��A��d���[��L��S����o�����1�g��+��n�Nda��<���Lk�
���C��Z�D�ޡ������+��i�t�w���x����^�G�ke�3�-��D��G�y��������ޮZ��a4UnF7��>��L���TAe��OLq�m*����G����[M�ҳ�-'9a-����_��ۘ#�,	�aAs�ʤ�������Bu�`�/wi�L�?\Cg���2�o�w��~�v�H��s��Ĥaеe�K��-*<��R�Cѽ�V��pt4�d�j��1"��y�8R��gX�(G;���fښ�<i�u�GR)�����_(�w9�w��q�6bTa���0�R�ZM(��%��rA�����v�;�'�V�W5AMU x%����>�׎H���q�ڳ�g�2���9^ឱ�{�0��c�N=�}�m|S����R�(�^hq5}o�����[Y-E!��9�ܫP1�T6��a�y�bj�u&�L0�L�Y=��"�O������f�k������[1��?	��$躸���2���Vі�V�a2�a6f�^����V$9�����7d>� ����X�����Ӽ���������^�_ E�ݍά�pqO�6�A� ����t5�zA0��<��*��oKt�����2�!��["|�����S�sb0�*�I�Ŕ�O�J�ˌ�@ZjZ	�2@1qnD����́�('j�B*C�)��y\������7�L���U��)3L6%��eW邅@�/��7��o�A<�)���8��%�JX�:_yL��Ujy'6��pw�%�r�U��ML�LjB�
���)�۱���6�_$ 	��f�H��?ł⎓H�>[]M��I�En>7*��?O�}��+� ��z
��+ �=mO'�[8��2�	my|�00p�y�#*������N�SbG3Gvb�D��P�6�`l0�"�C0��ĬZ&�����S��)���e�� � �9_=G�5s;���vp�[3�A��C�ƣ7�w3)*ځ�Z���9CE���C�r<
KAp��S.��J���v����-�MYXd9#���Df�Ϣ��j+��~2�����k�3�Ԑ�|��W˾�7\U9�*d��\dkI&�[}��r�	'�4o�D�ܐ)�;�ـ �"�%@���(YtJ��z�>�x���	��Z�$�j�m�)F���r����1{�v'�kս�{l�R;S�^*�
���̸8?E�^Ft-�JiR�*��^K
��g!��pyT� �-H�D4-���*d���X�beg9�Z򚈡���}:�b��RCC�R��*<�5�6q#�&v�͖0K���a�-�"W������(�8�:SO������kafSr��<A %Y��$-/x%]0�WΧ7�L��M7��s��c�B���T����P��^�9"����cU��i҈�зЕg ���y�; �3oՠ�%��j�.ZE3� qm��:����-!$Q�0E�=�;b�:G�߬w��M	�@��]Jh��^�'u�t� l�Ţq-%4��]�� )I��  �$��Ekb��z`�HM���$6�@l*s$Dw�S��P,�JO+j*4�7UY�����^�E�v`�B8�TZ��^KeB����ϻë��t��h��%�7�j�[�%�� d
��QD �����1�_n>�ެ�
��OW��d8ű	��|��V�6���>I�t�]�޶	��	�_#�c�=�{�8Jpm �c7)�1�.|�b��)I������l��R;���^�� ��
���K��	�W8o�Jcg�e(�	&�UV]T���i���KXy�����<<�K-�}BY�k]�T�ίnB��p)bO�4����|�����~���:7�oq��xO�k%y#��DHѤ�U���K�䙥��
��z�b�զ6���`F4�g{�,3�w�3X�Q�n%��h��L�V:L�T��3����v�ş�y*����X�	�钐��6�dD;8�;��FV�bsq�{0:�?��L��#(4��H�bsG��VJ��O��K��iw2�2'G�V���Q����;p�9Y��L��'8�~���ঃ�S��Dh��,mR�6����������5A�K���}�3jf��ƪ�y;6�WT�>������C�0���i&�4[V6�n0Q�έ�)��mbt��/��}MG���`��n(v�%P�1��D�P�[C�
lڵ~\>t��euK3;��;P��՚��a�Z��&�k߇�6�6HQ9���^����1��d��/���0
wg��(Lѓ���e�ȼk�A�`=f���Tp�n����)Dz1��=	L,���3В�7"X�2����ʴ�[��`X(Ds5�Z�Vc`�����������ؔ`�hw�����?WLk�nk��4e����쉏��i���S���kZE�ȕ�^2����%s���3���y�!aJS��I.�9��s̊��/۞�}��f���P(����"Oj`�V+ﮋf*\\���
����Yde,�Ό�NQ�k��
L��;w[dA^y�?O��դ�\�j2�r�-�n1�#X�����n6�Y�8��c�
�"���c˫�Rxs��$���s�;܊|/�fڙ��}	� �]Ǭ�\評jև�f�e_��%���V���Z))o�Z@�?���S�=q5t�xI�����Z�`���������S\���f?�$ �������ʒ�9�q�<z���ǀ�,���89������o5�O�i������L�b�(�pUߜ�pܔ��-���:lq�xi��A1�[|��J�}�yB(��7v ���-�tM�p����L��+��;4(5�ƌ@T���ϯ����9���������
:xhȟ�����.�b��e����
0VŠ�:��!ڍX1QEA�\>�ix�(XQ��y��j˙��G!���h�x�T�� )��K.�#�)ΈqDt���'F�<K�޸C���������OZ� �����߱�k��ƭ��毑vx�k���"�h�цO�,вA&����t%������^��:2�B���|!�Q��T�tڻJY�I���[�M��m�g�UG='#����w������!��/l�G2B-5 m�Q�IW\�.e�F�
y�)�-!ؐ	�jTK�>��V��)X�8����U!���������g��<�����ZF�;��Q����~���in�|M(.�IOcM���Xz��d�*|iqҬC �>V���>�N
���Aa�m�Q�(�<NX�Ŧ��1��>�D}�x��w�쓬�o��ۙ�����kE�v8.G0В���e�rQg�{��TO��O]5�Xx�j7�1��~đ�q+�w�/|�t�l��1ִ�����#"zQƛ4�1=��t���m��8�,Tc�Kȿ��]U6��?=��}Y�c��z^X%��6�a��u�p4�=�U05�h�$^R�h�V���E�0�/vdy�d���2s�쾲`X?Zdl�I��s�`���y��S�"�d��
���8�O �`�_���w:���S
-�'������ę>��pk(}*a�67��}'����O���T�6V�����)X$/������3�P7�}��\�xŭ��a��j��E9Fu<?A���a=���=�+G2g�L?�+gS��՘�D�-^�]�$V�1�4�`x�a����F�Rd��P�%�L�Š�ph�t��U������z���D@n�RA��8��]��`�z������|"��;NJ��po#Ix(&�-�HTfs!0'�g��6׈�W��L���+('8�"��t����ЎT����<���ܦ?#@-
O\��/�j,]@b��y�īD��&���[���i��t�JԵ!*@�~�-��� �e�$νx����Z<� 8���Տ ��j#Wg��9�%���G#���u�+m&�0�]��J���'g�1ܨ8�Z�fѐ���7�R�O���f$�ƙ� D`�e���=�Vm+���P�WV�5VN⡯��p���A�º|LQ�g>{[|�\L=s�Vop��KJ��aTܭ� ;*G��K�mR���]�&�0�g���/DL��o)��3�r�<y����@F�
D��8X|3��k]��b)^e@˼�!X�5����j'va ��]�,��i�I�Y=b�.p� 0���X[�l�����l�'c�������Lo#�T������'�O�8���y䡏�{�y0aj��G�Rmd�W�!p�F=@�M�ծ�S�X1 _J>f(!p��#2eb�{���Y�Wk	>��7�w�&�Z�����L>1{���ƪ�o�� �b�eBS!�{F�n�6V�M̳9�e�|����=ŪC�n�I�����@�@a2�;��̼k���m"?С�ХRc����wV��V��"r�޵=�m�?4|b�0c�G�aF�G#U�A��,�q���S�Wۛ�M��/ �d����EI�#��.8�B�q��ϻ���R��8��x����Ċ��@J�+���;��w�A��T��0��׍+�v��}�����{he1���|��rOE�~4����a����V�;z�׺����6O]G#��}r�~�3m���x��V=+чux@����U~@1�f29���/ė����o�s���-��%J��R�Oݓ0?S��R���8vR�����,��p���tr��W)�����rB��H�f�������\�@�1���K�ۣ,��PS`Fݡ����o<�đ��ۄp��Fl�n$����ч>�G��/m�p�k�u�N�f��Z	$������9M;Y_��I4\�_<Lw
�2P�~����N�o���'`6�����:��%��/:�R�#(�:a��S����M�!�l��r�|1�5�NzY}�ͰQa�U�@M� ��L2, on
R4���Ic���?v�䪫��A��վ7t.�H��bʄ:v�W�5hCw��3�а|D��A�$���[VL�ԧ��E2l���D��W穘�g��'\˺�!�c�W��̈`&�Eq�aw*-&��� ~o�5����z�C8���+��b%t��]�]��i'ׯF�:$�'!��9闂gܠ��J�i���?��c~"�ao�u��7�~���}����FvA���z�ĭv>)�
d] ���aJ6�$
��4ҷ��'K�$��l�c���h�J`lR	)���˵7���1T��C!ݖ �ϫ3�Z״��En�FGo�N*oI��Q�j��~��D��eG(�1�M]�م�h-�	�sêc���u������Y�����e��,�ؿڞR�EU����޺1�(vnW�7��h"|=$�o�z��|�=W��N��ò���r��ñ��#W�H3�<:���!y�-p�'�&�7����溂��&� 8OJ��:�ퟎƱ�Ƹ���s�@�o,�ῄT�[O���Kq�]�=�R���l�lA&�=�U�.�?hQ���/�r�ƙy�B˛�Cĉ8U�[�?_r�GQV�¹܇��P�2���21����吏	��)�쑻��nT�5+��ɺ٫c!�a�Q4�tOf���B�e�'�aMFH�*W36�&
^�1Hf�V���/��{?��H���w1&�b�s�{9o��7_��C]�e W7������P����Ẇ�PN��SԌ8��"s�&D��'b7UOBN�GcX�q�n7x����rS��B��:��%�Ӽ�о�4k��Bڢ�bEO�-�1���=�0<����|C]�yr��
@g�m����*T�#Z[�HV�-��Tvb�ҏ��qJ/�����u�2��g/,�cZ�s�b�S�G ����j#�F�=�ȟ�ybz7w�u'����G�D�z���È[����;���äf��/����Y�y�Y�x�UF���{�{g�W=�V�0�(�u^�\<<@,�ڦ0�I�Ni��G�fHi_Y�J��JF��:L��,��wUE�
��������4D���^}&���j�~ԥ�֤�)_ky�LKZ��n}�Jc�CUۖf�O^��
����r�'�t/;�9:���1!�*�+-@(�$t#I�\`�'�;�����%��|�=������z����}V]c���2=�$aZ�J�1�(TA�d��v�}��%y�6� ����U��@�a�����㾺�r�tF}^-=p�#�O>G�������#�<�Ej���,�h��rb�Y�L)Jo�})��| u%~�杨���|m�0��
�(J���ߪΪN���qqa[#͙|�e�
�x>���CPK˱�e�aaQ��?����Ļ꾩%I-=KvyL����$��)�pF&�11������΃�׭�q�1����,���W?����΄�;��0�X���r�p��9�\fƃ�V���4́���P���D������<ر�j���r�.��l�`"e�Z�}�@�"��,�XYRГv���aR�T�.�ȴ����R$1ׂ|` �d�����VP�ߒ!� ɢ�\R�m�\�dW�ui.m	��&�n��>�έ��� ���De��#��OK�ZdtG{KVy{��3�xNƪƆ���64k�%Y����fS���|v�2?kd�A�� �Ƚ��d�����S
\�E
U*�
�9l�uBS��r̦�i��~��hp��'��{lz؟%�9����T�5.,�դ��HF�g�?͙Q��S-
�Q~v{��
0X�<\?�,�_#�]#]��]����2�?�ՠ"W9a�
�l,|�縵�\�.��ct�xg��,�*ж������� D1)�����h�E�G�i�*+L�IZ o�L*��ӔKf}�Ť^D�1�����|,n�m�Zڟ�s������}���<����������k���>�'<��> :�Zu���ŤU�̭I�Q9H��Q�1�?6U3���=�%$Q�C���r�����r>�JH�I�b��O���&����u.2��:)����D���9�����H��d b� uȄJ�6�>����Ў������30��tx��������t�^���Ic������if�xM����IS���.5f�	�֊C����
ܭ:��F���Cl:�1��8s�=0�	���^ya�ϝ�*�N�^M[��LP��C �=ד� ��x��M;$�Zj�5�'ƃ]�M���Y�OV4�}��ۨ�F?}h�h�Xʍ��J�(��O�o�RѦ�C���zr��-������,�c�Ȳ������#���a	i8��^�����Û���ʧ���-ۄ���� �~!<���زJ<�Y�&C��cc�D�D9�,�;j�B�8���+�5$��1 Dbxf�Qj�U��P��E����C9��zV��<��5s��0��sgK�8�ebw����v2��-e��p�֔r�p���R��y���c�EX��B��L��:�!�(VI%��V[E|ˏ9�Lz��D��͙�IWk��ϴ^c��Og�5�o�����
��ǺY� �]�<�t�oT�k�loX���<	XC��g��AM9�%9k_�㠈�ԃ;5�´�-/3��n��ǫeq������J�Rk�y$���zz�^z�vXカV^C��1!�V$��z��`'@�V�����	3�w$><�f�|��W���UF�XL�﬽B�B%ʮV��l��ORN�mxF#�t���j����V= (k��	%�k���|�,ҹ��� ��:��ZV&��f�qPG�b�'0��t��1E�VdTV�-Q)M�1D�. �P�T�}�n���x�s��zh��9d9��X��cL3=笂M�V�8�r�l�+s1<�D+��B��%/UP�f7�#��#��F���~Gp����~�X���dU�D�Ǒa� )P%lN�����v�7�ڋ�㼨R���xBn���Y�����l/�<p�Ϳ�
���e�����X ~�
�;D3�C�~o7��֪���5�Dt�+f�Ɂ�����ߪ�6Ƞ2���9����{IF�䪑z��\��ˋ~�c3m�3?$y�PP��z��E���5.
�Ĩ}o� hJ����Q/S���R��oH�p��!\���#����-б�J,��5������K(����Ȏ�_g���a�'GFZzL�3�ZV�'0ͤ�B.�w^?�6���|���H����U�|aLNO_�33Ʊ1�$`<��_#�d�LL��s�(�l����1��Od���~џM�Z�}���P�*��Y�X�K�ք_�;���Ј;;E�W$A�j<����T�Fx�,1؀�"��?Ē���Uj`�\�PIܱHo0+��e၍2(0z��M*�OΔ'^�:���.=��q�;P��Y�Y+��E��Jp�����R���@l��u�F�R�@�gUH��0I��.ci,}מߋ~N�[�IOϥ�v�<�N�d+ҮHU=<��C2�Dޅ�#��`B��Ԟ0s��x�]����>��Խ䏥�AE����B�&��Bi��'t�u"�0�wί�-Q�u�
�3��O���Uaw�M��cq���q�n�b�,o�c;���0K8�����M0x@&�0�6/�k&����КFu_�X�yӓ��@���i�ԣ����w�*Z�t�a�Ջ"�a5r��P�3|�M���3 T/��[~��Z��5���'K�Ԉ-Aֶp2l���S�]|	k�'%|����4D�k�Vw��M��ul��C}"3@�c��n�M��C`>T�/�4�*M��9����;�oHGZD�Ĕ���sOC���Bnv5a}���ok����"�+ 0�>�ku���ؒ+�_��es�9�]�(o�}C��^��s��4�L�/�u�cg����d06�FZ�~�ց�`ȼ��ۘ�;������ �,��GgQ�B���
~w�dVm&.�2�6�Hv�(�ï �ɬ�ωc��_6m^������<��{���Иk�__F5����:�	���I|5�ÙK}c�f�;�\����4��|�\��Ύ��,��*��^K�)8&$�����֜�f������ԡ��4�?�L��4���O&�&c���AcP����������3��+���ڭ��xLT{HF��$�v���L[�z0E����4,s�/``��f'▫p�+�9<�D�j�l��~4��e �X%��GB�Fpf������v	���I���u?�ZF���Q|{���P%�E3��;�A�xn�@3Dt�@"-py�o�!�;y�����;��t�	��������y�IZ,4����P���b(L	��5K]s��Ƽ�R�)��#t�1�Kx�7��`�r�5**���5Y\7���V���}I��˗�he��xE�Q�~��d�iF9J�`��p�_󊙌�Z*����#ݫ�|L{|���˕w��U�W;d������<ご��Il���A��]��W�5�Ih���5>� ���u6]���L����j��H1!2�q��m�pΏ;JB�dI�7գl���Q�C��jq�@������W�[wY��|2�`)��q��k̈�U�C�ڿ·�Jg�4$[@BC�
a�W"v5p;��UM�fJl7,��q	LEHd�ĺ�ː��:.�xI�����n�#K��!(��yD�&؁Ta�}�0MGʵ���#�r�Y}�f�W��"�(y鹇Ԇ�A�r�sl���Z�6�Y�L!