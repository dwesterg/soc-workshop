��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�Z��!bJ�������z�_�ZC��=}y��a��"la_��u`��(��<ʢI��n��~Am.���ϼEAY��$��Ms�_jѾ��Q�^XP����g��P<������M�V��)!9�R��>J��F����x��X���p�$�Ws�u���d�Xj�U�!�; sX�F�~0�)�?���\�߸S	��Fb�hX��ǫz�Ci��+,'=?P' Y����p�R���A~C�1a�2Se��$oKI%p��f�D}yC²t �q�j�j�� !^�y�;���J	�L�a1z�12��<�/o��w��ð�����+����--���;7���+g�����g��cG}�fƯʉY۬ ����y^N��W�h�4����e�8H�'��e)~��RUu�t��#��յ�4ǐ���#x������K��W'
��h)d�?�{��οj��&s)�RG�
���4��w�*@���SCo� �Y?=�8��v�P3(x�Zk)���ŗ�ww�m���9�\ۘW�}:}�et��*
�fկ�Ω��#QnJ��	���$b�Ш`�>����^:���J��~	�$/��^�Xq��E3������L�e@H}��ahQ���E�:�VķT]����q�>�/�-]�>W?�s�	��=D��@��ȓ��̜�w՟��AӺ�ȓ�=,��9���6��pk�IfYt�L���߁�Rx�L�;��{�=f�R�{#��a7^��2��o�U��<�R�wT��B��9��|[�	�X0"P�:��9�U�8 �����7����4��]��g
�v��J�$�����뺭�%������jT免�3ɘB'���^���Y�L �p�2X�#v}8p�[W�
��3����<ɶ�]��lмH�=��M��v�P�)5�&+%�ҋ���b���ɧ5!�x"W,���6:�	 ���zgw���U�-j��x�M���9@̊/]����©Dl��*�d�>֤߭��
�$dJ[��-������W�����oY8$�1�6N{m3�a�t�%e�)ݞb��%��v��!e%w�x�⪤6D��.O.ק��{� ��{+����2�aKP�靲��g=ҵ� Y�#l5JH��Yʧ�A�8Q~��z�(�.ƅ��r$vv�pQdD�2�1ͩ���<iq����i$V��В-|\/dt�?q�"Í�GsR$�U:h��#�]��4�H`��>�е�Ѩ��y�Ư��h3=M>t�+
��X������^�t��,�lOh����챒VSMJ􍪜��A�2���bd`�y�z�Z�c���C�����VK�q��I,3��<pQ�Ir?Ga��'���C�L��{^�}�Ј��GG����t�%OO�x���8�J"p�b��&��4��랋��e�7׵~�� W�����1F��_#�`�ED��j�(�ߣ��]�|mp]��wm��yM�&H��$���̹��-b���W@*��AH�[���� J�֠:�%��������$��S"[����z$�����G
1���P��WXڤ?ny���v��@�՗��B�S�:pjѡi��}��W�xxP��!������æhG�t�"AV�F�v�0$��y��)�A{�C��h� �!�9:-u��7�wn��P�گ��;%.��p��8��`��)�������[h7��~��sn0`��֢ܞ��.]�e�!�|�	(ـ&5�5P-���(�u{��^��(�̙P���7 ��}�l�L����T���/9 +�<
�?���PY��w�;̨��Z.��VsoTE�%�f��s1�5'E�w8�W�v��cҟ}^��2��j�)��ȁ}ݱ�Rt���@%��b��H��q���H3S�hp}�!y���6�H�v �u��}�@/G���Q���l�x�UP�`M��
I�3���������a�s+K�9LBᎌ\���<�#�!�$z�NFm0۠�`ɘ���6��SCj��w�m���p��Y��؀��R�aa?�Rת'~*m����¹߫j"����� 6��k-4Hn��A~�dX��qw�z��Zw� �30;��hK}�iV��Pw�M�y!\)3�{����ܬ�'��c��D+�c^����Y
g�	7�]�������jmC�7��m��߱N;��������d J�p����9'�­5ki�����H�&v�T��oRМ9Z���$�