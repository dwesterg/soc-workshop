��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�Y�CO������_L&���L��5����V�5&	5��
2fOths��;w��p��(����� �c6ْ�}���"c˳oA[�:��yY�]BLg3�Yd�G	��t��I�?~�f�R��R��GN�0�@�Ž� ����Pzr�TM��A� 	�T@�M�c�yn����l��g������� X��/���ro�d�$���c��_��`�6A���ک�Wum�j}îR ���,�����i~D�?���j��V�O ����X�G��H����$��ۦ׷<�<�"���:8Z� l+O]Rc2�,T��buS]�)���Gl����]�(/}�Sw��K	>���q�l�"��c�X���oq�p}!�Nr�t��.�N �eb�j�Λ�����E�,���p7�_�"�qH߽���^�O�s���?$1�GH�l��\��Q`�4=<Ť9Z+��j���@�N��E��ʚTjl~O"�O]1�7���pMs״�8C��C���#^��m���%.)��Ń1�a��Օq\���wd|��j�}nE���3cS�Z˾���W�lgڽ�ռ��fH��4�Q�̷��\�l�N��tT��F�@U����7�̘pЋ��|��y�)�ԎnF�Q!$M4�I�ꭴ"]�ڦ*3�`�>_t�l@���+ZL(����v7����O��l�����zԜ�b�X�|�,����:c�p��|R�&z]�c���=870	ȭN�󖟫9:���3�C6O��t<��U�����:H�uS��?DX�aG����uM�!���k-u������v+y�J���M�X��^`�֑�N��2�,<����,��j
��_ �&�0O�0y�����������w�Io��a��@2�~�	��Dx[ Bu}��fc��Ez����BM'V���@��fBe�Jy|��*���(���5I�ڧ���� �e��s����J/x.�.��S�6�S"�L:�(aȌ��˃���u���,��Z����`�LI�P��T�Kl�0�	!����j�`dI)Т4�s	�}�1N�C����
q0����92|�6����Q��R����� ��p:kʻ��~+���Փ���PU��x�B>��I|vtR��%����E-%囓FT,i��SӁO��|�kí<��*���f�!��)l>�J�J�܄C� ��v����̨��^c�M]�1���� �AM����1��~д21�Sh�r�TҸ#�r��
���n��9p��a�$&��ʣ8ۘ�źB
�?U:�?����ٔ.-�lemTӇ���,�JU����S����;�����B���SeD�J��7� d�.������m*,��&�¾��(fS�>T#j��E=�2NKjt����f�V��7����n��?�-bQ��qq�Ms�QK���D�(y>���u&�W6,����H��I�$0�{�~p�cE�/XdK���l-X U�	e�� �Q�`��3b_j/���-T�t�)[�K��z������ ��:X�F/�-E]�=��O�d�T�����<�~-ByrK�q2�%d�I؃��-������(�ڇ����U�	��V^���nN�(56�����(�j({����N��)5���Z��ўE����[��<�8��b�|Y3�H���'�_���?��?,�xUT��o�b�2��؀IEF�b�����z��!�I�Z���~�������o$�܅ZC�n(�Y9�_�n�\�ܬ	r����v����!�:���>�	w�B���iD�f�y�y�n�*�^�+C���Uf�RJ.��K3\ż�o����ŧ�֋�������W�--#d�p��)~U�k�  c޼#���$��TI�Xݣ�-#�P�O/B4l�� �*�ɆѪnup�	�7n�M.bn?��:I�F`~���)']�>�Q��ٲ!�9u�g�S^	��Pa:!��2���b�LIxm_�lי�N7�,����a��ML��+�������1/���Y��m��v��j~{amd�"QG�|�T�1yv�C����� ,w��Kü7}Y	�c��M4_�'�æ/u�"�X1���J��0��Dd�͵A�����!z�����)�j�̦�f��Ux؝{��:-QV����lO�`2��+��ޝN�C]�*T���_�w3_$d	*ް��ks`I.n{�q^����al�s����8c>e���x�9T"<A�_��r!�����V��kDj�`�h`�����,��/���'�F=���7�)��j��]?d�~�M�_�
�[�����q���RU����s���f��>�sV�k�� ET��\ҵ�/B��*��3�>1(g{RA`6%�	f�ꏍ5�JT9��&��,L-k�ϓ��0NǼG"����Q�)y*e0�������J�ҏ�*�	�IC��|�D�!�a�|JF3ҝ'
X�ud�dV��ꩉt4\����r6~meo Mk񒴧HG���+�(���j�	�@]�|y�})���M��>�%���Tb\��[<��o��@&�ȝ��ŝ���M_����=]v�5\A��"y\���O��71(��w0BP����lm}�ds�܍j���"U��^�K�pB�j���KF�����?��.�,m�ԕ�������rɋMoby��E�����T�?��r���QP7��`���n|M�xh�E�4�'T���d_X���Vv�_ቊ��Ճ>!�Z��1�=�^�e�Vj3=��l�V��?��Iw��_`Z��b���S����:�>�i�� ��ᗋx�"2�P��4�8m���8����b���)]���TI�&�Ujߥ��ii�v��ҽ9�!�����t�ð�E����5l*h��$U�T*�9��:�����)�`�V���lv�8���c"X�k_Mn
�Hh��}�1������ța�j�][�W"��ŏ{>�@����%c�J�k�O��y�ˑ9]*������;a-B�8�t�i��β���V^��Tx�9��#�je\DP2y��;�A]n2➖���*�����ts�=<~�I�onZ���f%��=�A|�@h`��X���HV�����ݪG�|����f!	��e��i�djs��#R0����o�jxO����\nf�7( 0z3�]�1�n4��m!�d�ɻ���(�0}}�f��)vu���jW$�$���'<"(���3��Xt,1V�aC����^�����y¶�M��!�x:kE�%�f6�	�▥:�Y7�zr�Jt�\K𣎴z��n�R��dH0>l��oau��Y֧��h�b?[h���g@��Du5��h\�tڴ��@�F��ꋛ(K�C0�!��}�!ڤ&&��?Հ�u�A# �w/L�Eo�._��&�L�2�&����b%�$e�bży���?Z��J���{v嫦Ohb�u�ֱZ;hI텏RP��H��p�Ȟ�/�X߲���"�(�T��<����u��i����	>�Wt���L2�%�;��>�~n�<� K�]@�d�J>0ŊJ��"{'�$@��Z*�;�
�N�2�A��r�tr���F��9^�E	�$�G�/s�M��=������8� 0�˖�.H��W��A���!j�^�I��a�_�U�y��Uw�����40S>��,ÑDګG�ś�J�(�:dN:X��i���h�|�6�v���W
��xi���u�xd�����v4�؆�ʏ�������iK ��ךmڀrX}���>D�ﰿ-`�����\�[�v��~PC�b��1�!�!�KՓS�-9����'���.J됗/uЄ�*%�N��J<׉��LV<e�Ϳ��%վ=�_��������GF�����'�yԛ�B�y��a�K��a )��_X;���F�Cyq�B�LQp��ȓ����x�&,~�xe�jǤ�Y��i�H�y�>r���6h
���B��ߛV���F00���x<��zط��E޷|���
lK��dL��*A�WL�B�n�1��s�w���������,��J�h�w�M7���9��lS�I�t+�����"l���9��?������%%ɬ��*�UtTo�a�9v��Y#��@��q��#�����\�9
d��8^�mx+9q�c�=�M[����F^	�W�����ȯrf��S>*�ͭ����ʹ	tZP-���Qx>���&t������<�6��'���N:޾4���)ma���)�,��}qAqچ���sw�C����!%��"އ�)�~]��!��@���gGGq$�z��
���<�/��my{d���N�z��� ��%i�%�[c�(ڃ��p.CJ_F� ��l��आ��C���@�k,x��5�g:�o�]&8eDΏyN���-3�c�\�Ή�̰L�<?��T����]�>�g��ʾ8�̋�v���+������qn�����6$�T�ƙ�|��J=��$n��6j"�!�E_5U�!�E3���r�b�&�_~�w��	����م�Ǵ}�h�?bN�ۦk:��(�?R(��V����5������N�� 5��H��� 9�q�B������
�X���?�pw��R)����,"�佬_�XxѤV�E����:?��r��i�lz����G�#�96 Ѻ�N�ɝB-�E0YJFW X�O>�5��gS����0D��k>Z�:T���d����H������.6eG�7��+����J��%>��j��������!���Ǌ6��wj��@ޕ�J����ſ���!F��Y�SqJ��T��z�#�%�7�X4�[�Z�B/��P0cr�+0<��]b�ZWy��J��[��?�vA>����F�>k��gE����J�]=Ŕ/�z�7���ի��hS��a����@+�9]-O��#�=<=x��/��X�,{=��I<�G�;�1��Z��fF�.6".�Q-}(}��l�0�^���̀�>�j7�w<��ȶԝr�?x]f%��8Ҕ�§�FĮ��y�h�I>6�>��$bA����\T"߇����b�F�$�-;����?�p �	���㳎#��4iH����L�~c�k󈔡�W$�Rʡ�E7|����*��Li�{@lWQ��.v�(�t�6�9�R�o�_-
��|R���[~��«����A�Ui�ru���C�р��LD�d��_��*5��D*Qw�#Ӿs���\䡠p��ߒJ�0��}֣X$�!�������E�l�d��2������)����/�������6�3���������G8K���������#�,�&�v��s��.e8d�]NB�ky��𹜰���U���d��۰}�+w�h�*A/���B�Bu��'Q3����a���*�as:��JU��Iù�]��R2�=/�ϼ���0rXpC72��?x0�6pm����T����Bd�PB+�y"�} R�Cc���0�b�����V_h6�����&��u����*��N𞪨�s0�q��H�BE*�G�E��`�u�:)��~K��W��15WSŏ(���f��"0( F"*DC}��)�	3��kW��DY����de�a4X�Ft�nn��kҴ���
�?���%��;��6�9Ao�=;���4 ��m(��K�zDؔ���N��z���\�0.��T#���Γ�	7�'U,��p.mMA�q.���όY�_j��JT�2ha�{5��X��J�[N5�t�D>�Y��<������T*�@�$������x��d6���4g��.'�Nә��<�� ��=%R���#7�wծg���'��|ؗ�~;֪��L%l�Ή-:8��]Ѿ<�,_�Y�VX�Qƒ������zT����m�5���G��g�^�̓a��g$�Bh��T�t;����S3�hJs��^�n۾	���D�$W��2�E�EK=�!b)t>��$��t�b��7�^|�R�;��ʸ��D����ջ�ӵ�P��(Z��E�9}��J�΍u!ٌ9�i�'7���P��PH;?��>V���;�:��v�ߒ/X"z�BMn#�MW�بS�� ˈhɎ�ꉄ?��O*�7u�>Y���)z8m���ō�H��cI��IA��@�~m��v>c��oX�:><(ًr@j���Q�hV+5QxO	aZ�{m�uN.����Ƹ+�_������?����H6E�x:B�.��l]��s�[Š߁�h:������=�"�h,�	EQ�8,=˺���'��Hh	����z����g� Y��
�F4
ر<��wW��a�;�MԈ�j�Ďډ��V��#��uۃ��u/�:1���́ZtP2d�<7�jۆ�|�����>��Ɋoi��c W��4z愐F�I8��7���:Wz}���D���]�`�a_�R�s�v�������f�0���r�T�i��I.�(JI��,]^#��[[� ���c�4����#ݷ�Xi�x�8�z�,9�c�n3|�8��"�O����V/,䉺�3�d��Ai�sn���~���@��xrc�T�V��Z�_s���ьш�l��������g��JrS�&w�>a�C�߭�{���@��i,
���<�՗v�!e������ź�UU����8��f��_G-��>J����N�ʩ�t���c���y\M��kd&J��py6N�@ K�v�]ӱ�3������)^�M�|D!���ܺ���ʏo߽�Pg���ݽ�9���6�¨n���>l�Dm�AU��F�7��~�T���D�ttu~�g��*��-����E;:��G�b���;4���5?�ק)bwՉ@�l8?�ܶ��kH��8t#���ܩ�B1�nLԨY�������!�!����h�@�Pd5q}�K��]W(Ρ��^�,�G�0cGxmdm��!|��xP�jU)	:�e�hks���������y��!Q��K{��&#�H<u��8��[ ��W�Ō��`�U��o��&�uC,2Y�M��V�p�ɜ�"l/r=i��eF���j��up��:�4�1��B��]�ޚ��
����. \�POm�*�J����5�Weg9�-P[�s|n���A���ɯ*��T�l.f�?��Х����ӂBd��!�'�������l�`�5�T
j(%U�dQ�$r6��A�(;�:��~"Ki�fG��a�����v�R�h��iy��\��]6��~O�GZ�bO����_���(㇊�ՎŮ#�.�?6���K�?�|&z�p�w$��M��h{�܁�3� ���Z�7�K����B^�t.���a+��������o��!�������CS�rKv�G���,!�saW������4#�@M�\�mz�Ny��R}��T�/|�rx䠦`��,U�s]}���m�p��+�����2���[��!�UO$�#<8��fd�0�-^�tH/��)I��;�l���k�U���|����Ѧc��[DP �OKM?�oyzfd�Ke�Q�ho'��{H?��𳅓��Zq V�5���|;�]�Z�`V�!	�鈦��8S�M��t0�nW����X����H��M���S�h<}+�Y�(Z��g=j�/�I>@��^�ף���뛌4�e�^�
F��7JĖ�Iz�'Ӿ�ه4)xO�c��XԾ���쑬�KS�9�U�x����z�nݴϏ?��Rm�����@I��%K���2&���D.��ӗz������P��g�7Tq}r��Ջsq(�h�p�w��Xm�ۨ�5d�����JDst>N>%��:9�$�Y�4�r�����Y-?(�Ej�(+J��Bw��|yM���˯�`X�Fo��p��
/o��s_�s�L�X���[%�E����\�i�ςI��I'u	1?�~�"�=}�Z=$�]���#c8��i\��i�ӟ��\%���d������5�;ϋ˓�J��l`s�ʹ�	��N�1[�����(5���v�_�B�وE��t�ս�Z�CC���q@�"ae(I(�(-�$c:�?��w|��q?���3��nU��Ѽ�a������[B�wޅ���9��z��?jѕ�s�������O|s�S�6��ϣ� <(z���hN ��nG�;����Z�}��'�P0�C��	v���]ML^���i��)�||�9�
^�t�� cC�B�RA{PUt|)�,>k��p>B^jSv�3#Q�����mak�`Bm��n�蟟�*%T4�O�\4��D�U��9&�
.�9�ԓ)e������P}�,<O��M7A������v�(2�뢏<j���*0�/��}�>����2�
8P�QZr��L� ���OX:@������sZ��o��d��W,�ʯ�r>�S#x�v���~�t��h+v�<�`jVK���x��])��J��G���u��䉰y����"{/��� �O��gl��lK�HA�=���-�gĨ�o�Zd�^*�:L)����{N�#8�JSȑvp[kz:��y�A\k�������g�*�M��=�w���+��*���C(�kΗ�Q�Z0��M���?�Y%
���N���J�|�Ex+�N<���ABy�M���vL҅��r���Bs���{��OJ����/�7�<�7�����53�ʋ�{c8�3�ة����{�	g��t���r�u���4'���9��G��r���������(f
�enf���wj�FF�LR{�0uVc�D����7���
 ��]��s�*��q�s��79_<i��e	:�M�b�w�/�4���ā4K��{�2.!<ٽ>7�@"~%�������g�=c�T����l߁mw���GL�Qnf���6�ThUᏤ�~�捹x�*���H�#�|���NGBY��f��]����'y'��#�Rl��?.��?L3&F6�>c��0��YxP֥��u�մ_�IN�!�7�H�Ӗ��:!_��F`zW��f�����zF�MՅx�y���?.�>,� .Q׈�Z�"HFc�kl��E�Uyf5�cne�Æ����mq��"��Nj���b�yO��f���#�W��,��ҝVe�zyr��0��	���l�i�kM�D�4��;�����3Vu\�p�
:`O;~�XM���E��m���6J�_���"*�c�b�I�i�ksMю(�	�l�cqF��ίx����.�?y⽌?g1H�jD�DN��GȢ�i�'�\+��Ϝ��8�*��>��Ř��s�_gaY�|�O�|��	�n��0D�m�w�����@`Oo����#����;�)Z�>�:����J�_�mN��ղ�mKc��|5�^�C����ȥr��㷆�D�k�F�p���$O��������ŪX�8��%d>��ܸH^�� �%`�&�T�}�)��[00kz�*�����l��S(�����b�����Ϻ!�:���r� m��U�In�9�}W-����#f���B�A�qs��?���C��Jw۾M ���T+֑�L-��R��@4�̳*�-��d�?�%�y��MNr��h���K�ёa�s������D!N��J[�f�"����Ň�K7ǐ���TE��?e���;$�j����YŐ9;��kI-���ܶ/�ݜM�J1��B�+��Ϣ�8\�z*�F���@6�;�'�,����N�#�b�s}�w�9�����N�In���oN�~:_f�/�����"��A��U�«j�	���$>�,8lӲ�	f��GRE��k�&��:�]z�pp�	(I�N���r�����n�9�o6�%=Yo@���?�A%;��WO � �~']]�u�j����N����)��e���*�<4��

Qd��e�聓7�N��R�b���.��1Р΄T�t�HÈo�O:�݄_Õ�.�W�MS2�^��h��������s�;;�/@XY�XFx��#c����l�����|���{MF^�/^�����Z��T�k�]�t7���m��S'����t����0�Q�C�s��2R����?����n��r�k�w=r�&�K9�Ab4%E�V�͘�l�hs���#J5�i���q:E�6�����!qA����<-/��2�"{���ʗwks�)���\`��z�'	7����vTu^bJ���w��Ɏ*
���d���=�b�6ժ�.�1ۣ��@�ԣ@��c�)�����dWI �h��C}���_Cf�&P?���y�Q��Di��S
W�f�5��~1*���3���?����9����}�6z����я��x�y�O��m$���b ����a�mǡ�M�\��~Aѕ:�9y(	�7_c^	ۋ��AIgU�r���m�1p��Y�4tb{�w������>?S5��"`�Z�Xt]W�|����I��Uf�k-BlqS��)B�4���P@p�-��ko*H�ĩ1JB�L�OC�l��0�d#P�A�T����;����a�J���gz��M��n�(���O���S�u�E��"�|�U��.V���݀��R�K�6��8`�F� 1�?��F�d�5j]Yk�3U�?7�0V����=�^�<L�Jt�����/Wd&�V�#�cy��1�v'��:R���y��!0�����t����k:u"�_c�7�c�˲x�;S���{Yކ{M���[����A�,���M��݊���8�k+uvaшL�(M�	���\/���i�-�B+�����"�w��\c��ڸ�y
�
	�7d ���$�U4��K `��6�8�(nj[�)6W��$�JV��J֭K3)��ݹ͎4Fs6��`�]Y��K��#���^�Z3���j$��{`ʬ�MeB����҅ڒw�(�D�����R� �zpa��_si��|Gǹ�0H����� y����b\�@��ݩ�)^�{�t^;��{fY�ku=U3�dH�u�PɊ�WET!x�C^�R�>Y>�hh9� �AS�!�\��J,�f�>¯�	���ä�n^D�D�"�;�QPUf�8�OlYL��WwGA������m��!�8���� oJ���݈l�59|���\Lx���?���A`��s��zع6�vQ�	�.B�;�*����#6���˯q��K߬�2Z�i+@�	z�k�����^����ubTr��΄��D�Fz�tv�H�!t/����梧&PD�MT�ŋ�B~X��xM3R�A�l|ԎW"�/`�&i����w�O���<�!�)���Қ�Ԑ���^�����{c/L�4����L7=ď�O���O�%��Jx�,�0�?M �b���T��SL���pL|Η+���o2���,Lw�b�w��G�G��*��0�IU�˳{�m��?�	��%���@�-�(\���EA��9�x1?/�}��eae�F`^w�>���E��DՁA}Y݇BL{\�oMo�U�����Q�Q� �G]E�<Z(�L��qQ����;M�|1�A��S�d��a�KȚF�M��=&ʅ��rM�;?�jD����n�*��i��Ab� �&DR���D�}��2$��ǵ��t=���ه�@eV��+6U��m�=�諧��נbU:L�8˾_�[bb߷#+�y�<�6C���d4�F,_K�k�-cT�9Qw0�-��i K;ahjF�0"��ݖf&27������ �hjYt�H4������5���P���N6�#4btl�-�e�4�"�*�&��>��D���X��l�Y��{*B�*ݩ�b�=�o@/Μ���B᣿'�L�aS���[.�cr����Q�'F1sn����Ym��J�̥��'�$�����=1tzY�t�|���t�|v���?ui�k�q�c�
:(m�D!8����GW�'�gH�V���8�G#�ϡj��F�WiJH
�9��`�U�9٧��Y����v?V#~��6ީ�m� ?��ȯ����=���e��-�![�<Q�=<<�=��>6,n�DK񷽏^4�0T|n\W��ϖ���V��bo�y⟇�|��T;�Nxd!L �k��]�Cr�3�9��{�u���<:��r�q����2M�CL��� ����tvkE(�S���
� v�.W�x�H�,D��GF$#����>ݻo��t�#����� Q�.�E步�9���� ����;ȿ/��"Hqt3led�B��m����,����p��/@q[����V�1����$L�<l�dp��b�󉔚��i�/��)鲹J�<���k�S���w�ц$����Ͽc�s�D.�ڴ�P�JG
���p��ކ�������v2���Z#Yf*�*��\s�i3���Z����v��,��TH�>����t*P�~��M����Y�e:��0u����W���!������C0"�r��^C2��2J����T�{�lW���WГ{y/��#�$�|����ߑ�V�R?��("��ҞB�pI:���T8u�KNT��F�:�媡�+[�����N�TB���Қgf�.�?��A�?��;�:��R�en�t���K��z��Rxt��K���!VhR&��}e'+���j��@ �B��Z�rSk[��W��/���'t�q�$���+� ��_ ��=��$~la�4��2o�Ԕ�FT$v�Z'�%ӡ]��
�`�aV)TZ�!d����.N���������|lE4uY�[�=Ab���� �0�N&��(�c��p�Zg�[I)�$��&���ξ6�f����$���1�g�'�@{��|�zxp�{"$��C\�sPY��Z�Q��璺�'�"��z�~o�O�S 4�	�V�EfC���sU�Z5��61�@�%ŕ�s��^3��O}:�L�}'_��v/nu8��=�,hGxs��;X�<��Y��wDX ����:0�[j���;;d�i�)�qJ:��.��/Ԥ:@��6�<S���m��Q|���b���%@�T,M�k�3aK�{������`�߳�}'�2X-d���2�����:�J��4����~�,����[�n�[��L���~��b��a���4����n���ayoB����s�y���U\�BK8!��ňs�|�*��� //���عr�	��-namW��]v?QKG_����9�lȏg:���8�ף!H�Q�r��+徯ƌ��𒘛�����Rs��RoJR�Fg!]TΤ��_^��O;8&�V�A���Ҍ��xm��֎�)<�[����T�v��xm�3���/Hh�����݋AM�1��}s?��B��Q.��$.�^�`�B.b5u'����U^@D&BhQJ�2��,�[��4:=��p2�^e� '�5?��>��A�Ap�W_�O"<6�F����L�]MH��B��̉�G��[q,y�E
z?Ņ� s��Ig�C��"I��O�xx����/�^$��)��K���H�a���~��~����yQ�"�@|�V��K�*�zR���Ag��3�  �r�F��*�w&�םF$��t;*��
��s/��j���b�m���4��7�]��~�ز6=0�³Ϳ�X���^)�*���p���p��><��ܫzp}����/ɛ������m|�t�ϋ^`�:sV���|tl����§f�fce�+2��D�C�p3�	׼��r���e����)�)��Z��%	.�q҇��݀C�O.�w��:�V�-��W����^����.�sJ���,��
�b�D�]3��(�tb�0�ٛ���|��*0�clMm��U�_�<|h�R��� 
Nָ)%�<vem\;q�Ơ-l%�M�R�Չ�5�/�ԟ��dK��K�Bpױ�������(:r���%Ib~hpK� �$xY�T�m����ptQ�Pl(}>ׯ��#Ll��+]���r<�[����:u5~;v����Z{B�}쿮`Q����}��c��^9$ￔ�zK���.-I� �0�҂������p�µ�E ��O.$41�]�ǲ�"���fGB�\�_�a9�6�7��jdo��C���]-�n:,4�L��	���dY���M01r���خ��*l9Q��D6H� T��@���4����ݘ*�J���Ϸ��,�6���,a�$58t��im%}6Y>�r8�r�!�Z��H76+?;{`�S=%���*�R*���G�b��ep}(�+V-X��y�gCX�8xG��X��#c��%s64��琔����3e��4��"~�q�J�����y�n�E$�S�B=y8��х3�+<}��T�c;������y=Ƞن/�D�֊�� ��wC�)���/�a|���!1�����<�����t�g5c��ڗ'�\�^�PI��>�:3`O	�Q��!:=B�a$�_��`Pd�v��D�[|����Xˡ4}�,چ����W�>=+c+�Z[Y<��)���).��"0L�@X��h�����E�4�8������[{��IQ����x�r �a`r���f������JA��~��y����E��E�]�B�%8~�e�ϕ�z�*�,rE���L%��(�jO�ۧ;��_{<��i��}�nVX�S<ȱwd��38T�����
�hCLBC1��S:��9�vY>�v����d}*$�*�؎O
���|��<�#��O�Y<N#�ŞD. v�҃&���J�|��B5Tk�|}&�ָ�rӚ�ճ�olU�M�l�?����B�uM�>]���Qg;�3��2�L��_���;�U��ͷ &�Z��-e�:
,S��|������E���}=���m���0��`���!�:�}G_�V.��{����֝s�����ɥΛ��V)���� �آA��_
��o<�����Qon����b�c���	Y�'}5���)PdP�[ٙ �S��#ݒ�K/�=�0�HŠ|&��O������+ܜ��
�=�V%�>�������޳s3�s#�n$D�e�02�nډC�!*�����E֤�sW �5�N2'i���d}��Ұ����~��[�zؚ݃@��
�؉��	��Vl�ZT�P�b����`��4�\�.�E���Qv&�T��Bo]�n��iB`e�rj���?�ldZ��5���e�-otS��X-��[.��u	<Po۬���2Sz�����lY\4�vC�4��"�vͲS3��<z�̊��@��H�����F�+U͖�Lk�\�~M�yP&?�<���NIr2||�<ջ@��}�66��J9ӄ�k0J�}Cd��"/�?
P'�5�' �jFhhR�������˾��=o�:q�� �6�����J�FԔZa'�a'A�XRA��N��=&�gD+���C�55oad�-!$n�3<@�IpaX;J�ts*R���42 ɥ�x���\���L�W��oi��R��Eg�{�5X�]�x�'`�3hǂ�qt�n��/b�#|�W5w@��ܙ�h:�%c
��*/��x�D�@��J��L2M���>X`	��%���W��9Oz����g��������[E���9Ʈ;:]z.�}�b�@��c�<y�J�_0�Z]j����g�hg@��2h�{�&�ٗ��]�\���W'�&'z��֭o���H�Jʕ�l���#ŋ�Ti���il��͓�|%���Q����9U�!�@e�L���r��'���x����<�ԡɶj.9��X�{{�X@��r��"_(A��S��ia�	�c�౻ ��§UAD���|+V�[,D]�>�!A9ΏԷZj����Zbi��z�����u��vO��D�ä�����R��&��Q�Fp���:Ιc��� �Ͽ#N��n�<�j�I��`Z���O2�B��G�=��K�+g�M��LBu�D���ߑ�U���'�v��e��p=cp�x�}� ���4��;A�b;d��\��~�r�M5�0ÃIK0}��O:1?�v�C�o� ��Sa�j7�ܵ1�ؤv�e��r��-�<wq�>��B�3N�S�������P�}1����L�FP�td*kH/?��m����F}Z�#[��RHͩ�U�,� �y&1[מ�o��+��?F������2��w/�3�{��ܶ�FP��48��Tvy�����E��qw)��n��Bq!�O?��Dt�X��S�Ă�����>���8�Á!3���[�?�D�/5��R D�D�p�^���m6���O�X�IG�ӴwK7n��]�4�Cλ����R�K�@y◧	����Z�~�`�5][�������C
g�GQ"bXBhl�5��|������}�I�X�z��]էv���+��o��a	Z��X9�_�G�[2��#r��"���1�JZ���&��[��ү��0�[��"��y3��n���ϐ�)��� #f�~`�1H�������\���� ��b��V�����E���I�X�y7|'ՠ��rB!�п�V�����Y�բP�����H]����Q������ȱ�J�IY��\W���g
*�GU���nvO�o�ј;�`���s�c6�Va�Tכ�T�����է��V�?;5v�7�Q%�����Jt[%��dg�b���5U�ɦù�6\��/��w�]�qq����
�ܴ��[���A�)iq�o��S�#4E4�J���h����'-X�۶�2҅m�Z�Z�'���=mȑ+9������#�̽L-��#����ǅ���)��Q���&���E�ނ$3������oW7;�m�,_���)V�#~o��X�,
��f��?���S_��KcZ��pؖ�
�`ɑu]�s��-��F��<m��R������E4~#�Z��8�C0
�����b^=�-p� zv;�V2j�a��z�-�k��T�i�h��
ҜG�sH���]4�8�k��f
9�vJ�@��q�[5c���F�
l�li��z���@Ƨ:�O��3�-���q�Ȉ{3�,��T��������@R�?[�Մ��qM�#�Mf��\H#/��a/�������;E�5�D>���j>�r�}�{��ޘ`��{`��mw�%x߿D��)��3��������P��/����o�v��w�N��iZ�i�4O��f�աv����@#"x:�e��wY7�v�a=��ԣb���Y(�`' ��q�P�bT��	��yYŻJ3v"ίC$�B�Dѳ�`7:p|Ց�j%A��(����@��=(�W��E�u���|�X�qI��Z�E3A�K�9\10(b�&��Qx-6�3?(D��@İa��IRȇIO��ڮ?��b:��Sd���p M��|nǵ��׍Uv&�ш)�6
%A �Jc~b�D�2��L��ZO�Y���R0WYl+��� ��ͥ�"��lw����Zġ�7\m�0�=��b����&�B��^%8�]OS�|\���\�y��v݌���9��>;�If(���o��&��h�ɢ$0F�0$��z�O&N� `�:V�������DiG�>v߭/�������j���v��:v��#D��A��C���?}���d �����YpZ�}=<���D�#�G���[z�4�X��:�>��A�X���4^��oG�7Ţ��I����[ܾ��{���Ea/G����	9��XQ������J�3�O%�qS�,��NC��Q��o���@�2#�T�5�N��^�ͮa��S�i�j���U�ry�{��eN⿏���E��V�32���C�A��� 7���(��g[%�G�wP�un��ئN0D�|{:�0?hD��N}���")O�p���T�	AY�Z̙�lJt;$�6�G�����|J�Se�P���+D�3XZ� Ȉ��MVq��8��,���|�t�ç.���ߗn��e9�Y�df{="��$��Z���:��� nK�;��E6v*����1���� Қs�m�+�9=�b;��h-�4v�?ho��~䅀�
�O�o�'_	�Tq/J�����J�V���g��6*䔄�[�-��O�OC|<Ć�jAk�;�P������ŵ,?����*�K��˛�g�V�zy�41 ]-��y�zBv�tJ�܆��ec�C8�j~�i��\��1�����E*ܲ��bfT� c���LHY�&�[ ��vS|L�o��<b��&sӞ�V���՚h������Ж�+�>�SJ��wp�$����G�ͺC3�ι�W��$�}��m2�p�@��p�8���R&gbՀ�n�h�a�Wg1�6tD�f&6g6D)>����G�s��A6��`���Ё����飪�x~�P����R��IhH�GpNQ7�q�y����V80mz"�D( l���a���M��T��wlf$����^�����pxô��8�Mf�N�{)��N) фlF���������AГSN<ӟx�	̬�W4�j;�W����_�\�G5����$�ϴ+����yP�߾q<�4hOSYl�C"[*8��j�V��%$s���U�1�hutY[:�ޱ٫��VK9�4���m
���3��Zj��y,[��.`D��:mG�ZD����*oE�i��m�������	�#�&e
�Xfis77A�2�d+r�eU�ul]�GKџ�׷�)��-f�M2L�I�ɏx"2�
Ӡ#Q��$aA���v�b;VAu��z�CdB[����a�R�8��U����������2�#�~�:��{��r/�����J��r�ٍ�������:�-j4;0���E���%��l���c2(�J@p��B;t������j}���>/���-�\�Sp�\N%������1-xR�sG���Nt򸽒
e[�uz1�����]!�QL����'d?��3?>\��U�@#Z-F{�98*���=�݊�þ���~x�O��L)�����*��ͽ6�b2K񒢹
�3B:�_Xl���C3TX'����q#�E/�y���9�Z@%!G,n��sTq��"����5��P�?���� ��vԤ?��i�]���vz�F[�/ch�R��^<�� ]������|���x͍b0nhE��:�}��չ��HB�O�ͼ2r�ߛ�Э���<O���O9]C�,������7�ڮ4���堵�j<���Ub4J�lJ�T�
خ[�73�q����T�D1v���mnH�����k%3@�_+3�f�)ĥM�s]��lIwQbVJU��ZC�xO]��
@	�Xz��I�@8������ I*<+�� ��ѿ�`�A���Pʳ)��MɎ
 ��h��"v�y�;�;~A�m�D�9ˉx��Z4W�,/"5 t�癮�F�lGa���vyj���;�'�)\ϔ��!�[y^;(������t#Q$�h�a��I:"0杽E79��͓��=������o`�5tNQ�}K2��-/I-��>NR�d���?�"���,/eù�i�oz�G̫2/�]�w	Y��`��?��}�I�s��� ��_ǻ��{�hD
�<TQ�ήi_\�	&���بㆣ�xJK�9	�_��Q
���D[��k����mU'9ߔ��� �B��"�Y9��?L��6���.��/z���Y����`�܏�p��mӟ�3�H�<&z�B9_�P�B�&���-��꺲����1�1�!�F���Z�1%aHpDOz���t'
�$�����^4���so#����x�3��ˋ�dCԙ<��a�/Tm��ZHm6��;�7�P�(
�j5�?�^�c�6	�{�����-p�Zԥ��f�9�s��}GT���&����#�F+1��w0R���h��<<%�-�E��S2�4c�=�*R�2#��9ȝl���̩شW�8d�T��0�-_�b~O�6�Yn�恄{G}b�d�"T�>��.i�ݪ�^eH�q�G�E��mPɍʴ�l=����aڛ4��C>�5�|�X�#�����U���imф8�!c����D�irB��qx�f	ߚ8-恋��1�c��q|��|0�yjX�,�GR�L��Ɛ����U��p
��84��G��2�v����:7,:��4�vwb>٘��p�d��KR��ʪs����]��|�}�ڔ����llk�s���(��8��� ՠvK?}��j���a��F�
D��+��
݁;H�cE*�d�[+�����4Qg��K��r�ӫ��A�M�P��>����X-�m�0j����*1�}r��ص�|�:�ΰw%���yA���>�4�S�ƺf���� x6{��UڲWM(�Vz$F�!�[�\������U��&[���xy��<��������#h�x���Y3ܮz���`VL�����O+c��"�Sgqp�����#�<��_FüU��oMY,�Wî��备�'{���_���f0E�4Վ}�囶�4j2$J��7}��UI�@�i��!E&o�ⅻ���n�)�I�r��M�b���%zhu&��F��[�$������'ܢ]-��R&Қ5K�C�j����钛������6�X[��>����lK�W#���uZ�i���γ�1��^`Pҧ���̚��z�&7��&��C�I?��UD�fjݬ�Uԁ��N���H��;�]�T�5�F� W�5^�q~���X�ަ�H"�Bӕo����~�鈉�S�X`"�p�3�輊�cp�a,�b�R\�{a�jW�)ۈA�O4��/ Ø���Sk�0�r�J���Q��dv����\W�V�Wki��'��l�E��sc�｟�8�・,�������D�ȴ�<�4��`�,o�9EV����L����	Te�`�I��,�Ȋ�.�l���d���'�w#���k�Z��P��؃Mgr,�zW�����A\XK���T����n@��C�ҋ0�:m�z�V�FE�X\�T����o�I(p0w�w*FY=���_��ޓ"�l�-��zw���k�]�r���7%Q��o�#��@��a]T��z����է0#o�14[�6�Pޔ�IjL�͈_z��jgp�/�8��sNˤ��}�%���������X�']��C��2�yV�FU�c�is�H�����(�3�e�l�A5�φ_\l�q& �>�C~��_���F9���[��8)�2��㩇���J0fY����ŞVޮ�L|�����L�9�]����{��)�.�щ0����(!ŦCH��Fl�6(����^�f+��g�<��Ɉ1C���)���V֨��:�
��Q�O"h�j:� �ш��-�����ي]�c��:L��
�����"��fow��s���X�ý=l�>Q��B�qC�S���Q�S�]`���,b�<	����U�M�r�؜[��E��e�����r�ݯ��V���lHP~��}��C���>S��K�����L���1$�(��(��ϸ�!�|�P��0M���5�'A�y6� u\;f���s�å��ݘ�Wo�p�$�?�'�?����"�徐-� �C gNQ���9��^�X�g�2x�Ҽl���+�T9�X8k�0M�
��j�{���T������.{�Ҩ<�S��h	\���YEw�R`��tj��5��Ę�D��O�X[VO���sg���W�>PH;r�Yh��G�H��zWrn�oaY� |��a��J�אՅ�����d����n4k-�ߨ8�2����Birb<���Ƹ��+�8{�R�S%�B}S�q��w��D�2��j���rGrE�2j����.��V>�#�/?�`	�j�RBh7�t-m���A�!��:t�q;RU�]� �9
��&׶�����䰢���f'}�����+$���D�p��jJ����;��{�;�=�Yi�ȥ��@=Գs���}}tⶔ�)��pX����Pt�&��y&�Xp��߷�@��k�x
$�P�_���-�n���Z�O�/���+q�� ���|�b%[�X�Sn�{>�-�Kg�3�`w)���Yڲu]�­�� �w�4	����0�p!1�5*��Jf�,GjO,h�J��
��\o��������n5�l\�fB���o��8%2�:`+���ռ�g�r���,������Lv݅� ���홇oY7�M����x '��������E� @~$O�4��~��R��J<�)�~N�&���\�`Ba��:&tQ���j(=`���6�}�J�ov0�����^��2��kD�qX\4k���~���u�&���OLl�&�+���>�M��7�IL6�1��5h�$�yc#1����=N:�N�@����l�=?��-M��t�����XH�uE[#�g�Ϲ$�ŰፕO�a��;x4t��ؠ}K���ZE%7/���u |)!M�����