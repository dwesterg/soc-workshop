��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�_�L�=�g������x����RI_�������=t����z�2w��.-wx8N���(��ZI9:\UC1���(4�k,���$
�`[x�B��*�jo�KZ+�pĀ3v<\ڵfu��5&v
%��
��� ��^"8��6?��OV�l��fv{Ĺ�	O�8���j�/ř��WXkK+�kf7�Z;p�C	x>��	&Y��.�e�5D .��䓃��wW�-�AP��P��Q�N�	�b���TȀ)��(�h!����#˵+lG�=_��.+�ա�]k1�N �x u�!��rZ��P��ΰ�tl���.w���\���[�ɡ+	���|bU�_N=�w�CG���b=���H"�O"������(z��H�*$����_�k_�0���/�`�. t�ﶇ�>��0�unvE�����y&.�0��Q�e��\6#M
dj�h~����dL�a]�:�'gPk��<��9	PM���k|x�qZ@���W�V��EM�u5�MC�y�o��`'�Ж���8A�K�+�s�
p�͂�*�����Cy���<�*�3�Y��)��j�唓�5C;;�cG᫓�kڗ/P�P[��dtb��[A��q�X�]�0���(�:�(C��yB���4�+�2S���ʶK�~���2u>����~I&R	`ɐ��u(,C���7h}���q�cD�E,=�q*������8�T��D?�eD�&���M�.���T�j���>6�WUN���t	�nZZ�S�٥�`x߱N�����/#ܷ̅P����⊢�/Ȝ�ڝ>�4��E���7���#W�'&�yI��Ҫi�Q�25��;Z������ۄY�P 	yc`A���;�~�g:��;D����V�Y({��6��c��=��W��Q�	�R�������}�G_��NH��������axi��n.iȎP�/�\}޶���r�����'-�+޺����/�d>u"(;B�x�=�	����M� �"@�f���	x�U�
���l�v$y�e�L�:K�W=WC���p=�ɛe�iw�hvޮ����4O��f�$�)%>���x��C"ɝ��ᄡ^�䖁���b.ĸ�ƙyw�0�[ؙ �c����S��9���n%t3�E�W��7KM�<�s5��x;$Y��ޘ��3�HS)���I�D�lCG��xĉ`��@��'���Bh�Zى��-���
�[qw���������q���������o��m����s�a��7���h���s������z�q}�zYpk�������xu#��D"��atd��D3XwrM���0�/}	A�Z�hG�/��e� th�s�{�S^ƛ�buM	�����o�O���W6���|<�~�ԟJ̓ӓE�-�"9�_�y^�����B
��~��`Һ��>k�57�Krd.�B<��^�������!���Qo��ת�أ������C_��T~"����u�eu^�R��4���҅(=�b��C�A�?��sY��cyS���ZV�����Y�Wm��lx���,T{Y���r�sz.��(�D#ԓj<����<��w�r�_�0��V?7hS�ft�e�'���u����d���ǃNu�IE%<N�zb�{�ق���w�E_E���A�kS$�rjQ�r�1����� }�/J�����%��I�[`bŔ�;�U��h�I 3˧=�p�����և�u�sM�]�Jr�\e6L�a�@�u�<���h	�mK�o�\�}��o��P��
���X���H|G��y@� �p0�
��v0Q_*�5SC~��S<�w��ѭIPM�A9C���[1t.�-���.�ql����7R��J��_���h�՚ �f,�|�Jx�Y�d`�ZUyF)o&�c%�5Y"w-uߵ�V�X�,�d@��=`�aO���
zpH�חbkJ�# t��ձ���o���]�;�UK;S��T�u���^�"�lМK��HmqySOĥL�bЭ�uu#4�ٕAr�c=6g�+Z)0�q��c�4�֜��,� }��~���ݿZ�o��-����Ka)f=��O�؂e��/.��tn�+����C�@-<ś���;�7}S�5NwO\L��^E�=�0{��A�5j]�AUH|����[f��t8��\��o�J��0�u.e�p��-��^�	�񹟭�U��zw�h���B1�ݼ2���}m@�a��^ui�3�Do��J�n�z��ȇ9�(.c!��g_ʒ��֤_���1����{oV�a�>��R�9�u>M�n��ݻ�Qڴ���X�lOy?	���ً.NS��O,����Rk��e�g���l^�K�y0��ݼHR��^���*�XbL+�&Q��{TcL NS�����Thu��{=�s4����X�IH�yS�ϗ8��X�RX"s�K��2R��_K�+�f��e��=]���6{��
�ߴ6�g_p�,�W�Ct����䅼=`��[V$8�!�(�eO��L1AΝ�
��g�L�>�K@��@��ky�Ϡ��'\�����1?B��m����Ns��J��a'#{{/^_���8nVNH�d��!	Y,j���� �1 _u֏�E]�6�n�l,"�Z<t*���2�b
�����%=�����k�׮�H�䁚_���M�:x�B�Τ��ʫ�����<��w�5��	W��R������j��h��ItݍkuZuX�q�����+Sā�M<�8q����Z~mS%l������!�ĶrQ��Q�ƥ`&�[�ɜ�橾�TJ��in*E��D��@�H�����χQ��ʭ�~'�E�^6=����g�����4^��O��6��*D����^c�_
�d���ǉ�JP�����QE\�mhf�9ŧAM�;f�)b��sm�ի*5�0�UI!&�5u[�Q ��d7��]�J�k�vU`Q5T��� n7����{��,?�7�)�����#�qX��	;eG5eLb��_���et�O�n��y<���:K`��;f(�hJ�=����.� �&nں��'i�����L�m����'�|�i߫|���8�V��ѦG��V�콞�Ҷ������H8�$�BZǹtb�{/�k-$�+}�e������ob:��(��d]�`�;�/J�JA�}�v��j[c�n��b���(1�cd$P
��@�rޤ[�i��Ֆ�����<���b6��H��PQq0.mZN��pSC����٤"�w��@�,��N��o�	��Y�E�����~�'(�E�X����b���F�C8�d�[tJ	ؑ��mR�y�ϵ�/��-E���7����H�
�"���@�)���[���zz�-7�R
<�p �H���_�e�d5�qF��=_W�O��lc��ΡAf�!�jjG�`�ٳB�x2�	��?WT%W?��x:�,+5 +|���V���Z\��׍\�t]s��}��GA!�2Y�但����+^&iج�>;���~�E�M�z��s"}W&�S������^��W�FL�9�����#���+G�����~O���#l����&5*\L�d~�0�BL��W��}~q����f��:�p����!v�L"tT�L����p��|��d��\J�ŵ9�ɏN�:�p��2���[��I�i�����1�ꗡ�ha�����W�jn1>�`�]��l�~E%(Y\�;w�dڢ�I/������'B�_�%��_``����Gҗ�?;9[�{R�X���j����]�a��!�b��f��_��,����ļ���b3�v��]Q�̃;R�2�ֽhCѯ�7(�|s��͖�y:j\<�fCl\��3+":&G��-�Z5{����Z�z��Q|O_�n���	ǩ�	W��RYZ�~.�D�QlD�7�[�{�����ǜ]�M?\ڬ����oKK^C��ٝ�בb��qۣB����m������X;H.
����I��mb!�h���"=����B��p	@g�+
���0�U�E�{O��ʣ�>���|(�;k��
�מ�	r��Z�Sw��(Y$�V��5���3�����ޟ�eF+��{�|Q@�Y�·�p��ZY7�onr�x�bs�|�r�]��Mϼ��%�,��ǥ����OHA��na�'z�6�j qD
m��Th�����#2&ۿ�ZjqBD�í���E���}�d��8l$[��$�>@�����W�-кaw�x��dp3��FVb�,�K�o���u/y�D���	RM�T4�4K�\Vj�~���|�4=q���T>;_��q1o1�#��5�ў�(qzdɘ�����/�
�+�F��F;���lN�����!��2����3�Vday��̆�h�	F����`-�eq�����Qk!'���>�W���8�&T�j�bjC�V=m��1�X���	+��&ȁ��,��/�3' ݿ�($>�]�_x�*$.���1�z{[K�Զ�s��ON�gכ��}����+��xI���a����g��o�Rb�1&Da7�N�����xI��
���j�2n���1��d_�B��0(�Zhw�H��o~>�X������,�Z*�9�^~�Q��ӌ�����{f����&�< 56��ӃQA{}����[�F����'�'���o�j�A �*�v�A��IF���>��[���r�*9S�]��оU��է�?� {n{�%VGD�'�`$n�nN�v�%���(�sF����|}_6��W��|�����+Ơ��L=O�
CL9r����&?��f��F���2>B���h�x�GX�asiϮ�h��di�2m�|l��b龑l��k�A������Cїߔ�n������E$�1��~f�����W(������X��h���Ѩ���u�����1,y��8��h?ƞN���l�?g�/��� mQ��f#�o^x�)Z������ٓy��r�j��q��dQ3z�5|D1���D�ÌZB4V�.�}+��9��~�_�L�lX!�̻���p��r;���y�;m!�ɛc$�K/�|���|x���w�9ʯ�0b�DQϦ��|�wb���A`�� � i��+5Q��\α2�jxi�S&bUԴ��%�s�4�BǮm�}���Rd�&�S�5�8:�o�{�ɼv���NU9]6�q��cgc�~=��]ɧ�ԝ��9��g���ƾИ�8P����PGa�����^o ���̾3z�5*N�D���uDh2*�aJ�`��i���ku��PeL��J�ǜ�m�#��w�b�:G����n9.��8*���uQ�忦� �ȆN �],Փ��OϑHUh~^Ww�Ƞ^�<X,cGk,� ��[��8���XJ>B8��!	��*�Z����Ҋ��r4�U�u���VL��g��|ޣ����QZ�9А�Zg�Q��7>b��"[5y~�OeK�C�pђ��
<�b�g��u�_j�+1���<�+XagЇĘ�d�m�Er󫩤u�w�Ah͈�K������W��v��	���8�A������F��x\��1Ga�ɒ9���į x�L�R��G#�$SM(Zz���"P�3�\���.Ž�$��t7,�����ֿE2����T[k����Nq�P��ت@���n,�$�/�(׹s�;��ZKDĔr�ZĬqſ�lc��OTU��?���{~��'�����uI��W�{wPy�F:C��'�]�ALه��l�V�m��������&�Ԛ-"��xD��z���B�� ��y���=�H�F�7>�GI�$m��G�����6��c��وI��Lm�_�#W��jY��}Տb�J ��h Z]�c��j��㽲��
K'��\��Ou-��~e�Z@L����#�p"�sX��ݝɹ1�{ȕ�>����\₨.�f���X򉳠�(j�'���
���G��A�%�E����A��#���"Ub���Z�1��҂G�d=��l5!ޚ�4�~�`;�?�e�/�)���je:��3�Εy>�j��x�mU�:Ƥ�,�;�^�鏉�0�2��D]�[��L�~FULݒw���4�N�/�o��o2M�	�:N
t����ff�����1㋐Mڐ�3�W�x�u�"'�����ɭ��}�FS��b�i4�ppr �j�A���"�c�)gU��$�]����9E��\q���|��ױ�q��Ǆ8�x�2?���6�J��L���5�;�[U-%d�.8���Ɖ�����w�h�`gW��Z	���G+H��I�x����I=�V�a�ӥB�A����}�w3rXI��wغl<]#a-A�ݩ0�O��,��%=����9R
���<��y%�c���p@f��h���j��:��3�O����k"�Q��̋�x&����x3��:����Ld�o�K�<����Qe��z�:����T��_^;D�8�w��.;��.3-D��q{?m�u1�����S�7[������J�n��nM+�.�Y$��1�H"����H3�#ݚ>p��e�-�3sRs,e��d��s�1W�ĕnb�(̨muB`��q���dJ�F�1WgW#Lo�S5%f��Ou�g�D\��\ؠ�!���D@5�nawW�7���H&���V���,�#'P��j�TSlH��vf�<�$��Q��,|{�B@i�[�P~���z�V�"�(��Fk�������	��Lf�� " 	֫㒳"z�oK�G�Ej,5�,�N�֏Q�U�Bv�u(�����H���"3���4���!�ߟJ�!9��h������^|��W@i���@v�ڰvq��g�h�Q��`�
����S��Uޯ?�FY3�A��J�)�L[:k`\HG�u|�z�a))�se?���w�LRq�쀩i��8�B��[���39�g��6.��:�5���`Φ�?��S���`�/h�����B�N5 Y���C�
4WQġ:+S+��O��G��e�9v��ëv��p��Ja�L-�P��ehwn��$� ����� V��Af�)j)H@J��EG���(�)tn��K�F��
�����e
����"������1:'�0��\��G&������7����H��y�c�͸���<���:Vc۝�#���d�U�V���B��]E��]����}���>qI��3_���`�2}���Q�RY�mP5�l(��X5n