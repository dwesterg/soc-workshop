��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+?�9��"qzC���0��tb�%m�o7�(Ɏ�u�l������`ڴgQ
w"%M|I�ۀ3c�m��r�����&f���v����f�%��i9>�*��6�-��k�IZ���Mڵ�a�a�xfH� =�A�oR��ɼ�	"��
��(&-ͳ��֬Wfm�_�+�Y�rPy�2Q��2���V��y�����^�^�@��=��,"�W�����7�݅�̧�E���؏���_ū̳�)l�ȗ
�,��V�н�C�7ג�(�W�T�YFc�l0�΢�7�&v_����!���2���$b�k��?'(@SI�QrQE$^'A�Y��yic}f��!�eyB�J���@�W��P�O�XX�D��++�Z��B��4�!�W\�;��.����r!_��9G��@����ބ�X�<ꮪ/.���.��H�D>j����V��*�;��h[y>�_(��!1ݎ~v�ZjWm?�G[����F�m�A� 5�);gȑ������d�Q�9�ھb;7A��d��a?���	���L7[�����
��0��!�Pm��N5Y*��y��+�t���0T.���I���a�g�c���I*�1t�g���B�z%uՈ��8ؗ�ca�	�co�ݒhZp��I$& ��<;EL[���Fu��9_>��GW<r�LYK�!ػ^[���P�<�*��lC(���X[��P��_�`�� �-�W6��ٖ��5�
ѿ�Ԯ��l�Prc���{6�|���Y/"r��@�	���}��M�)�4�Pxv�C蹉!��p*��-,�� �*����=GW k?�āY���4����5�7%�����	�*��VA�g{�,r/L~�U,=Z6�4�bv� 7�z7���W7���"����䖚%س+�}f���C*�v&�l�Cp���+����̌)ֻ=��5�S�H����`����� |0T~{���$��Ѯ� ���\�ٟ[���ḐX.X٧ⶎ�2cyv$@�|�,�@$�[���B"�7O����Z��Q���[k�k�.��o�Cء���w�<�����ָ.�(Bh���)��A߂�f:t�Y�Bs����,��Nd�`�׀Ja:�C$\��,P���?���ovK�������)���`��"%��,���b��%;�zh�g�$\
b&!�0�ܻ�����e��@?��t�*M,?]H/I��ppk�c�o���(2:�������^*tToȟ�Т5��@����،�>kd78��>�6u��3��NHU�����z ��~D�z�Z� �-��&��~+�#�� kq�?����`��깕/T��q��0%��N{㶷�|jP�Yc`e�T�!j� ��_߼:��$w�Hmj�D��L�M��o��*���m|]As���{y��|P�5wߟ�鎎z����p�_�5ϩ`�p��f��{�kia.5�_�,�8F�Q��"�|��~��3 �����!�F�ڇ�B$�4W(�y��G^��@��4bN�R�	K�￼ڇlDCn^
��b(9�q��F��@1�US�r�4����B���o��W^H'�i��������]Ś0e��i�\�E����,��0o�.���������w�Vq`pZc}�yJ�\��;�M�`����v�$^�7i�yTO�%l�"����8��R&>�����?+��L�|�����Z�3��h��˲�����3@C������C��w��l�B' ,y��S�C�5$d���önK������Vm���LH7N�+�"��̾ԩ{�299w��j�آb/0�Ű��^.��b���j�w}3����Uj]�E���-��ENa�HtVq�<o�?�^��k�)�i��I�Hw�2�җ��QY����7�q�(z�xm�L��F�_��P�Z�Hu��t��c�����UH^�Iھ��m�����j�p��H� `�u��Xrl;�e������5���ADs�J�+����$\v�� إ��탠߱v}ϻMM<~\�É� �tF�!��C;����F�����)�X���7�T*#�'��kZ�ݻ~D���%���O�C��N>ϴ�s�7����F�_ɥ�7��%�8W����-�7� '��&#s�Q�2ۀ;c[H�q�Q`8o@>V