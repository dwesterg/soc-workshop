��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bdc��NAs|%�;JN��}Oݮ�L��-��Pɾ��2���O=�lǁ����Jw��ʹ���c�����j�)T;k�F�XHp?<K��Ǡ�����4�� s�3MT���<D��{����Ֆ)�$�)H����`�a:�b��c,��Ud�S��+��`g(��2����dA%������B�nV4J��_|��)%�7f���-����|Y�G�5��am�>,Y����.XXKݾ^�_}L���e+m�x�`�j�Z0ww�p��0��e�xY#���<��h�n���fti��zWs#B3'; �d��1��N���,�Mb�E�ů|�|��R�u��c�"bB&�N�vB���H��I3~F��q�qX�D �4��4��R�(@ 5��r-q���3�8P7�+�"��xm����|��ߚ(�[m#�19I�?a�?Ky�2~��]��������\ �	�|.T�1��F��<L��Q�������?6~r Qyaɮ�4&�ڰA��%��DY����\�k;:�!G֑�d�
�:R�˓�W��o@7��\� �y:��!���O7��qkP�q�sbǜM
�\�H�2Z)Q��4��Ğ�0h�p-m����[���>4{��mP٘j��61:%�tx��Fyᢞ��C��2�
8��Zm���Pft"I�,�X{U�ɡhq[�P����2��+���������"�����f̈́��QC~`�
�;�!X�z͗��lŭ��~Q�W|$���-Z���x~GKp���Ǉx�z��%t}ɮ/�!#��������@�좞e�(��v<*"J��tm��V �DG*����4�?�J�YZ�R�k^�]B��WX<E���5�h)�!�z�N�J
�\����S7�Mv���6���F_x�(T�k���}A��7�3�����1�39ر�E������ r*�]z�E\�Lw4�7k��(rcʉH�g�L���iWYl���\�~w-�\h^�t�W*�g�P���>��KB�&�^UۈAd�����SjCޕ4�0�M!n���'�阐��҇_�T�.����Z-�F��#��o7}�i�<�-L;����xn�����ŉ�"��t���/x��_�i&�{!�CNe�Ҿp6���C�D�	�kF�buw}����vGH�no!�㛴�ԹT�Kn	�̉)��U|�$1��7̋>�U�߆��A?�K�HZ�>hM�qS�;!3D�*��}�%!c�^κ�.�*Y��^�0y��q2/��n�2��YBmu�)���w�+�N����|�lW��5�2�@�r0�\�kb��^����ܘ�J�m�7����ó]B��2�b��g����@3�=T7���㩣��O9���]3�� 8���Զ�(����t����c={�vK��i�����ph.��( ��[�������z�;�N����!�e�l�5���_��QG�}n���&8Q7Az+�M������#�{�{:�y���,h5D��I����D#��"A q�`/	�f��֎�r(�]�>�������������_6B��0�&��AD��f�,���Gkc42%����	���O�sU5g\�׽�.�r�s�J�!��¼*�v���x�8��qq�1�����c���{�t̻�!��UI�����,?�ygFH��:������e�\���:tV��9@Fj���	2	��+��R��}�1�I�?����\�f揅7�3�,1fI\㝄�^^���)�2#g�'�6!��?�8�
���{ǙӭR3G�gK6w ��������O��+�XQ�����;-{�p�6���h�%.��Kw����t�S�91x�L·<�{�F�;�Klv���y�^�y�t��VQ�2��Y�����	���_���K��i>(XT�PvT�q�e͊��mӏ���a0H��B\~��{ceT��_�n�*��cE�k��!>�2 X9�ʯ4�^v�![�䟯;lJ�$�L��0w0| ��U�y�Tm@Y����8.�T�u�7��R�.-�)�3?��@���{_�2�s���\ >ɭ'N��n�KC�x�"?��fDӨ-�?BO�(�H?v}�.�`MlY��|�zNUU��((�W<!�E]gP��b�돇AR/26��_��M���(p\p��61l�ԃ	���\��,[�� �Yu�)"������k  ���a������ny�L���z��b3����g��H-R�+^��Q@|����۰H�'�����U�{�e���o ��F��y����1�����V�ý�-CB߮mC�1��ƿb���EI9}YI`��!A �hi�;�N�&}w�6Lx�4���a�^]�8��
p���m����F���Ǖ��Qch��)F�|K�s�+�	?@�8�Y.	��iN�.@8c�yL�T�j*`�sq�y�EU�g�w�nM�Mx{�e^���5I��׀��YA��"8R��c뇘"�x�Ff1[���F�@`D�; �x��,x���ߤ�[��pB2�o� kǃ�5�Ў����b6�%X��G͡n����8�F����Ħ�V$�/�ڇ,eP���lmu$ؘ0�9���'�v�@K]��K��x�������lQ�����qE2���+F�v��嶽v����M�����KG�������|��
�?hʠ����ˬ;cF�	7nՍܬ�R,�IT�/~}��8�I>���鄀2��< �U����W!d���X�՟ޱ2�y$߶B��V���OŊB���)��f:���#�'�2UQ��	��a��w�<@�V+Nλ�Vm��$鱈F���q��	�1���ګ�L5��l��9�O
l�NlM�(�`�HC��q��ʃ׶�b��9z��R���+���EEw	�tq�����5�@��7�=�4*��!֞8i)6�(pbٰ��C!Z�C�0��Mz��YjRq�h���bdЏB��b�聏�h��M����|@��K�7C"�B���xޮ�����K����h.�	(�5�@����1�X#�EQ:�lh'�^���	~�F~��xZ�!��Y�-J3�v��ǰ�k^����ع�~�H�;�X#���o��t� +�\A%�0���UK���Q�gQ���h%��1�G��Д)���nM��1��\�"�˳ ?��xdW>F����	�1`���3',�����Y࿫�h`�p!���t1�41S-Fs��cR���l�´��*Kn�\H ����9uڬFJ����Bl_�XQP�"��;�'~���8�%ڰ�ʚ����Ȉ�tΠ
�M��u#�����}tH�<e�&.�{a�{�C X�b<_��9��w���Ъ�s�M�_�N�]�����%W��#}�� qI��ig��+.$�?
50���h��־�� ƭ	A��\�fŬ)���@�1�|���9!�n�
�B#�	C?�&K;�5e'i��ȶ�����z�P��`k��տ~K��sԘ���Y��F0�-��5b�<?@����f���|8�T��;�:�o�_�e�3��>P���F��6�S[����qT�l`�Ϟ��*�f�>��Cp��� W�S<� [u��b������͵�L@��0H�,��ٲ��j�,Ф҆z�gn�u�~��Ou+;	'�~EI|��C��VΤ���b�|�%�}�� <Ɠ�uU��:���s�:���+�l�W]O�د���>�b&	hnV7�\:�&�[ڇ
wf�a磞�}y�C2�MO�&iO~=���;��/�A&%���2,�Y\g����ެ�l ��KN�H�V6J_�?i�#"n��aAt�Mv�8T7���R��g&[��̞m`�݊��ǭ���z:j��]�)?�����Oxc���i�E쥐<�% /|��e���F��D����Ýڭz {���sp�8!����΢�T�DC��g�  V�q�k�9�*+�b�ސ�*�["�\3�@���4�nll{��/�􅺉���L-���g�4�[�^0�|����-c�a�њ�p=.�H��]�����c��ѳ��NtE<,pJ@�R#M�^����,c�v�g_���Z�d��?Q�r��c}`�����U:��8O�;����	�x��B��c��>$ّ9��DB �\r+����й�C�|�
Jm�]xЂ���h�!<ҡ�RőB���i�'���Oa���	Fb�������Ṹ�p��<��c���؜V:��E][�=Ĥ,4�7�E8�{�p��ƾ�ט�fg��"�P�����|�##"��O3�;�`�U���u�u�F��'��^�pJ����	:t�+��p�z"�o��8=�jT��S��1�$����#n&W�d��g�[k����� Ϭ|3��S�i��/읪��B����P��^N�w%��6q\E	ϼ�����FҠ�D�X6�6�JT�%[*�! �y�D?JD)�EZ'B��l���Z�ȾuC%�"�Cm�AI�&a�TF5xx�T�~D44��ؔ�~̠�t���G��L+F��DnQh̀�zrc�E@���Ž���D6�D�t߭(��/�4?#+�Mp`��F��9`��)9u�x�(RE���������E%Q.O�
�\�XX���,V/L��1�4k�N�ئ�(%
j��{�T�B��ή�쏨#��\�N5��������--{R6�b� Q���g��׵5�I������'p����N�%��7��w5��0�%��N�S����XԽy
V�	^�8�B����k4spF~r�[�6�&H�G�vs��&h��G�`�/��tC�^��GrE��Z�%���o	�_G��ջl��:����0e������R*�J�;�^r�3Y�F��9N�8_O�:	 a3L�
�p�x+Y�o9��2ň@�?�4@�*/� ��_�
�kGmA]w���t�b��5�Ȍ�|�[Y�	z:�Yx)���RR�b	H|C����a�):�,Y�e�#�M���#`yp�z��|��mrYq��֒(!����	ʨ�3UY���w�tSE�@��1���K+�M����:v��Ϙ\ű�M���� F�	�(KG��h�G�0��XO�خ�8�F�ĢD7���S~�8�T�Җ漎�)Y�~��0\����T�(�䅜&�-�]U�\��s�.����D�\�z��1'�=$xVT��Щ'&,*X��������v�pTz9��m��NZ�P��r&����M)��p�t��H,�"��/9��{U���Unj�'��˧�G��$V��y�ش a~�#_��#ݛ}����-�g�p���0m9�ƥ��[We�a.����n�N�~���,�е�
��;�'$��b�M��ua7�|%����.�wK�0G�S��"MIŤ�ڃyj˼�����GPuhP��k{z1O�/W���@�&���Pk!�ޔϳ�G՗3J�7`0�v*�	�+�>�S"��6����5�)JqE:J�;�id��<�<�#Wv7��y����
�����Xt�J#�;�Vܢh�
S���KD����/
h*g��N��WWE$/_wR�K�ݟ��h:Z�4h�Y�Q���l*/��ő{h�;55���;�U�y�;QB#���t�4q������(U�.����I]7�vZ��`��P!�a��霁�2ZTK o:|�����Fi�5���\�%��$A%��Q�D�dӃ�1�t�=�sD�'��6`5jq�|�E���E�!w�5T�����υ������)QC �M*�?���g{�]��ݬPh>[xq���x*��I�ƙixn\��n�����h������ed�-q"@ux���?J>rʫ���h���"���\�?`XC����\wM���.+�t�e+�b2+�J#���z����L\�|!�0��R�̝���m:��!p�y�V�~�K��Y�b���_�e��cZW�m�7����_�w��#�J��X삉�j/Ĕ\)y:a��t���x��������kE�ab�>�