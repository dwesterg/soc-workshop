��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���2_it��S�����qR	���f>wd��4���&V�*�b�_¡rc%�׉�m:�G�[����5Jd$5�&�t�O�,��yp���i�j�W�y��{���Oԕ-8_�7TՇ}!S���V��,��kej�)|�L�{I�Zo�8J|��e��,'^EoKEז�O�9�K~vK��M�5/ʩ� *���*Ǒ�ة���i<eR��nM���Qjv�k`�4�#����o[#��PF��n�寧G��G4��P	��~�\��:��R8�~j&r��=߾~ tR�9�G�)�~�~�#CS����g�^4���I(����\0m��3	"hw�n!t�;��6g2�)`BT<�ݴ'��;�O�6®���lٲ�/#�
9��l�cov�v7g��P�H��&��\X���Y"��`�f�����j�f���a�2?�(���ަ�<��98�w�X����+��%�6� c7(Zˎ�DfE;�g"�qo�9�����I4�g�f�+T�!_Ƣk����F�dӴH8U�pJgr{3��M#E���8Xˌ=������.�`�O�`C�4�SS���^�:F	����/�=�:�8y�7��RҘ-lt��N"��f$�l�������I*0�|2tAݿk����w@��L̊cI�̈Ykj+�l�	��<%�<�r�iİ�L?�qxSy�LÃ�x��L*[��d�28�x=����s{5T�<�GK�P���|���ˋ 4襏W�M��n�d�d@oDL���@���n�K���(6�]1mb�<��u�2�l�mB�-�-Ў��ċ��<�D��.��_p��9�~L��J~��|7h�Ø�,ۂ�t*<񣈞8���&  �]s7I�*�LU4ؖ�$���v��?�R5fP
@?��7���m�x��#�vQ_i{
WU�ٿt7~���9��>������6r�\��@6(�K�򿒁Y5��Ȧ4~I��CdAQfW1�g�'������Q���y�҃�˕؛Z�q!%�����[�^S�ы�������è��e)��������(bG$�yכ�)�}kݳ��$BX�q���&��L��(���E˙R2;i�!�اB̥I��/�Ӝ�&��.8+/�C�rQ�:b]��lS�B��=��	5p�^Ե�N}��L`�ĝ2!)q�o�0�K���>s<�� ����"�puM舑��z�f��� ��<RG"s��W�j����j��.`o��̣ũ���)U�����8�I)�}��w��0@�9�}[�|Cl\�mǹ+�[����@T����t��-�mn�n����:s��� ���n�b��N����Sgx��ã$:�=0�f-�vj���=N?�=����	�e��e
(x:d�G�B���r�v_<1vs�B��'ߺ��tq�����q������ւc�̕ST5���]:¸Ү���.:-u�eI�
��X ]f���=硂��6~Hd2D������6gp2ZUz!��U�ak����d(� �:Gy�p����g��2�� 5!Puǁ�t0�{6�Xn��g�G�K��W��Hc�5��'�b�Qs������V.)H��5���O�0��5���{��:�ziB�Bb�gˊ�j�Q��|��6��� ����{݀�����ko�F�$�DrYm�${Q����ɕ��Q���F h����%*���:��vo�di��8�!���;����o�C�W|-XWZW	�<?�e7�%3�K|�����������f�A���&�jT�w�BX�-����iMf�>�U
�(��=�"�����=�T�+Q�M�g
��P�H��o��R-r�ʅ]"	������2A��@�G�v�����=.mi�s?���Kgf�����c�,�+�����m�z�Ӊ�q���v��>�4��Ii.��QY�ӽk�����u�� ��(qRyb�s���En��� (�Dt�a]j3��V��~J��&ȲO�H/��;� �mAUQ�N�����]��F�{�j����	��7�f;��@��*�,��F�nսM�.X���j���[���U�q�C����Ċ������~X��9��5B���(#�y�5!�En��I��,F���Y>�k[O�b�{c �8���W_��0��R��ޒ��¬���ZR��O˘X����InUe���V���#��m�fK2�ᐶ��fq�셦7gl�|FC��v�ߑ���:`d5�yBu�ri��^�i2�H�t90	5�v��#Q�}׬^�r��f�l3��q����՛Q͛�m�Dv����g0iV�4��>��+N�<j.Z��LC��n@R���L�Ν|���q$��䪛��CXAK=_�Y�������q����$�,���H�Pbg�d��16�B���!G�8����v�a<n������ 4�KaMK��u�dv�.%Dd;���x�X�>������h�Mt�%��%�ا��.��:p�$��U�� ��S�)�9]�z|d >��,��e���vȩy�h�U��T"��䏛̀dX�iГWq��nF�fqѬk]#R30���5u�NnŅe��>E��D�{���l\vLj��7cA�����Tq�[�_� �/T�@�p�	�<)���?����>��f�k�7�����霘����ʘԨƄ_���Lp27Gx9v��J��X�pp�.3�S�=�n�7؛���g�u߻�-�R��z�����K�ɿ�z�r#cB��y��p�G��H���J=��)A:�+��
AȐy�	��3H2B�f��n�r���D�7n>�I"��В�X��Ɨ���v���|gkM��s8��/�)�<�f]^�B+�t��9��_�i7R�(7a:�'J���i�_�TJrLEp|�Q��f��.�U�GGg$�i��J�;����Et�k/�?n5|$���ZM)������ ���.�6{��/Gm�+��� �K�PY�*��-��ڞ ���藏yG�k�4&�������l�jƾ
w�C��7��/�Q<��	�E��La��K%���QH~�$�Py�$�D��o��u�(����!��f�Z9��"#fZ���ӱ�'?���?�,h��H���i�>�ಁLV�{��@T�c��#؞5��{��K��[Kk��&�
ݻ��W���D]�P[�Lp2.�4��FniT~On�D^BV�L[z��_��L�M���gUȡ�ڏ��g*�����yha��:�\^�Y�[�Z3����PD<2!��}�*�����P����mG�i�.�&z��8�	m7@�u��n=��y�<������V��Yx2��7  �r����b����s��q��f�y�ple���a:̚y�^��vJ-��b�w����@�2�ħ���X�qYawW<4r_�	�Z{f9IwI��BZ��C�`s��ɏ���(ɱu�l�&%vy�0}A�(.�' �Cf:)�ў�Ҋ�Q�TxFm�7w2��
]��:ӏ{��PU��ڭ��l
��ڢh5:��ր=e�,?!�H��V�5������u���+��A����4���!}�w[.��N@�XϒO"���n��C��T-g'�_�M�iɽ5�Ť�}"�V<Is��+����(eT�;z��s�	� GQn��YEd
��h�r�ˑ�U$x��m�"����̨u��k"A�>��� ��#�a�V�1�F��Y� �x�#C�C��f~&p44lÂ�����v;�������� �u�ؚ��V�X(á��~��K�z�@&�~@,�HO
Qp�غ�Qxq���ɞ
��q)�fk�m㨐��rI��H�n��oD���q��Pŕ��L�I�oE�POOʫ{���o�ds�E<���:��EI�(ܲ��#�ȥ�J���Nb���`Ȉ������~�u��#�bK@Q>��3��Zg~2Z�Q���b[P;��~P9�>�y���z�f�DE,(��7+��M���v�J�Qح��d�z>U!K1���CI)eɲĐ/�;q�L3ُ�3��o�(�n
	��Q�������NL�#����:��p?��b� [��O��T�_+f���m��^�<��F�G���ڛ\�}���8���kr8�Ҿ����;�J6�/7&�w��lu�_�>�r� ��pc��=/ưq4O>���7��L{�.��W��6�O���������L�E�V���3w�����z���8?V��L6�%=�*=_��ۥm���a�MM�Bه)
��"�gi����X�+*��e�"	Ǯ+��V�!�
��F��qA�_�	law�q��)!0Nnݪ,əl��e���8b޹@ɤ��u� ��KKh4�&�ǓYJg��fV���d�J�Ҙ)���04�V4��!��z�����)~�ܣE���A��Yj�nT�����!N9�AZ�;��>i{{�;�$�^��'PL$,~&���ε�����'�U�r2Gl��M��x��m���
��#�HǄ�`^��~���I��H�տ�+B7���}�>����%
�$�WTr�94�c�ё��A�c���͕�T�S� ���l��G��K�Kx����q��Y� �屷�{t���T|v0}~"�1n%
2�of@*������gi�R|^C5�W�
L�"O��K��N&OY�b�ӡ.O��<���<v�d2ŏ�^��X���x�ta7韈�~D��,�B�#��I�G:<$I�u��q�Z�~��G���T� ,����uu�:�S��*8L�~EC���Z�O$�YD��J��)�bDU�
�9�η��� tY�H��nQ7&JH5����=+~�!��4x6��	S_�e#���}.�*	.�$��;v�g�����$��ū�y���^�Nk������$����L�|��4���?���G�s�ɽ�i�@)y��ݡ�?M�Ch�����W;�yܵ�E�o���LB���W��_֓4�RGt�Hy���=T��J	3��}��T�x�F��7O�鄳��^(�t���~jk����܂�q�t�_:���^�'G�h������R_O��Ø; @��?4����#����^᚜1Dɍi6�ڪ�+6!{r8���لR�'��K���A�@����� �ǑD%�U�4�Z=�����a.)�x�7"9~�Q �����_��Y��7�g�tVJO�X�r
nĆ�͟�,����hЃ����8�c,�z��D��T��B'�	���X�wY#b���eE9��(��� ����cX1D�jv����	��'y�B�@Sx��S�Q@��a&9��Y{м��X��I��.f4���S�	�*���P�z��e����н����@R�����v���iDv	�b�ۅ0����E�P�4۽א���f��BЋ�����Iõ��^���
��̹-8!ͽ���š �_4��%�r.��b��I��F�|)#@m��8�U��'���E�C�@m���ݡ�7��k����G��L��{�*�!�z��{�3~�}�d�3%U�	��;�����]�%Lr��nM>�+�v��[ ���}��PFp3�?p�D�Mߘ�G���L���T"��Ek4���V����B�z����>��iG)+�Zܮ��S*2Ȓ�	'�D��N}���~�̐J'�q���
P��n�y7��nz�|"��# ���B�]��a�֏M��t��+�f�%R����X��&/G`4oD�e�Wo� ��h%|���`�۹;g�:[
��j���|����xc؞��#P]I�[�W�x�M�\����BN��+���(���#��ь�Y���J^0A�Z 4���i%u����'��g{
/�5��`�,��$�j٦b� ğ��Կ$�AA>�{n�3��ic?Ȱ
�%��_ы���21����c�lS�m���� �w#SE�i���~:����,�#^!�5>KU��:oO5J6����e+kR���^�8oXC��^׎[��r�������(��]��	��#���l����yt+A9<�҅:yb�����I�^cr��V�rI�?2a����f�mBL�lJ�P�����~�!�����i��	��9n+�
�د���7X�&5򣠼�eǀ`/d��f<8���r�˵D�����>�	X�W;ԕP�j�=��2X�iD9ިӞ�giI���E�1j�}K�G��B�H3�}�8�̩Փ	�����-�pg�:��e��-�t�[���	;
dx,�����6�4�N, �_Ď���?�Ty�b#�ƅAΧ?�RB�rS�r���%�%D��,�YH�[G��v�6w���}��G��T�Gn�Y(�M-[UbwH&9ؚ�<r�����?��cо�!	/J�.m�p��~�i�M�#��@h� �9O,7�)���s�"m��ѻEpm�{Y%�ֆ�9A	4��-��ĥ?��ǨF������ g�\d>�h4���4셔\03�~�� ���� �|��lw�\�Z�H[,�����7kn����eU�e�]6��H"f���}>����/r�����.���OH*���-g����d$��.��Q��#r�&}�}�{�TV���O�ђ U��4�B�oM�=+Zw��9�(�Ѽs�b݂��$��=����3�$��	n_�֭�$��x[P@��'���u4fRX�&�3�ݔ���HT~��Zy�8u$�U	g�>ܼ4�fZ
������}n���G�t���*����j�S ��^%��m��cPkFY���o[��C-|���旇I�4�S�,J?�i���d�s)m.���ҡ����t�=���͒�ͮl����
��Ր�컗��yq������ăҵ:Zͥ�J�C����x�^�vJ�$�m���lebNrS<�M��K ��.c�ώ4���k<Y��}��:G��8N��v�t3�b��t���ꕒ�s���1}�Ō	�D�DdT�gH<�	w�h��/�^�����" �gɏ|��X�o|ꏸ��S�r��V�2�_.�����D�
0�F���?/s��p4��~����:�T���ō,Rc�
!b�7 T�P� ��>?�4��H�۵˟w�<�8��D�ډI��Q�Ћ��!w���<~y�1~�@yd��w�]�)���@�~�{U�^ \�&d��|x̒s<���P��vOpfE���	Ml���fS���m{�VD��#b����yJ;�y������3>I��/�<�.���f0-�;�,6y?����������*7��@ʩ:"��J��34�G�"����녮'�K1s�*G8��^�Pt�_@�k�A��q�Ǿ���>�D~{~��I��sS\.� <�����p��=	�f�+o�'��_i@_>�W�G�5��'`-�(�����#�֩ �B��������L#wJ�s{�;�uy����]�h��p-�4Ĭ��[ߊ�t�4���hݮ]q�B٧G)(��7A�v�O��t���6t`$��N�t��+ǟ�$i�E<뼄Й�L�޷�/cj�A���^����Af�F+LfS[[�'/��jFI#�Ø�=r��8�,J����us�ix������,]�zYa�E���)������j�OY�F��v��RX��Sg�} ����������}"��Mj+�h��?4��4��v��H�0���2~�!��G`�P��9I4��A僩�x��^4�?�<��"���\�!���
�`4O4C�ȿI�����y��h���*z;��z16$��Z�"�J�����H����m	^�� B-�"[��L'ݴ�����J ��W��*,�
-�8s�!�z+'O�uڠ�@P$��o:�r�k�.'�b��,t�������̶g�L�����;�ʺ��S�r��¸\�����6��>{eI,�mv�h���$/�F�Yۢ�ϧ�mΐ ca,��38^Tע7�,�3ij�>���=�&q6�Mؖ�L�L�,�r�$,���qǀYyS�xgK�)F��2G�|��#R�-q��Ũ3�H8s���!�O��tZ-Mi�b\��0חn⯡�����,@�zM��1��xv1ڼD�]|#�퉯��	yTd��Wﶍ�T<�������U�c����\��'�{"����-�>�>[�� %������#���I�����s��[9�X,�������Y�t�j����Ӆ��0�O�ӞH%W]��U<��r��"?P�%�6�#�n�ZR�-e-;������NZ�(�f���e8kkGp�8���	S�����Oe]Z���|3b5��y���3!lh�y@�ܢ��4����簴N>mL���j|$hI|'��.LTՇ6Ʌ\�^pW	����ض�>^�����҅����nε�;�,���_���8S�iV��S�{��X�A�����Y��Լ�
F���_ƚ 3�U&�������S��}5�BB���$�.�C,E����Y٣AZUI��U|��G)�t��K�Sr�5š��-"hL���!�f������A��q��$kh�s�`u'Q��1 �_�!�t�������Ru`������ӹ$ң�^��@��u�)�h!-�6JU[�(ee���Z����wX$ψ����gI@̦^��KƂ��±�ק�@9�8�	���q�&��=�`�Fa�+%~�7lu��{�r_@��&S9~=�!T����T��7s`t\GOÊO�q�������p�?ԶOX�����p��O_�9(X�F��i�2�F#�&jOG�� �ɷ���E�{ ��n�g�{B��,tTD/�@qi������)�^ßA)#dg̮�Xp�[g�)ʧ���c����L�f�>P������YS�x�:�8o�� (^;/�_��[K��H��
��ȵ� 51#��٘�sySC2=��:�T5B��_:@�5��^$fO���<tKNB������-�_��Q/ɞBM��`#��zA4	W:=�ŃI� �9�1�@=vH���ȶi< ��η	#� ��i��["�u��tD����\�	!�b��H� +�&�n������CɪO�CG�Q�b���{b.�_��
S��B{��K��������<�#o�P����B�i�!,����-f��I-W�C�?ĭ�6��� 딣jE�}��� �IW�a�?C�'?�������i/�Gq�QV������b�X��MnU�hv�R�n8w���>/��wG����G�����4M%�~����7�G��:��q� E>�&�aI�A�E���\ann֙�0����d%���jy�<���m*�٬y!�k!O\��GX�&�N�\� (!%c
���&��A�̣LS����ĝ�E���BҮ�	}�]?j�"����.k��͜����X[gg��x�_&s(p�e�Y��`԰
�8�|�9������;��I���p]�-t����G��������|A�xH�����1�)y��?�s��5
fm�b���{�1�Х�I�pFw*���6��_�4�堾���DAb����h;=�Y��f�V����2p�^�ŀO����WN~r�c$@���9�+ϫ�*T��kD�?+`Spe�*���eq7�F��y��e`ī�6{\�7�yhR�:'�j����U��F�`]I8�)� R_G?��,�m���
���g�/?��kI��(H���ƠkLs�E����,AL��8�?'⏝�<��{O��w��]CM3�1=-.���+iN����T�z���h��C���@�i;X��u��yl(���g���9�n�-]�ݢ�z�>��4!�'�n������7:Tl��, %�����A���R�!_{�����%�����y�C�ݡh�p��w���3�-�7�S�K������y�����z�EL����[�O�tPc<+����@�u���;&m�i�KB	7QW�x,Ū���A��V�Td��<�|l><Cj)З��+�J>�*p�����/Qe����Oީ����8��hM�G�ﾣ�Bs���z
��_P��o��ei����Aq�8r�f��y�o�շ�φw\rY��5�ၟ��9b�l���P�R��D���5�wUC���a �`�^�)5(Dd��r!�5�Sfc?��ɋ(E��ڷ"� ��.��'�PYFD�G�����#.%��]5h��V��,N&$�Ll�e�0�����J�׶���Z�^D����hᮡS�KLX�s&��Zq��몀T� ��ܸ-r�:2�� r��<A0��d�@�!�!�Ip�{��u�䠮�F����V�O4%O���ZӃYG����K��º+�N%��/"@�Q������].�Dƿaq�!l�L/>�Is�m���ў��Z�貲� Z��w��((�\z�}!�@Rs�MG�(j$7v]�*޵7S�O��)��,��fĚ��� ��Y"�p�^V�~��J�*0����/�*�������)
"�L��a��Ec�n�٪�s��� )�!)��_d�������L���/N4�l�����_=��,C/�B'��P��T��I�o�&�̙���Eђ��s�t̠��y=��&Ѣ���k'��������I�Jw��K-��	�Q����	+_��X�{Q�H���m.@R���1�����k��2�>��<\�0�̍%��mNk�0y)yY
�?KZ�ۜDW&ԍ���������ȟj:��w�I�Mr��9�9�ߜVCψM�n:s���I������{?�r�����[O�Cj�v���gXY��~xS頢|�%�~����3=~��I�m���xG%�y��H2G��<4O!s����--�il%~�6���X���jW��~&
����?�+M&h=G�Z���'&3)�~���/�h�߸SJ�о��kڵl&QYv���0@�]R�p�rD�D�!6�W�UP�#Gl?��y���6�sF�`E��̬T�;���£��:�5��>һ#u���x1W�S2�XѫƉ��#��7��.�a���ꬅ���@�Q8?[&/i�f�c����;�L*�N��V�`_�Ǣ)����7��ޣ!�d��&����@�N���x�WZ7~^$��S�=D�9�(.\�0��Lx$�7�Q��X$g��c����� �u[+|����$�v�,;��W`�cէ������e����;���e�����W�HY?e"���ե��(*\\`�O��?� s��R�����0���8�F�[��.���|@¶j:��/*͜3A�-4�*m�dbvy��'=Ye�{Glcp͐���pc:�i.�gۭl�?��$PX�O�&�װ���x/�����H��h\�����?�T8�9��hCp@e�[r�Bt�d#�[-Ue�qM��/��޴\�C�r0ڥ*��ۨ��P���Zu�]��51�\�@����	�\)��0�ޅ�."o\�:u������_�Ĕ�ՋE#p��쯽*�E���zj�ђ����Q���I->�
:��3ƞ]��~�^�Yp ��*��nՓ�j�*��d��p�xa�+Ѡ&]+����B�ք�q�ۑk�������!�~R�lm�m�N��]��>�W��G*�L"��p����� �4�aե���pD\n�	��/>��h��{u%��ɦ�M�T_��I�PJ���)G?B3R� ��{�-�PgxD���s����# �
���We�t!�C��E?�[�cz[*�~I��qr˕zr��YU��Ï/+0K�0��ԳN��2��c��w=����Wuf{�����G@��tn��U��<)�"q�+W�1���g�/2�ٿbִ�5zȦ�W��{(��O�G��I����§��hu���V5r7�eZ��JC��� ui|���3�(���+qny2��ɚUZ;�}�r�=`��P��bZ��d���k�#dDWC-������0��{�lCU��鶢gz>�n����]�65)s��j1�am]����!��_��,�F�8�5mg�|��f|C����)���I�e����4�<�-�Z������W>I uR=��(O�{���[N����|/����n�nDAGc�\ڶ@��B^�;��&e�p (�wS�����N0�9�O�7��p|�ǂ����Y�N7������:�u6�m��"·���i�Pn��.t2�a�F�����.��?%}'�f���Sѩ7��#�
��c
��fD�X{�Z�0��Xg0�~��B˹.�9� �ȵ�X>=�*`ZV���&(��+�+*��9�1h2��捣A�eG������)9Wtr\�>Q��N ���z��T�pU�m��* �Q���$f�ȩ�x��,�jQ'���.�џ�'���1z��?�]Y!K�L`0�<� ���G�e��@��B��Ƈ��aR�D<.k���H���B!��;D�?]��	!�[SFjGq�yE��:���TZF�ho�=Q���#6G[�J0�����A���	>�wmG�<�0i�\�}��Ĩ-���->K��ļ��vh�y��w�W��@:��o��FRިYT'H�����Vw\�-NB�d<{�F�^x ����WO��F3m"�Ã�]A��5cZy��73�4���>�nC,�	uJ �<���(v0����?�S��օ�bx:@/�����I�@��eڴWj؅�*Jq� F�U{�mK�0�-zo���lf7�?��?�܃(�u�~<�؇�Z��H��=EOohC��h�T� *ޯi�qh@W|̨�?����b���s�)�	m���D�$��F|F��s���#Ar�z��gVB(���������	�5.WJ�"󾿰�[�n�Wz:j�i��	z�˛ɫ�2#�g���%�,������T��{���c^����z����J��l�!�T��?��F�!Ξ�p����{N��/��N�{��=�Z�$%�'����Ӷ����CWF^��D�h{����Nd�����e���s���NP]���|��V��=�$|}d&>��H��u8r4�4'\c[�J���9�89�(��A�S�|2���bCP�|j�F~���h���p��Ԟ�s�XJǧW΃y�C�$  ���ЇÑ���x�F��&^G�͑L�ۘas���N>�mN��K����|K~��Gl~g.�y
ҕ�]�F+VHlr��S����ᆵR�9-������q��h0U��`+gJ�r����Ipّ�L�q MFH��q��<`���~Ab�y��Ӄn�t�m(�;�:hFD_�����ز�E�Wue�6����6�ه�I>!]^�磩/hs����n�ٴ��ſ
�CWF[��g������P�H��(��!�9��T|͆AWg����Bo�^���tP�%��ơ5:�;J�
��-R'�מ)��N�m���h�������j����U����<Y��S�涂���"}����w~V�H�h̗��3��7������]C6qR`e�> ��yYݔ��8��ac�Q�>�݇8VT�~���X^������"K���\���q�#h�U��qըG���X�ca���6t�59�V9j,�����#��Y۝f̶[��@|HtK$I��Z`͜����H-%C��oެ1
��K�{W�@����̐
�#p�k]�������@?�v$;>΢�\)�Q�=�`\7gGY���vK�	�=�x�����"�W�}~�۝:Qp�YV/:��Z��R�#�e`c��P����Нx=�6�*�u-{�������5�<���ϓk�XA�������<��dgʤ!�y��iB��ګr�R���sA�}f���m�	�{蟛�'��h��Y�>�56Y��ϝ�m7���ە�t�
�O@p>4����"W�w�=�'�!"�$��b�r��h�9?�R+u�l=�_2T'YHP\��E"�pR��ׂ���,��&��i�V_�`�%�6X��'��<,xB
s�����>b-'����^��'��w��4�_����谙��qm���¿ey^���K����dI��kQH���̼;_�.A%��L5�x�KC/������`�q��b.a�y����_�Xɐ��5�`-r�eR^^+�g���6<2��B�n� 2ӭ��y�㤽zᐏ�� �**���/�7�y�7����얥7�(x��c��@!
F�+eCN���:E�A\�j�*A�1����"��Z��6^�Iė׈�EOr��O��^7�zäyU��ѪW�m�&��]��wi����K���4n�8�`�Tb��L�h�\��n�S����=�	c���ә#�ń}��;^j�׹K���߼�?$�0j�o�W��m�tGژf���j��|Q�����8#!��I��El,�'Or �����pĝk��8��v+R\�em���Z�Mjߗ�Wt�Ii���wR�B72P�x��p��/���⎊ ,2X����p��H?K�1���˸���/��!89�{Ooc�DZ
{��v���0)�kƾRKFt�!� �\��\�*���Ó~yK)gZ-�0Ԩ�٧�'��"�Ć���%�>��.�M�Sro<-�^I�m3��K�D�v��mo~���9�����p�ɝ�_WX�ϓ��f�U��jo��`$\�u�ߎK��~���������]y�rK�f��j��i���p*���״��<�^�e� �dÆI�=��ōc��؅�^傫ѥ�[���3��/5F������N+[�{��NP�Hr'�#FE'�_�ܪ 
c~��:)@MR���4�-�lQ�5�9�e!���p6+!����+
�,H|͛�>��Ԭd�.�A�MD^��kxV������Í�?��b�[�A��,Ҁ�aj��Z�%pxg/�%ZrЛ	+�1��=j�>���x��}. S����G�J|�b~2��x�m��F6]˭����,�G�1}zoG_�m>�;i�/������϶X���Qx�_Nϔ9g+��%��<)[ܺ�F�Z'�;1�h��l�t�Br���Uh@ղo^�o��˚3$��H�#gM��C4��{N'ԎĢQl-����^�5�5��� {�YAQ����� ��q+q0K:����i^��#BM�.Z��laO�K3U��� n2�,]�(���$�}�]��;���@�����&#�D�y�wL�J�<�&�[,}��	�n�ɷK��o7����?S>�A���pG�JX����#:uN�\���14��Ӻ!${�����l՟�>�}��Sx:�eRY��b�nrW/چ�:Yp�����V3����&�f�M?ޫ@z�X\��3q�ԗb��t?������w;� �}J�(��çbx������w��XA#k(�5��&J�Ӝ��Lr���j�x1Y�~�ە1;����b�_x�kw�7��y�n��2Dl��p��]:=��{���/�k"��|�*IuL��w�ۋ��i������7)NUr���D���W�K��p��&���bo50�"���>Y#&u?�
�`(�����Љ�lF���D��`"�?�WC�!>��Q�]>+��Aԙ�M?Ê����P�����xY�$B��_=��9���M�(/;����;93|L���i�@+hiq�qJT"��d0}�"�-'g����a	}�0E��%CB��3�j�B�!$��ʑ�L7�
,�C/�d�"0��g��JR�������V�}p���
����� \e?�<�`|?j���lY��a�ݸ�%�P�b��BzL�>&��w�c��ah�u��y����K�==�r �7�0���u[E&
�Ҹ�lpm���Qi���ˉ�2.��X_�#�/7���/�p�6�_�#z�/��� ���r��cQ��� ��f�w甲���`b�H���3mt�p� �Dw��s���ꮆ�H��}{��øo����)+�bǐ�����RS/d�+<Scb�٪7�i���m,�t���m�oL�����
B��(��}_V	P;}����܍��yɦ8����B�9eQ#�r�"v{�U b��� ,~�l9�1�a���k/V���3j����;�j�L�A����TڝKQ�
-�Đ��L���;N�ȆGג��{�Ny�Ԅ��.Y��OZ�?��Ck!�3⿖D�m�=H�����o,Oc<_xwZ����S�4������
'��=N�d��p7��e܁�(���~�r�E�+�H�T�!�_7I�S�/|'u!� N�X%��g�,��U;2�
�k���Q����ЮԖ5�A�:M�� b�4N\�)-*X���[�	��Az�i��/��Zr&���BI�Qd���f���/J��̶V���O��(͂=�S*�FD�K��;<��.�m�GG��C�R��6�%x�������r�px�����{<K�<{X(h��SК�1�uI�V������$e���C4�p����rݘh�D�F�K#��e4���\��z�A�*荻d�U+��s,h3C���^BB�Z�	5l�OUlz�f�6]~Rmn���"L��Q��c@5^���x�����H���i�NǳQ�`Pk���V7�V��~������S[�]۾��4�E����^&�d������ �qX}1�6����,�'���A+K~����c�o��9���8�w̫���jd��L���4���*y���$o�� l�K�V��DP�f<+�F��<�!xCw���5�*�������-�Nx�(7�z��xY�e5Ҧ7���D��rZJ�3wڃ c�׃�ǝ�N�R" �6�,�"j>��T�g4	����Zht�߾��BV`�c��@��?2���d/|��Ź����K���(	,>�J����3���úQ��Nm�n�flØ�A���#���_h<:h�1+I�i�:���}ݻȟe���J�����l
f�_ؔ�8];P&��֋�p���d�f�=%[��ġ���m�TM�.;��!�I1L~6�e0.�m��|������I7�4�0��6�	~���eR]MK1�Ҭ(%rw��v�ۦ��.+#	��D	k�z,eU�0�3�ur Ǽ\0q��fUt4:�(S�@Z#��x�FT�~m��e��i��A�����wB�ms�^B���j�%bv��p���k�.�}+�9w�;�k%��Î��xYW�� ��  ��5S1}z#�����:[�ň-�*e��+g�q*Ti>ZWЁ�����bA�G��tu���m𙚚��^
��m��}�F���x�|�;�5O�T����P*�.$(�槹	6�~�OC�y�Ԗ��>B�;�EȊ{,��N�"W#����d��Պ�EK��p,��\pT��J��e�Ͱ%K`��9l��ET�Cj���}����7.'�9�cwH�4�.��fg|Y:�������l'��i*�3��7i�j#e�r	��a�Jʍ������o��&�d��!ӝ�x�|�"bcc�Ĵ���
�
�	7b�b"f��R�>EY~���4��)���� >��8A5�������H�IJ�l�!�����I���z⒤h�����ׇ�$�������y�� ���+kr�UZ�	TWO6Y2yh�}/�H�X�6 i�n�vl(x g�*�]2t`����2�Lf,�UJ�J���js��'�:|�W��6�1����]���"\���C�.]��?~�*��?qTQ�i�WvY�R�W+iV`��;�`p����E`&fx���ه���v7��BR]��Ԧ�!lRo�D ���E,{J.�����i�J���ܻ%�/��o��O���	�E��3�����-�b��P��؂E��f�C���8���P���h�wN/P����x����&�]�a�|/��f�%��d���,Ume�G��?:�a�������H<r/< ����3��u�>mtv�y�i��%}��NuƐ�Ʃ�G�d<��v�<bu�m�i\�k�UO�5�D�.	Н�4������5�Q
�|3������~���IHV�Kvl�[>{���DUZ��>�"�����Q�U$��5o��U:5ʞƌ'չ�M@��K8� �Gp�^i�$��4�Wl=w:)��Q��?�W�k����e�<�����8��dk��۱"o���ׁ�Zc��Tc�i1�Tn�U����L���r@@�B�&s��K�} _Tv�iQ��ȼal��9�-$���B�g> +� �mr�0���^^�1ݹ�}��0ՠ�Ԫ�|i6f��E�H��
Z���p<�9tX� ��E��&�bAZS�7���e�)F=٩$����$��_X�Pt2���|�K�̋dD�2�ٱH�?�Z�L�'�q�� IX�n<n�����GBҳY��
�kHq����7�Ę8�u#�\�[��� ��)�G�����o�>3�:@ɀ�f_��̾ �1YV�d<�W{ޔ'�B���̂˾����[w5��Y>�ޘ.>Z��\�!�����G�6#�M<0�#_V���2�	#�ri�X����t�c\[xHue4�����e�uB!��n��JM-n>�eoo&�{Rc�1���T���y�Sg�l�>#g�����(p|�$����:��1��ij�h:��L� �p���_���tk>4�'bB�`���0�����	��������}
�N��O�>`�N�"[;��������Dm%<z2�o�$Pyq�%�=�5�'�������G%A]���^H�����WWL�W�S��b�ׯ�4 �k��,C�;ʱH(I;�	`毎XM�o����r�+��t@Lo�y�����X���=��L�h��C[�llD�QL���$g��;�H�r����n��������4GU=崸�9��ߓ�:�k�TY�ə^C�M���)��&�>�\�e�����e�߄z�&ps.��+|�^��P��fXh�6pi���K�
^����sY/n��7�"�:dԔ�g�j�d]�u\�,�������t�w`�=,�c�E���Za��Yq��@����;][�����5�����2��`߭�X��E{�9��Wm�Q�݁U`_�A&���*�^46*����m��hn1�m�ئ��w���kf��������%��&� ��f>d[Q�8��\�K>XȞb���+��h�.S9��J�WA�;�֓��q1@�.z2�)i�k}z!�3���[���AyJȅV�����2���-gr�[h�գE�`��5BI0������
�+�e�͒WP�����d|]ӊop,�)d۰0���W*���1Q��xu!����߷mIh��%��9a9��f7���������'d��>F�����8�<�;>�6el_�r���!IƳ&ă0ٗ#5Ug��?DV�T;T��j��b���(��Y�l���P�>ֵP
ղs�sz=��SC�lH�կ�O��V$��?y
�WE��x;u;�F��r_��������dW�J�A�Lb���э(�AZ�\��!~("��� ���ۑ�ʰ�[�uNQQ2���}h�JE��`�S��~��5S�vż�[�:gK$k�G��mi6���ˀ㨁4ke�C��6�R�8��ßIp/��_1n�<��މ�琜8׷;q���,՗no���返�������"� O�;!z��1�A<�\��ձv�k�ӎGA�qZ|h�N�	�=}�ɐ���� �J��aW����Ѣ#%�O_	���d�5��M����](��&F����^jf��
YW�o���ƽ�[E�P��4��gH"\�B:�XZ"���ZJ�|e%��;%j@*4vyv.����h�{�C+��}�QX���XƦ�����L\[�0`�?I&����E�L�/ה����%�:���	�*�݇t��I���jd�{�A^��Z'S}[;G��)��h8�KWm���Md�p$ (�2nx�*�	tST�U���z�bX���{�c�s����Dڳ����.P��p�\Z�P_�C���X�@��&�i&��2��}ڧ[�{�~�N�H.bf~5K�Y �������� K�"���,�C�='�w財�Y�9�#�ɏ��9 �5�`���Ig`.ߵ����ES�lc�����U��8�B��,M��A,1<;�sd�J��{i���y�m����I�Z
��
��1,*�N�dj�-V/�q �q�$��>fn���p�������+�3�|旝Iz�!F��9n9D��܃��0���K��:���p^��£��e�5�&5�C���_�S�NjЕ�6�|�fV�����(�g��BAMF�m_:Uj� �k0g��1+��������7�����B�0"D��	�M��U�SҨ���$�J1�bez��m�[w�4&��HתֵyR8�a �{�<ʙ��=�E��D:�e��"q�bݿ��m�	�#]в�ʖ��o�� �낹�	CE����.n)R�@H��$Җ@�0w{$�o���]�j��G{����ƶ�Cl��	Tku4:�L����6]�{����$��
��(۔S3��j�^�n�>�����{�r���٭輲:m�_��Kox+Kˮ8~���_�v��JՓn���wiYu
��a�2����>�s{��o׵ȏ�\M��U��k�?(���q����ǹN<�}q��R�ۺ���y*��Gm.y��9<�N�צ�I莂ʚ�9�!��B���U�|�d�[�L�΅�q0Cm���{vD��rßi�+�bC1�+��0�%,��w�Ȥ�1W�f\y\}��P�*'E��������3����#��sVZe�&�¥�J��ƫã��~����T�*����^k��LV��������.�Q�3��g��as���~��-@/�b}A��J�W���㆓�fc}G>���Z�iq�*J�ڂ@�͖�ؖ�*�M�zc���Ͷ��T�JqZ��PB|�!�W�Z�I?����sA,�����nx�?����نK��K�=~t��D�#w��T!X��H�72�퓒u�m;���� �[��5pV*�?�֜I�#	M&����� L9<y����	*:�&�Y4���E'X��Pn�w3��z�'�㞒�"�`��(�g�1��Ɛ��П���>�3���}�;Ŋ,c��#�կ9�F�O��=�[^�^UM�6g5K�����]���z���ύ�o^�ш�5� �;	F�ՠ7�o�k�l��u�^�o�%�6�CQO�zX2�+4m(?�h��)+������s.�/�E�KF����?��D�l���Xf|N}I������^?c��9�=���a�����G|nO��d�� �'����
�kM��EQ��q�M�*Q�p���hG��W�߹V0��hؑ�y˽n�?�L9]�cS1�I��J1MM#%�����O����}Q9�3C�UO*#`K�P�X�{���^94C�|���t#Q�K�ń�#�r�]�n�iz����Ad�[��3�#\�L(����Rӄ�]rc����T0�Ӿ�
�O�j���ǌp1j��(>3w���Ғ�7��U����ά���U~Uu��U��2��P���A-�(�
�Q����T�G�@$�\j��e�¼�����nM��0�èaDV���Qzъ�lx (0)&P7���,�"]�$�!�G�P`��3Kճ��m�Kw*O=�����)��ϥո��QU�aЯ�:���7�o~�bFx
��~�HS��Ce~�$�����Au3�7�2��"ﲶH>�:�['�:�՝�ߛ������a��w��d��% ���AͦkI&��?�1-Z�8�ǇX��J���pK�*\ln�h�U���2�T{��PsJ'&SP	���m�&}s�uP��ᨚ�=]Z	�4|o?�~��^J-�jW�[�"����S��d�ۡQ �G�I��̴�bh�!>{h]�ab�i�4B�nk�ta��'|}����$[�<��J &O�|!��^fEGU��:��vN� x%����vy�+���s����b��9�m�ͨd�я~f7%�ބ��U;��j��G��s�q ���3��k�H�S�U�E�x�%1#��{��q�`���e:b�2�i2ж�l�E�F�ӥ�'��V6��2�F����6`�ɥ)lZ����x��1B��,|���i}q:�����t�@"8n�_�$AkQ�N]�Y%�V����D�s��XkH�hd�z0���U�5e�8sE�/�:�-Vr�*�G�[��.н����k�Э�R��;���6�J����.�6N;�)����t����U��(3��A��;��,y� �w��	�۔�b%13��I$+�����_�����9�#��,���O��
88H���b@��A-��,#9d�r�m֑����-e"Ö#�\����r~�?�:Z<˙L���Po���U�o��Y%����jrQ:T���ʀ�8��ۏ�yy�h��8��d<���������@��tƖ��	�Vum�$1B�e�4V�n�D�M��`v*�I�帾�t�VL�bj��ǣR*)m�s5��i�d.��*[���Ҟ&pˈ�V��	�^g��\LL[)��.�jv�b�|�D`Mhb���E2	�FQ��	́�⪜�J�uK]�n���x${���$��?�-����]��s�G{r-Q }�E��e�>�ʣI�$MA���L^��Kp��5t�o>���u�:ϡ"����u�l-a��a��G�Q�q�w'4��!D�g<�Lk@�Ȏ�������Kx	� �BÐL6ֆ�����ٖ����Oύ�Mn��jR�*ǘ[[�5�^S_�� ��O)��DkIX2��4'?���d:ٽ�ao�5^a�e%@0qF�j���n�o�, �c5�D�ɵn(�䂸��׌�^M�� 0�i�Y�	`�L�"ʍ�D�J���b^+;X�M?����J�(A��At2g_�Cȷ���^L�� )S�}�|�_���cUZ	�R�ic3 �g����&�(y΄��P������>+�hH�5���:�z�� ��ʚb�-��4)ģ~��ii�[��)!�3���ÆA��\���{�@p�����v�Z�t"�qE���8�^�Vt^�* >j�>�3�����븞�FwD�R��-� �3$�$Cxwru�q� 1~�w
zsW�:'�s<��e��p;�o��J���~��`�s��W��(7�k(�l	�nCʝ�4fFfs)�>�0���i�kml�bΉnTQ)F^��a�N1H5�$^�b��)����� �� ���,��<�A/�8�� {��b�!b�(�[C�拴i�u%kǗ�[b�\��y�V$yb�������Go��/���K��I`����0V��J��U��5�M�T�[��	0(
��K65c�3�KN�*�H��<m��� �h�Xݗ ��B>�.�
�e�Ei��62My���#�πQg�}b�~S�Txp�Z���l�"���jk�r^�:xW�E���?=<��Y�3���}D0R�lBԊ,B�^uR���[��
���}?aT���%U5	DIk��J�ϓ.w=�(M�T���hE�hYk�n��c�O�7����3t��8�T
ϋ�Gg�;����z���=z��2}2��vC�n3�����]2yt��]Ϝ�&� ɖ侾 '�N	��%p�C�`����fB�Ge_����@Q�0��Y�mkF"�ie��+��׫M�ݳ�Ʒ�u�\##������u����$��T)[;l:B�2F*5h�V��I#�x	��/�Zu�'G�|�;<�~�0VnI.��<��=,V�&C2� �.�a~Eg��)�)l/�����F�,⹠�ڍK�f?Q��$ё�H����8ZD��FD�҄;�Q��]�	��{5�؊�u�����6��46�W�L ��K�zCt��5�^��2w�r�x��x�}޶�>�q�+<��9��&cy����ۤ~!�t8w���>�K=M�4�/���a�$�4�6�-a��r��,Y�F5C�;��R �Έ߻b��Tf����V@j?�eJQ��F�V�sM����;��-�zS�� :8YX�>HL���<aa��>���6��6VX@t+�)C� ���K�K�Y� �dQ�E��UT�G~t����~�qk��	+��R����)����O��{S��O�!��>��zN�·�
QC
���y�ʅ0��`^�������rIb"�)mƱTu���|Z���]���������,-���*�s�o-G�ñ腬9�������]���Ɠ4��$_��η]���(;S��{��s�s�`�DYE��jX�Ow��/��J��mu&2ϔ.�)�LI�b!a� �����9�rV[����U?\�Q�O�I�R�v�h��<`���5�m�#��^F�dgP��µe ��\e��n��h!�Q�Ǵ:f7<�%ͧ�O���{4G�Z�-�9��ޠ"Z'K ��AF{��0sh�o����'��h����D}*Э]^����)���D,{��L�UL"�J�w��󨙹}����� 1�"����8f�^�]t@���c��3���k��-���[Y@Raq�%��0S s�D7c�k��D�Aͣ�h<�UV� ������L�H( !�aba"ڒ0.
�-L�&�*EH7�Ŋ��tϭ���T���g��tYA��3x����1�2?K�_>;�r��WGQ�q2�rz��o���� 4��/l�vMt!���G`�.�lX`g��F�JU%�*r�G�
�<��dO��C�;�+V�'�~q]� T�q��4�y��C�E��*d�Cz���G�\�TA2��xfMa�&v�90H����1�l�E�"D�����2@�\�s���h�i�P��#L��p-X���x��	�H���I'� ��J�q�X��~��3]Ƿ�L@�.�)X݊���\M�/tYq��=Vv :�h���Bǻp��M����iw�1HZ��hA4����)�Û�Z����@�ڏ�	��N �j&�%(��� �uq�o �D����V�����jv��P���sv$����=v�u��BN���:�q��75�jB��j['uv������#�lO���G��
_)�O�Ę���_���.�[P�K��\?�8¬P���]��H�֕#���@��O:+,a7��R<87n��f�LtC9M.m��ؙ��"1�
b��	mm%���:m�g�~^[�E/�����φ�=R�n}�Ct�UA3�|Q����z���v��G�ԕZ=h�}��jPF�B�8�G��O�Ϳ]��b�����.�U�݅�R�Kg[^�ϳ�!��R�-	��#�$8�I���/��d'1�z�50�� SM��(�l�H�_>��C� ��Pf�)�8���`G+�V�H���7�N\������o�C9̖��7o	H,�U�{��6C��f�=�_7Z㪴�!�(�g�?VM�����X�p�n�!m�;
���5���\=�"�<��b#W��G�������T˿Rΐ$���j�u��(_��_2�fWp��0�}nk �GX�rc��j�ց�8�r<I9��,(��������z��(|_;.B,K�!�2�ũ)�Q4��0d���[7g�<����,��6u"M8A^x�3��T��S�B��5��C�@�F�A���iM��T�)6%����U?$�������&�(�o���kجč�M�:�R`hQ�AG"N�e0/hB��yq/��ڪ�{���
/�XN��3����}\�e���;(�e��џr�r�7����j�����.�<�����Hg!-��c�@���nh�8m>��5�˲(�0�"iv{���ɬ�-�P���c�SV�{�+f��T+D��2Z�	{i������5��fl�1�E���*}2z���9Z��*�U�h�������2����ᯥ�=�l
yB�A%j�ɫ���K�W��6�7Z���L�AAǓ�Ui���Kż�l�"?�l ����w_�E�Z��j����:)B�@�TE�6D�M�ݱ[r�_�2���0��oh$u#3,����&~{r�V��F��}��чr��7;�ׇjGw?�ZD����T���ƌ�~��&��F�(D�.��9�[�����#90�&95�DϞ�k���r�WxT�A���.oo%8�tkg�������ؠAp5	ɔh.+|���?o��rl��&=��2����{�3��^p���țt^!�������!~&���A�׶��튽�r/֯�?od�F�c��8n��ΰTN!H�sK�N	cgG���A�o���\��l�
���:U!�W����p^ �� ���»AoV��$�����P̝r$뼙O���X�<PHe�
�4&�<�����"6�8���v�e��c쓝�z@�V<%iK~�A'�ɸ��F����2F�WB���T7�Ab:��P���q�.��v�<����������:)�$�k�cgs�">�i7�48�(��Th�?�=H&��d��d�*Y��SB�ט�o 7wJnqg2d ��;��h������� �P�գ�.L�+q��e�����0zN�3�*���#5r�;w�T��{��j��\w(�I�F�{�у��]w���F�2@8TuբRm
�Z�*�y���Ы�-y��X��Ӓ�P�Qy�[(�zb�z�L2� 9,{ٕU��]-w�t��?u�ck�]���}�4e���ݑ {����:�^�b�C�Ջ*(U͛��TKH"�Z�`�on�#�!��F�slČPӱ��r��#Ro�9M<=.�JY����W-���\*��.O�+��|�M>�ؒV���n������xk�R~t�Q��I�X������C^[a��ԭP���>�����|����0]kЛR��9u}�Kk^.M]��#&�1dͬh�dH�����ݎv5 ����$��bB��d͡��k��eD�����\���VM`V��W)N�v��K��rC���|[Dw�TQC[���z����s�Ǫ=�H���?>n���;�z�{h�ZBB�H'6����J��-P��m��F��N3dŬ�{07=FN56Fqf;7ިĔx3+C�m@@@������]į��,n��5�`�]��S�;��l;�K�!����ˋ���B����"z���r1#́�-� ��B�5��-���Ἧ<�c��n�!7��c��d����:��P��)�1*�r=3j��T�@&��5��P��x��}郮E��BNP�(1�w��y�F�(zɤ ��p˫�<���S��=oǍ*=eʥ�>Nl�]a=A��B�P��ρ���k ��S�il�њ�D����u2�?k ,��a�B߸�y1�d{us@��Φ[\�?�D��~p�Rǲ�f�G��p��b�
 J^7�4��2�F�ZN�1��c��ɿ/�;�� g[<n���ik`�-�nN4	����lSGT�U��p�2ӟ����x=ڥ*P�(v��;Oٰ]�)
�zb��z�q���G��""�Թ`��՞��2|��+jA�]o�E���''A0{s�P���z�Lo��&��4#�k�.���u���U�M���.�u�e��U)�L�8>���L��i�D�@V��K8�p���{C���zZVD�_�"�]v�^����=)���En��a�J�8:�	� �ԯ���ߪ'�����J�0��^\,sn$J�@La���ƓB�b~ʿ�;ΪW�f��/�}�ۣ%]�;8�S�J�R)f-ԓ�<kSKr<*	��J�E��^!L$/z��V�֛��z*�@חŻN�>>z/�����$���=E*��������X��ڠuӄQn�n���M��n��RĻ��'��/�>U���5��}�,r��S��������!yMƃ�x~�7�2��	FxP��x���ma�ވ��F�s.ka���b�볝h�D^. �ߙј,Fi�=a"B%��>���U�d���]����n��EcIB��Z((8��Db�,���sV������1˘���`CH�Wh%���}*�%V*��]�$]��*C$�$\'?WԷ��l \ĕ渍fB�szi
�6�A������w���_Mƭ����;�'.y� �k�M��W������s��7��ˆ�b��H�bH�0��{��2°Ӯ1O�vM�ED�u�'e��I֫S�܌��D&�1�bA���Tfw}���N8,�xl�.?Y�������;t��� 22��.��)ǧ�����KB~���$�c0�L>x��['�������M���>�D�x�(v��D�['�"C�S����VT	��18�dC=5J +-��*��Fݿ}�@��
�1��~PtH H� �k�sN2�,}�}��j�:���$%Ce�U����3��1���s��ġ�чm��ɮ7����+����Ϋ�i�y�� ���-�E��V�V`��M?�����m��J�NYЛ��d�\�{�,0J�7�Վ+�V�Ƥf��]T+�F6��63����(��8���,.Y�QuT����fhkڷ8������З��SFx����H�m������)�G;���L5���sE�|	t�)�OW6��N�kMp����8E�6�����X�W��14E�T��z���b?XM��W
�4��y�I�§ʊ�$@����0���e�3��
��н���p�qn*�Jy���?|[�����c����P��S�Okr��}�V��^^F�� ����e���G����F��S��g�$�\���ۨ��0�P��F�2y :ց�k�c�h3
L  ӕ�S[��~���cl�H8�/�ױ� ��Jӝ��`\���,0�b��uy�"�X(����� �h��
s�]�1�j���@(|tj�":~|p�0����e��C�{��bl�0U��`����p-�����-����n��k�����X�R>�D�Blj��pf�c�z<P~���؞-�����I�b'����-��T���Ӻ{
Uի��L�RD2�B�z���`�	� �r�Ѕ��)��)���F�T�hl��X]��2�F9��l� ����$������Ũ)�fi�SH~#��|�����bJ�$ҥ2� qz��	bf��N�1�#�=��VM��Ka
������z���g�k�!]����6��]�-��H����̪ܸ�k�}��b^�^���c[�J���7z���h����I�/�`���Jdy�wz?��У�����*�P0��"��jXWe��w��Vܔ_�F����\\ ���u��D��p�V�%����?e���%���KO�nܘQ��?[-��w1;
��)���X7�O�PP����c�3�X�/t��X��f�тc��Qi#ȸ��5���,���+�(�Bѫz�S��$�*�UdB�|qs��<��e���\�WC��2�70�"i���r��F��t �|�ӌ�A�D���x��+��L�D�Z"u��euk�\�o��}}�!�;��ͩ�<C�Dm�
rC�SgC�R�t�ͳ.`_�΃ IqRɼ�����[���4�
$ީ�9�V�x�R8���r�q��c,����I�mR �����x�E�Ok�0�SU��cȒ�ۧF%�D�֗���X������S,*K��1%댓��Y<e ;+أ[�x
����k��i�:iUKǋ��`N�p[Y{����	��  R��݄�[@?W�k-�kK`�K���l�D쑖%�Ek]<�E��@~�</���8���_����M���6�8��-�F��i^�����YJ��hH�@�L�l�@Ȼ;;�{DW� J>�)�R[�'��0`��W�5�:"��߈�p���(�C�Y��80Yvv�^���#���x)V�jb�S��m,��R\Vs5�ieA'$v`&�L_.�}/X��P�f��Re�f�����$:p��R���w\k1T�O�n�I>45�#'@�׹�#��]ؑ���޷a6Rj%	?��5��{�Z���6�&�����F�}��BQ*h?_�@h�~iy��ڒ�-y����J�����'S�:?C��Y��y�c2�[B#7�%��B�x=��_a[`M����؞�'җn�fq��ѝ��/��3ѱ����Ĵ�^Q籽�E�K�+���г���W�] �w���n�7���C�V'�Iy�L�R�x��%������s������$+��D-G����ʉ��R�Ԯ��d�O�:.m��L,���W��d��ɍkyM1�i/D�\*qdm��<�؞h�&͛c9� 2t� ?�2tXM���KL�Y�#���}��~?�i޼K[6X� p�8�s���=���+�o_`�W��L���23{Β���H-e"���������~;��>�k�ߒ�wz���j�%R@]/
�bz\-=E�33�U+�2{��D:|L[��h��ݛ.n�0��`��D"�^1?�0�l0Q+�{�n-ڴl���ꥳ�E�p@� t�b%����]�>�1�Hc�U�5��N��Kj��h��"O������c�F7Dg��խ
�c<B>��8 ()WJ�0���_�	�� ��o/*�~�Zp�q�T�n��E;�?�Bh�������b����$��t���o-b8�2\J*�T�E֠B/.�X��["�'�_�o���	?wŴcG��oH-�.{C���B<?_���')�!t >_[��͛��"�'^������Yo��D>ҳ��[������g\��}�CD���ds��dx��Z��;� 5`
��?s�ܻ�БxT��9��ѻ�lR���r�:Kh�����ƭǒE2D�.�*l��8�eAa���q����S��v�d�PZ��@�/3���no%|��WQ�{�����<d��$nr�'� �N���C����T$q~��k	O�G)�͹J�R�[D���1�F�>�sjW�v� �fn��K��0_�l^^ ط�_�8٩�7I;��ȇݸD�iQh8xCWy�[A蓬ۣau2�5A�(��G� �GQ��ƕ��	��t�Iv#�t8�p�#l%lz��vŔ_������%	���'��y١�ԏ�� �m�p��?����C�mZ�`X�lw-J����.aS��Դ�ii��6[����K��>�ų%/p�v"ð\��Ƒ�_�X�����!9��l��+�w�� /D3]+f��.��؉�(U`?}�3(Z���hq����F%<8O=5u�D���W
 I���n����9���4�8%b�6Ķ%��ߨ��υ���.��̡�`;d�4�X�o_��i�����:R/���ѥg�9��ܖ,~�y�͹Ă�2���PKŅ�
�Y�(K5��dA T��c�{��M��d�c	f��l"R��!wH�y�S붝(��*ĉ,��&Fl�����%M9R�![��$�(�h?|��(
, ]2�_�H/ŲÎn2�C�gU%ɲ�L9��{��z��]�Fb֣��Yf�2���.�$�g��p&4n�K���m�C8l�'��a�)%��$!�u�`G��Zq��<Df�˱�Z~��&(��61��^�2vX��D.���_x���������HZ�9�U4�D�>�9I�>�?m�$ ��c!^���I��"sxv�&�/�y�����w*�R^r��h��z�R!k��~sYƯ2ގ����FԴ����3�Z�U�P�b�J,g.Hs�uU�+�}�ZFQ!�����h�,"���$c&�������{����L�r�U���U�r��u7~Bt��	��0��,ƚ���ȡYEhh�`A��S�U:ë�����ye��lM�J���aZ$~�r��A�L�.��������`~�t�- |e%�-	�?)6�g�E��N:���P=��ŕω�	GG��M�a+*tV��h�L������!ۓ��-)�Q=�E/9V7u~z�EJ"���Aq��mV�J7����A����fL)��z(r�6���^����-~.�X�:�&<�6_�����V�f��ޯs����߷#	Z  �rXd	g�ne��M	��	����@����ڽ��G�4y��6Įr/bx	�g�t�iw�Σ�L��W^���'�Yv�����P�O�ثd��b�̛��<���$Fc�F�����c������j�U���RK{~@y ݤ�A��hu�!J�EY�旒������濊Ԫx�#���>����t(�#�e�($þ"6��0�H��n�<J���0����HV���0�����/��ɕk��v��*�)=���W�Ldà��+�*}�g*V]_]�j��� �o}{%ų���������ip+�f��2$�vO}��"n
]��I�?ۂn��fE��(ٔZJ��MV�/���|���y���zdꖢ/��l�6fy��]�НP�7'$TGqf��*yޱ��!��Z����Y�C܁≀e�ٗF�-��0���ڲ{%�tK��>S�*���~�U�BM��-��$�[�׈b�ߚ�6G{��s��f�7���ró��_i���j�Y��ۻ�!I�nS��$F*�;W�{XE�E]o��!�e��F2��׳H�{�u����q��c��^�(�T��k�ML��	��o%
򉃯	�Z#lV�m9J�0 ت^����ɯ�ńgg�͠_�ӵZ�.��2ᄀ>2UuǴ� '���S����Fb��8�@.�8�ӆTa��ᖨ&�P��	��G%P�):��3��cu*��#e����{\�iܩ���u��#�Qt	͘F��X2��P@CͭĴ�����0:�R!�<l1΁���0����1#�/��q|�����+��rʰ��o�*N��-S""Ng��@*I�W5ka�o|��f���P����"5�u��3V8���!U�сO���	�]�m	�{�Eۿ��?LW��<�J>$,Rz̘��{��L��
R+���`��Xk}�Đ�L��r[�o�i`N*�D ��(�iXɎ�T�ZR�z86`&�y!�.�%S�xlG�U���1O���P��?E�Ѱ+[�e�8-�c�3���M��A��Gٲ�%�!�*�%&��'(�&fИbXO�:K�Y��7��k�C�')#3}	�|�R�E�!w�0cÖ����H/��ǍR��ρ�ϥ� �I�H� ��l@E�D�xr�l�eP�Y�8r�%O��>f0A�i(3�;7o�9�����}�ӷX��aW��V��a��r�^�J@�h����q�m�퇯���%.<�-��a~,�51�~�b_T�C�LwJf��fY-�Hjgz]+��kW��g�!�β�v�ꠐ�/d��l?0!��CH�p����?Q��FMqv{`�X����4�v[A�a��s8j��oD��K��4B|��-�~�`R8�8��x����ӵ���xNz�ȳ�� u��{�QbNL��!�fpv������j?����r1І��T��iC�?gؿ�����;�����3^�U
3�G	�%4��̳��j���y.x����hĎ(�Y4f�ň��)��]u��"[�{2*͚��c�"j���r�á�B�cp��go�)0-��-e�Q�z���~3�Q1йqe[P�@ڢ�7�-�w�Y����;W�W�w���[b�D�W��g�OlGzt{�Z"�n���.����5��HNY���������o�����1pC6u|���^A�i���4�"����J�"d&x�1<��Ӥ�t���^��_��uF+�����5��H�oI-B��'|�%H��?(�����)k.�N��׀�=�O ��H*��<�!�S	�y�/�-R6%����}��De<�xgY� ���	�ʉ4�eE��Lj�\�0���,����]�ş,��D��#��z/ '30#���(��1������r��O ԧ�1s�:�OĿU��Э{�#�s�ZX��L'e��X���?[v�~��a��^P#�\�B���H�-^,.�	q4�<��f�V9F���L�V������BY)����-Q~�O^�XB��s��6�[��^L�Uv��]��ޏ�u�_��n��J��Rc6����h�<޹h���=��\��v���̈��aI8b��t�~#�^�_��A�,��~���]n<j��z��{���O�[b��Z�>$?O�ȃA� ̒���C�A3��%���m�(e��?�t'�&����:墟�ܸ�k�%�Pp��$�e�T�����k�*i�fN<;g#��{�s��Q Fw�'�y�)\S��F��|jX�|�N$�M�̀�?Sm�J�c«h�^,��Ri�9��؀T���Z�,��g��.Oذ�5�Sg��9	�ʇ�FAH���A�7�ڂ�[+̕�Ef2�B�"��eQ.r.Ѕ��^)M&�#B�>�ů.rY�l�����Ã��|���:�k2�ɴN>�hv��ZD���ZJ��#Z�LN���H� ����4v�Oj��X�=a�M��puK~P{,v��P��-�.gh��>2*����O�,�Y%UPa� h�� %��k.p�I�3!g$�%�����#�J�G�}�y�� ��&u!!^N�� �AU���������C��?�mə��zz�V\���d���9&
ߏa���On�r��Y�D�����D�v�4��ܔP��3\S)(�Iz;Z��| ��P��V`���*�+="��L޳�9<�$^2;P��-�r2��^��z��$��Y�"�ܸ�V�PWbs��YT��;����<��4����v���͐�8�3�K��kG��;����F):D�B0��B�ҩ�~in�N�����?L�n�r8E*"��ǚ.:I�{�wr)S�6��YEW��r�o��w����=�B��MB��Zn��š�avM�O�[�?�a3�
#*G��d��eB�>!����%��ʨ$9�ν�[���DU���^3�7�zs����n��`D���p\ �"w[�tf���!Im5��n�I��7����N	�R�Gk8�$���R��Y���s�ĉ��2GM�K�v��o�d/|�.I8hV7��e5%�2n�z뼗�
`{?�� �~PZޜ� �i	@BЗ�(x���*�$B�G����h���16�d�C�y����)e�M4�"j�O#19��	k1,���8�e/w1���_�ˈ��j���e���Y0G��74(:�躻x㤲�����Q��dtg�o܎���}.4�`{�a�}�`�]����-�A���%���U�M[���AO�#Kd8�5?EU��R��O�A��?�s���S��*R6G%xA�L_"i�:�>�=Q�!�P�t ���r>�����u�Z�D��C�<%��V�YmJ����[^��B䮓����$�6�p�*20咦�B�`�,T�G�*���'"I83Ywbl�}�J��]��?�o<,Q�Ԡ-�idϩA��*�Tu����m¥��ځ��}s�|����}a�Jq�K��$b�!���� c��8H�p�F��0�0<����7��m�?�3{o�n,P�i�������fn�jY�L��+���;Sx����7Y4]�"4�6��Ǡ��X!�
(C�0��w�FOX貭FM�T�%L:�����8��[q��d����Q?����pK�t�~^K���� k��ŦY� q5���{�t�a����r��ΟG�����G�1� �.|ě�s�x>o�ǿ� {��i�n˾y�ꦟ�;��U/�Vb1�����v��=�Q�K2�O]�(�3��	� y�����YY��\��F���5�����D�p�P�H���QY�Qu8O\zZOjt٨Č5�L�6
*��_i��}(���D%Q�Y<�#5p6��6�ǃy�ޠ��M�HVk��)���#�,�dI�����N��7U�p2����ŸԚX��6B�]Q��� ���{�*�o��}�x��o�T��ߏoQ4x�n�[�5{ oS#��V��&֚ز�65gtP�O�e�R����*��MX�d�y��{C�q���X�\�N���a$��$ɩ�a��6*A��8�n{�o ,��q���xH�2A�^�I�X����qE�\��PA(��N��p.eXaN���L�C}w���F���v�1NI����{����t�puH�k�}c�o��\�c�HǗ���� !���ߚ����Z�P&�Q� >"˛e�!�\
Ŷ#�_`�/A|�^�T�0�-� j��2+4P�K��PIeYJc��
���� +��%ȥ��&w��/��:�EP��P4xQ�����H@��Q<�C�/��V��th��2�V�8�;`�&���%Sw5���v߇�j_�Fgz�2�p?,���$�qAղ��nlVB�/(���`ֻ��`~7
�Iq*e/�y�gq�Nf�Ȁ-�&�W��`��gg��\�#��=�R�~��syg`<3��l���g�^�:�ߥ6XegֲԜ���Q5Int_+��<��I���GRAZ��<*
j a�Â +u|���B߮\x��̬�s�%�]�spw�W�|�ǵ6<�V������LJ?��dK@����faB�N?)����<��K��LÎ��~S��+}�G.$%������U�<?4�$���x�N��-��W�9�!�%�Xa��5BHS71�:���Ү�CIũ)�E-:�q����B+��z����`��(�7DV)k��8����X�j�{S��v�f� �d�^T�2�0�e����/L���\͓�0?�1�|�$�+S�Rz:$ёp�,qJNl�(pc{$VI�O���+R3�]�ɽWA�Z��5�=��&�L�oE��ڨ��V����$q�!��g,��'&8= H�KX!�Z�g�i l����#L K�1iN���wimk�f%\"&{F��"�*�b��K�c�����L�'������aM�\+���fR((�(Z�T[��]���yq!^���6���ki�BH���G�0�[�}� Q&�Bْ�4��
KNb=m�Ŋ9D��Iw�D?M��5����7�Q�߉?���N��C�^��E�4L�f�)�ك�	z4��xfЦX$x8�;_� ��
����Si��(S�?ʭ��yF1^K���E?����$`���\��ݶV��'I�#/��=��j ������:ke4Ġ`��M�54���ّ�+�n����-�o���.�iƮXL� 8&�[�*㐧�y���E'�9b�����C�{�q��S���US6mN�FP] i5��{���&�����6��/:�<�RK*�O/,
(�����c��.��in����\uΤ�C]�d��8R΋�Y���lfZj�z�EQm��y���v���z9��-~H�̆rѴv3������\��1
gt�l�H���Bd�CdJw�c��In�N��2�H��D&�.]�� �Q�#�/�M#�C���.��h���Z��~���KZO �:�  Q�v�.��E���Ga&Ty�ò:7"y�5mc���y:�dL���5Q�]߹n��Z.�n�}{�8�������d�4I�8�!�@Nl_��0����&
��eI�͉�N��̹��KAw�NEE�+-��`ζ1*w8�f��()��q���Jegh�ve���$�|a��v��3�@7�)�Y����O�]m@E/�QI����E{˹�XDT֞:M�v�MO��&��Myq`G��%�9��y�F7ɈL���p\z��26G��������Elc�K���lF�o�x�%$�p&34p����zO\4�_��R�zL�Xw���z���� ���q����ƳM*t|ņSv�7�Ąxdn��",��f�n����}�.��u�o]�W=�Ul�	97Bp��
��Du��J�Z�IcD��X T��%xRu�:�	E�
<��ѫ���Ξ�!�}ְX+%<�2����Dt���y��<0�PǇ�1�th���:1��G���]ǡ}�5F�������" @"$bx�6d{�~���׏���{�'���Q��"Z6�OZ�!|29�r_���H�%�ل��:��|�]�{�̌2�����L(� ��ΠX�~����$"�z�Fڟ0R>����)��������}�I�bndC��] )�	0{�o��C�7�� T8K���Uǜ^�bEޙx����t�{[�HM,'������OlO�~�;T�_��ݘ�"�;�(FT,:��M:X�2��/n�r �Tmd��U����4�3�Na��Q�2yh�¹�����}�)�n�j9��@��sHB��%�':ZjQ^�l9�?���Bj�ح��lq$�QY�O��O4\[��[�Y"�sW�|�N{4�:{EWy�oF�R�S}���K`�b/r�����T~M�x�{�2=�\�6W����8��χ��Sw�5
���H�N����`�� ��o��I���S�d�bg�������$�������l��UG3*��
��~�g�64����A@�_>B�[�œ�0����Æ�<׸�b���C�@���cøt���[�©�sx�Z��P��sF&Ԋ��y��K�V�-R�u���T]=�W|�.� �	_�4�kVCX��Tp
�5�N��{��z�<�aos�9{h�_/���b. �c�sA4d_�'�����A*��20�el�2Kp�����􍸂!PD,�I�}��$�����D.9�(%��>�*��J������B!w�u��x�_��<X�a�������������� ,=Y��	2ރ���0�>�׳���ǐ�|�f8�P� j�U�ќ_z�œ7i'�@�,�@9��LI�H�f$r��s���b�ѢL.�d^���[�=2�;�E#Щ_�+����S!�n!�+����tY��z�$a�+ݫ� ���D���C`��SJ�p���{�M��l3G�Z]���(V�>���30�]�!���F�������$���Dn����^|��ߑ�e>"7��g2��7;�/����宮
S�5��0�vO��79�u��g���ف#/����S��-'�i��Yi���2�Riõ���%U�?`S���s���J:�_���/o4��̱ qB�X��y�r@�����cz���1��~r�����.XR"��Uxs+xi?��D��B��+m˳Ɏe��!�#�~��:OT�~u���iwB��WChb�W��3���z��f�Ĕl�IT�� U߈��O�Zcf.�B�jF��L:�����"�'�h�1W2�Ȋ�m%�������e��uZ���!f�*O���:pn!S4�j�i���/s��%�8�����{��@D�!
N��7ӹXCZx��ߡ�V�HL�J�׾;����5G��F!!��\�	^(YZ�	Clt�
��C�M��vސ�NF8��Ѥ��;�\�q|#iw>�����^�̣'}�U�tVɤ���H���L|@�a.�%�}>�H")�f߮笒��t����mgJ團��*�㦶��Լ~���(�w�6�*E�'�G.�˟���<		I�0�e8P�gvU��O���`��A�'ޯ·�0y�ce9m�_,/�Јqk?TׅT�����:v�;�M&�C/�_]orbZ��Y��:>��uT�?�03����i	�1�A2ns7hä��>��T�����Ѿz,��^M��	g�i��e|����s�o�л�6�w��Mχ/�	�8�N��9�rd���5�y$���@�`���F'��6�v���,��OV��7��U��OY���CG��{�n������-�Ff��J$�ʯ�U	/���+��GzH�tתݡ���_�x)\�+0�a�A!�l%��)���`8����l�;V7�*��!'���64Z��74f	�{��,�J��RIgw�щ�]OΘ���(�'�9M@�A�f����s��[��9+�sǩf�~���sw画y�-Ri��!��z��n����!a�
nN��s��ė(5�K��"%i΍��6W5܊���,��8H]r&���@lF��.�M�:�)ɱ�FkjN��[�U���q61���G�)6�L����3����e�����f��6� Ȭ���M��ޗH-��]?ȔU���=������졥r��w9b�ĈR��#.������l���t*�$)j~Jɷ_d��`�_����@� �?-e8X]c���0?��{�����u��TԖ+: 4�}�X�r TBA��5Ո�!�57,�P��=�>-�h��/)��!�H��S�n�i�店@�&�2KG=�$61���� &*�|��nW�������Q{�i�An?`Q1�~PXe� @	Uk$'��r�j�S_3'���s�{����C��=�Gͨ7)�@@��9c
$��#5���|	&kR��P֪��hS�U��q�����$BA�x���ި��r�oa�nq�	�N^i8�|����,"�.e������N��dn�$ni��u'�gX�˪��`�+7����T�VVv���L�9�ߦ�5��O���{r�oN��#���C�#E�Ox�>� "���XH++�A��M�F2�P@�:�nh�~�)�r��תF(���Q+�F�� ���J$�B0��k$�S �z�379��1��;z����8���m�%��H�M����έj���:Ժ���vy�Ynۦ��RgWNz���]�j��	~ŋ��i%��\����(���d	�����Fr&0v�*}Ed6�Ӡ���$�#c������ٷ0�(�\�ԟ�ݾ�bj;�a5k6p���xh3�烒gח���H#�Jp�j�Y�� ���Y��u��qk�`�������z������^�u����5H���>�C�ȴ��7��јw��b���4�X��(�)	��B6#��6J��Z�IS��	p8���w����6;��7��SMM�:��=�fݵ���"l�\D�M6)'�blW��se.���՜���N亴�eŰdfM �:������54���T��0*w4�8屽�/
��UB�IwA���qk�؏AX�W`F��n%���`Z��?�嗴B-k�֗��4��G�:ϳ
C�*ó�R~�����0p��s7��tF��P5g�?>cu�\B��	��G��أ#Xx��A:�5��Z����Xۨ2�`X$-ACؿ�|���Co5lY�����m��V;�+������\K}�b�r��C#x#�ȅ�u�p"8@\��H��(9��C���I��zB��^�iI��9[>�	�L�\�2�O���^�#��X�K���XO�eV���9�u�H-��,?"�������|2�����e��m�-iTԜ��yHN���s���x������^B ~m5&G�����r&5ӿ0��ȡ���ҫN9���G�aZ����[T��a�/�Xi$ώ���ðD���4���W������-�9K� J��͈O�.�e�h��2f�8!��-�i\{t��zxִvo�*��5E���:�.�Yj|��8�N3��i-QɇS^�����y�0T�	���zQS�-<]�5F*C1o ��6X���&s��0�bً���aHo���y�Y�.���8�&��@�����R�gJ��DbA-�����q�j��#��������k\ze�Ss���s��^���D�7�4]�p3�p��T�[D��w�,BN����R5D�����W��".�"�����o
WF�\p��튝W4�t�{�RN&�C�$󨫚�vɾ��k�a濙������ԣ��
l�M���K������9�v��1�ԒHVp�����&�*�a���Q-�V�3n!w���C�d+��jS3�f����d���ŵ���_�b�H��Y�؞���M�����kī!�)��e��{CT���x��r�E �9�bA�vtb=o���
v��V}�7^���8�?}\vx�ы.d�@�Ü�kw.d�߀�����%�!��}��v�"ak5BD'����c}�i����h��=����@��?t��q��uZE>=5bbw8Wl�%��.u��V����E��|�k�N"���{�}�R���_+D֐�%)D��2����y����2�
�.}���5��zO7�Ɗ�d�`�ȱA2V+<��&$\�K��3xi4��?�$xvh��1�/Q��lw�������O�W8�E����YM�G	&��ON�^ڪ~��I���[��C���&,���`3(�}201ש!/�9rq�І�9s�A[�tmh�8^�Cm���
�{Ma[�^�d���[7���8��~Ue="���I-*(S~=d9�;/?%/��`�{�ӛF�9yk�=�E��]�<|L8�5�}�Aӎ!�~d7�L��u�K��G���%02k�H*|a�?y���}c=�/T"�<�	�-}�a�y��6y#Y��-��m{~����d.9���E8�=�pa�U����%	�����S�J��h.��U-pOS�Z�p���UMpoI�w��׆�3I��*u/���LD���w�Pΐ�x�^�^﨡����Nt?�5W �ق��Y��{�\���)�*Gb�P~7��y�B<�&�7�X_?�-���%&<�BɊM�Dw���w��Ά?��p��׬x�}�4]�[#�6�B���F�'�&�'�}G��>\�J�U��R�uw�@���X��?:Dـ�m���]jNK���`�;��4 �UQ�٨����a�Ö��߆�H�̊�9�Dsv�6����ȡ+أ�G�w��;i���9�2U�P9��t,�|��c���M�@Ϝ�S�k@�$�Isb��xBJ���}���D�v�8x�_�"�e���St�aOR��فD�\����W3�oK`|3F{�U���z<��IK�2ѭt�@ Z�B0pa%B�z�F�m�m~�YV�g'
G�S��N�#�+:S��Y���i�Hn;2���-N�ß1�DM�	�@HH�STd�Gw`�T������ġ���2��nؗc�^���u��M)i��^\d�D��>h��)���:u#��rL�P��-b����p&\U�[T`���U8R O1AY�e"g�Y�΋c6&��9�I��p�T��������_1�9���O��6+���o�*F�3����Y�~{T�2�贱u%�09��c�q`��,��!��G?	Ȥ6V��͍ŒRzÊΒ��zol{4�w-��"L�d���$6��j��'%]�:��w��@���:�1���_+KO9�A�*���_��[��0��J�I��)*t-;��W����Qfs�\S�w\#�{Gg���'פb5;�vy0�tG?��^�{*JmA6V�e:c|�D�Sְ����(5 ��N ���YR�T�z��.,,�V�bD��P����1�r�g[.ڙ~l���2z�����=�;ΐb�Jp�Y�d��pv̈́���m������w1�է��=@T,�,*	�� fVz"� ~-9TM�
Be�a���XO/Mw�(ii�������.T���ڍB�ǫ��،�΍>aB�`�Ƌ��|��p������9
�}�	%��3E<����i���)Ct*4�h1��LྱE����D��E����(��V�X]��a㉣f�
6;Z(@�/}H�?�a���c�թ�'] 	��Yy����F�T�+�F��� ����	#��b���@����,|羖KCF(�M�Hf���9����Hf2!s �u�����͇a�	��N�as͗��l�R�h�q˝v�a��3�"�{�,*�F�Y�G=e��է��y8G���@�*��\#��{�\�Q��<G	�����,���Ou�'��Y�ī�we��;�p��9���n�w�ɿ6�m��=��o�G�������-|#��ȳ)]cm!�v=���Z_I0�H*�SCM�ɿN7�����X����@���Z?�_{`e�O�� ��wN�U�'���C�XÙ�Rq�+��Z�UH�jػ��W*� �O1ֱ��-�,���{�v�IQ�1��ֱh�Y�.x�֓��˽V��>]�^I
��
�k	6A��[Ėv�^�Qێ����΂�ZDjX�,���^� �y=�"l�f�)���QQ��)�'gG�O8�}�>=}3Q'�]D��!��oy��)�Z��.���+U�������=:��;P$��R&c��NE�8��z[S�vb�U��S8��z�U�c[�"j�p���X��W������ڍ{}?����1E)H��J�u�iiotyC����řl��낀w	�!�$Lz��<K�Z�(cnUuYk�����h��.�S"��������w%�����~���y�ف����2T��H7�6���誄:T{�����tZ��SBq��
c.�-Gַ�կӇ����f�j&����_�L�e���T��������W}�B�w	��g�}{����#͡0��������a� B�<�M�t�)��b���T̆�/���Pq���@���}}Q	��9L��L��)]_���A�Y9(Uf4��{��N�'���e߉��,��*PS/�ݼ�|��*R�@(�Sm+��^�:�I!o+�;�"�b�7������US�����` �n�}?�p��ˉ�(���1�"�*��[%���I�B��F�� dm0�"4 �G�'0�нz_����W�&^�ˀ����?CJp>W�Sñ�zA�ͮF&C�_�οl�˵�1:3��5��<��EA*�����#P5�72o��TH�+*���|�<Z�����k��G�Kl������8�8��Ab~֭�`���M�3�5Q����L�/b��i>g��ejrK�A� �29�c�[8��;�'٢�����e�`.X'M�ϭF+����@s;l����G�'b��{gm?�<]v�&ܗ�M�6���C��<�S{9-luQW�֌:�w^-&װ��{��H�k�[q��O��)W�j�g�5��O<�F�&��{f��ԝ�aAd��l��}�ʻ�p"8�,N�&lC����xo�1w��k~tY9=��91�}]��RB W?f���X��b�L��y�~�i]�ht"4�y %��2��2[BL�IXͳ��`W���8}�J��C���5%p%IB,hf��lB���r����T�j���`M���*g$w��5Ġ�¦�&ZQX)���Ñ��i=���j(�rS��d�qyX���{�ʑ�L�j :�h{��Y�g��ಉ+���kz�^]�c�8���V+������
4�OE��᛫��3+Ā�ʘ��C��N�DI��a�I�#%��x�gN��p��������ͣ\hy9w4�Y��<�s����e���n�:MO�J�\J@�v��?�7��.���Gk�0�hoՅW���_(w�7[ ތ$�G��9$�m�#�O��ǭ�-=�=G}�hr�IP��_�d����*F��D:��إ�:c͘w�U�qx�"��b�b���mH2�W�F^N!�p�7O�N1��*O,~��D�a#$I�
�;�ҍ<f�W$�1M�-�ڄ���Babr�X�&��4������+�H�*5Ō��Mg��YL���i�shA��� ^�Z�5�L���^�����l�\5aK�g����w-�灯޼<��D�8F�ȴ &�V��� 7(�$8�if��'#��l
��O-�SAR���'�W�!!l٢��O�5u�D�_m��*����MYY]��S�����pD$�qH�=�C���\8ʂp5�d2��bk����]�E���~=�y�!#iOW���^�R@_3eB\�_�d��nP��hD.�,�)� �w�G*o��f�.�'�t�
"[\�*M�Ӳ=sMu����	�^@G��B{�u�*{��i�ʙ.�=:��ؘkwZ�AaG��8ݍo�c0'�%���5��%~?F���}�|�K��RmQ:h�!�EnHpf�~u��{�וGJ�)��Ȧc��I��F8ւ}Z%�l�0�1Zʑ�+�#d_-�4�����OR�$������{9A� �
@h��;�-p}�\�N�4m��bg"S��G94o6A�3���~�y+ j� f2��<k.�½D�ؼ5S�	�"���͈w?�E��V\�	S�����5�h�>m3V'����R��K\9�k�=*��>�`>��x�Y�-�B��f��((GW�k���:�D�	@ϱ������|��p��5D�$����$ߥ6SjX�D�p����������k��\W	1<��E�(�i@;R�aƏ��q����/�%~C-|.29��i|���U�ٺ��`B����1Yg���E����J��`m��&�]�"�(�1H�G7��@��lԖc`kY�?>G�:<�fJ��w��@{b����ߟ�#}��9d�E��Y2�i
�w]g��#�R���S���ְڳ��x�o����f���j���PG�l!8S�7�S�BR�L���z�B6Q�[�#�μ�?��9�Eb?U�I:ʅ��x�*,�5
�P���U�F��Wv<4���Ȣ(�B���ё��*2�0���"*p8��r��x��~��|1\;]	�����Xߗ��lj/:N/��B������d��2��S�<����D�,Pʲ9�#|�[����u�.��BE�ٷy����*]�{��[W�����?�YƤ�7Izd�}�jS�3�"%��<,�H|,] ��ᬇ}F�A��@��R=�G�p�}(��FD��O�ᵪ|F��-���1��6��2l��� h��_�Wr� 8��1W�.D��{^�qi��1z������4�<��3.�x���.��Nc�]�:�,��⢹��*<Ĕ���鑣���ԑ�x-��K3/�~��rM����o?
�a�`��}Rж��,�L���> AI�����E�)F^���x�y�1a췮C�I'_c�p�mvAh�v�����|Jq��X�'���v��k�ZA*S�F�����c���m�Qm�����?�����R�l^Ia��Fc�"�h8�E��#6Q�����#����Tl��ũ�d�sT�q�,S�\��L��,�y��^}�6�WF(��F���sFU�;������V@�����7���Fo�xœY����fAq%�a��/�T��0��(;j/V�*0�pO2�?��?�aY������"=a�M���-����K6��i�nۦM�v�:|�Sj�q2��699����)j�j�x��k��L�^o�S�>vo��x,IޔT`��_��9�\�ջw{�p��,��3r�U�!L����h�J)�J�J�Q����談�)B̚<��w2<�X��ی��E��H����T)���(7��rK����r K�,���)��5�(|�	@IҢ�-l��'��T��_̹�������ۈ���8|h�l�Bk,0��x \}���%�M6L�p.+�\�8�Oڟ۵eޢ�m9�%ӊ��|J�����e��P�QQد�9r���]
7j��tO*<=����\D�A��9<e�N�X�j�q���'1a�(�ʺ61��-ߨ���f(�wI�[�jԪ&|����jy5*\�0�D�+I�3��Xt���cm&�5q>�X���-��[.�O����G]�c��e0z#Qki��BYH�@���4�$���t��R-��c�jKb��c���&E��g�u
ޯ�����&M��'��,����[��VY�J.���?[��i�/��f�^9q\�f�Bn��<���	����\Si|܉�4����_��0�0:�����9�YS���-�!�c^���-�|0��*K9���J����P;���T[A��f\0�Yf�=�������B�)L��"'>i؈)�����8�6Mu��X�����~Č��9b�GJc�*���/���AS>���.BRj4d�#���P콱�Eg����7c�3'�3�d�z�a��H��P������,�a�?�a���y�1�`^������%����!q�^�w4N&�\׾�<�Y�<�
|ʝf�� VR�W��_6�@?_@/��K멋��K�ؠ�En�r:@���� ǌ�η�A<3�zB�����c�yS�B@4;r���/�Y��3+�v�~�H��������x�4�p|ővi�b��Bvw��N-�.ω�p?.<!?�z	"���zz��}q�Y��p#�@�Y�>�C�|�VC<HUU�(���+�OCŢȢ��	�{lֳc��0ja��A�@�Ѱz���"���uA�.�K;��R��A�*E�[�kP��l+qGb������ye��~x��PƬPz��ҁ�wxx��/�t��X�p\�[R���wf&|����y�4���{!��;Ն���#�a���L�x�����<��G=�ƴT��"	�P]6̈́K��V��uY��t��e�9�=�b`��V�����E~Y<=l�>��v��3e�Qn�T�@8�>] t�̷�(D�W&���
W�u�"D�?S�ޙ���+4����!��yV��I׫J\$�'�$���-j����/v����;�y���]� ��yZ�}|m��E,� ��[Yhh��"�&tis�x���ػ��S�k�	O�vkaQ�5�74ŵ��T��~��q�4퇪l���1��IO0pH�ru�A���cz�I�}9Д���Dy������#F�&��*U<$�wE�!�ϵ:W���|�`$��Ř�@2f�d�|r� �<��Q���њ �ɜ�O��"ϭп<An��#b*ck_`�d�%A�X	�@�	~9~E�$/��s��X�Jt�n�[/3Wۖ<l���o2�f��1����	��+�]�O�{����s��rP�ـ��F�L���X�V��
��.q��u�����0�e�K|���f.�cs�\��Ĵ���6|a�oLT�;eȁuŹ�u��$��mL���v.��k��$"�J�0�f�Q� �8�\��M4�5��~�h�Ӭ�&,@q�6|�V�p̣��褚fYWN
9�;֙=N�����Ә�����~���%;�m)��V'�_/T ���w5�����f��8թot��z��%)���#O��Qnt��A1�n�k����/�HO"��Y ����Aa{e��so�ږ�Q���f�#-��.t��wՆ�2��i�O4�L-�U�3Κy�ʉ��C� �Ω�˅�S+���}���uҨ=*G������G=%��2TsS��=�;Ip8�Ў5�`Mʫ���eפ���X� |���x9�Z�ؖ�� *�d�4�=�6Vu��$�VGK�6����(ҨuWO�Wg��Ђ��V�	�%n��3l�,6A�K5�5Ύ�%W?Z���Ґ��)"
y�2E��Գ����@����e�Op�dq(���`&������t���9��&������葻/�X΃�)���}+,�+��s���>*2��w'?-����E(��N����aӡ�,��~�2A�+X�dn&�����GV��~���t�.���&��e;�y8z��1�9��*�(f�A(�:4����?��t2W��_�ǘ����.<2&������'a�E���-�Ta�`�Wmn6�=�"d�������c�;�u���:|@�;������Uz	�&6}nΑ]�Z��'��T�����P�qO�����J	�i�>�b�&�6+7g�$j�JJH����|a�ˎ�HHK�-5��羁������bn�}�y��:�^�{��-zs��
UHk�KbZcX*�����P�G@���Dؤ�.�M��۶�4�\���oT�p"�h?!ݝ����WUfK6�ѭ�|�g���MZ��N��^��H�f��ny�e\4þv{����WF ����vn>��M�n{!�U�-����Ys!V�yt"p�r�l`q�_��}��l��OWA�.�<���ei�#>���A�W��Y�y����3�x�#�:�<�O��A?5�p��xٶ.o�1E����C'�(_h��)�\=�����Y^j[�G3�tX�N{P��׃�A��B��υC�PE�G�b�RfӴ�0�ɭ;s �5�9Rlb����������e?>i#������L��N��O��$a�^�0��ĵ��L,~
�̵�Z�5��$��i�GR���?�d�k�4v΂��_��X�\{��D�W)#p��kMX�y0*ήz>ze�} ֿ�0Z�"�od;���y�В�{N�_oD ��"�杖}��T,��+�B /�HZ�~�S�� �nN&��B�#�T����_�C�1�]�-{\��z���vxK.�f���PN/������x���]�T����,1��G5�e�?ܜ{�.@��!�
�ٻ���O@G|cj�U�LiJ�ɍ��8�<|�ٓx��#
�)�h[ɋ�gQg�a�����
���0�Ն���D�\Ϫ�@Ӽ

n� �ƾ�*ϯ���X �|t,a!���?��x�W�;�+�m_��6� e�5�Ƅ_�N Y̘�|��N��|���Yޔ0t"7��f�L2{��c�_������,��9x;H�%��Q+"���i�"��N]��!� t5�I��IӴ	�L6?f>�5u?�&O�k�',��Sʿ|Xo:���7�����"���0�B�����+�7A�vp��ݳ��,cF��}eY5&�z]lv�X�gxw��)j��ny_����`��.���s��)|�0n�ȯy���*��PQ�ԏB6$�2�6[�Ax�n�bf ���Z)�h�ݩ���W��:'��v���iX�E�%UӦ���XΛ��͸�T�{�n�����.^M��$�=Ԑ�~��/�p5e$���w7b<�4d���K��M��UA�LWyl�A��U3E�9i�J��Kv�X|��I��T���z��c)��]��%wW���߹�����h`���Ȁ��"VgH��ND!�y�I*/����΃���M���e�l0���FJD:DX �q~�v�W��_�]+f���	��R�i���*��p��u���.M/����'���w�#?m��R���J`�7�n��LV3{�xz�\�'�vL�.Y� X�"4�s��?�ǒ���0����(;���;���x�����	�+.U�{V�kg���+�0=NVe|*�ZBR�'Cu����	��Wf�埻-z��1_xd�n�屇5 ۜ�_��͉�NL9M�i���Z$��LvY2O�ptGX�"��uw�R\���l�2E��m�إ��&�|ha8I���Y�!kS ���`�6I�����Hz���}���c 1F�x�F;��w���־�p�o� ɋ�D?�T)�q��Ō���`��ʽ5�ʓs�x�@�����Ρ&W�2~}�퐛Ա>�hr�`�m�8g��������>V+ǹ��"�	��`���u���nS�k�;�[����r59�