��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	�����:o�R@9����7�Y���dC�%�&���2=ڂ�"�k'w��W�����ǭ��,��y �'����Y���ewY�L,�wNfAXg<J������ ��¥k%|{�����cO�wWi_���<�'�Xb�����}����d�d�veэ����	�JB%Z}�n�+�l�M��"�`�aZ����c~
��O�J�/X�Y�Ȇ�ob���ۈ?�]T>��\$N��Y=�|t�z��h��1������whA�d,T����4�l|f�z�ѡ�4�~v�Z⭕}!��E��9�+,�$�����є��q]���k��B.c�dx��(�ń|!B�Qm�J�p�Ԍ�z��H�r;	b3{}X1�����������w�ւF���+��w� �嵔�)[�jju��#B�"�,��Ӽ�4I]3s�̤V��������rWh��!�n��g�Mq!)[U�y�N��~s�m�f~�D��{��NWN�|��d�����8�;�'�����g
��q6�4��V�����/���K��X"�8�ے��W�A1�}],x��s��zOc��wQ*(N��x/D�!��/',:������D�(M�ύف�Sc�m�Sf��iW?q�1�ã�Sg4��A���T�fs\=;wL�]I�ON�܈�V���֯���d����bC�F1����U5x�{eU���-<ہ�Gm��䋷�ـ�L�̶'�g�e�$��:N�~���l�5ke���Ѵ��S7
�h=Ko�S8P�z�-Ml�F]�?�$~�2�n��}K��?..s�b�b���RG�"[�v���nք@+	��1�������\fc�4V7���7{N���U�����zSr���՗��6e���%n2� �=]�t�ky�]��,��3�Y	RY�F�������\����X�MO�S�F�!U�D����=�G"�܇�ȓ�Z>��������{��hhW�ͪ�H�(��eb�v�?�����ԍ0����6ANz��q�m��_9j)q����p��,��̂[%�P���D3����f'�c)���GL�)�v9�,'`�� ��� t�s�<����M�)��q�خ�C]�dO`p���p��'͵�����7k����8eÃ�lF�*� ��AP~��U��=�-G`��L*E�)���[�
�N"%�������,�c\4[Dg�G��V��<UG%D�xn&4j|A8U��w��?�v�b���y�Ƕ$W��g��u�c����ʋ�������j�a$���\�������vS�||UBE\,]hFȄ�����%�$)t��%�+wqt�0�W�IG�Z-h'x�|y�%ي��?&>�ҿ[$�5�Gլ�L�M�Q&7���5�L��z�	b���E�?�ߩ�c�7b�TP����4+��Ka�Eх~���v�M�~���8V���Î!�"���)4��ϻp � n�ب��9/w���"w�d��V��E+��oο�)��s
����Tn'���Ɯ�i\�9_�
�����E����ู|�8#n�5���z���Z
Sp���lı�u��B�p����;W��J%8��r|����+���d��?@F��K�ֽD��[7�^���7g4����JU�Y�?�l��OBA���/���G��S�5#��9V^<na�](����D�
3>�㗈��%���[�X�}���;���'T_��l�*�a��f�rX����ܵCj"ȧ��W&_j�����O�eT�(n�80�\&7�WB�9\E����M��)���2a�Ї#��kI]��Tt��8"��K��x�tӡ�L#���W�j*ѕe�WV,�3Oج)�)Y�qU���Xs	M�b�G�L67�M`T��H11�!�1�,���SY��1�]�
��j�2��X�\8��ɷ%ϻϘ�{�=��>&?��I�C�΍�0�K�z.�_G���=K(��;R>�w�I��"%�/K��%!]�SH:���=�{�fF��nu��'�6�H��jŉ{/�>����4w�H1�:ڴ�K �'�"P�Al��a�ڶ�>��ԑ˕�@g�K�M|�q;�� F���Fc(���2 �4���� �{�'�_�*�ys��g�˟3�z�*3�pQ�����ʄ܅5�\b܂֤�Y���v��ݚ߾f���;����?)b�]�ʙ�����=��)۽������>�L�K�RԶF�	���tVV��L9�{:$yk�L���[�1�b�luqɗسlGv�	��ˇ����c7��+���?��8֮��yx+$�� �[�i`N
WS�:��ɉk�����%`1l%��/h�BQw�<��H�/'Ӻ?2�?c�D� �l&҆���eP�<"tH��*+O�����D9��f����X���>�>u7�0SQ����&�P_��}�\�L���T�+��|uei?\�H�J�j>ĸG��Z%٘_���c��0ݧ;)�3�e�ݑCܑ�ĴZ�}dL������=n��{
�p~�۔�?��E�D޼_���֍2�����6�AL��B�O����;�F�.��Sl���}��B�x߲�N.��D����
�3�zYf����bt-��8O�v(?��Tp����0�	��k�n� >�n�ou8��o�ghyQ[˵��/�au���p��F)Y#-�&��t�N&����OV���{�?m!i;�y��T1��GH��V��%�	�����@Ɂ'Q�0�L^{c ��=)��k�!��©.:�3��:x��F,�O�sm�2 �5x5�s�lʍme�4����mi�B��}�Љ�� �����|������ �RdB�ں���b��+�{��7���'��ē��IC��A1y�K!HF��h�F7��t�F<cY�\���A%�D�7j�������#gs����ze�Q���t8�RT:7)�Ȑ=�b�����0.C��f��rY���d%Y��\\X�&s��?k�E2�"���w,��Ϩ�~a�O�kiL�`�7�`�����L�s�Z��y)U�C�AljA��ꋻ���P�?��J�,�5R~�a�/>�r��G8��ϡ����V���1�@V�#,�P��Q���@�?����΢�ZBSO��hW���� ��<�<�8¯�%e2h����y��~�4���UE�ui_�8r?	�����y��@�T�5�h�.RL�:�dp�`��J	|'Z�v[q�Y�9j�(v#��ƈ�Vw;U)�'���~kR�W��?4*L�b��B<	a�zP�hQ*s����x�Q5��輎�2qa�+�c0��#j&ͱ�ХL����\|�,�/�?�/��g�Cr\��� ���_({��VD�ɦ$��|얽���͙�+�(������G5֚�ԁ��n��1
M��/׆��1O��f�H
-4#�6���ʷ/0�w�H?հ����H#��:��ʟ�-��t"�0N) ��U#�j�i OC��;�9!+�PD#���&tu���7�\��U��5#�� v\�Ňs��_��Ľ��r"kST���/S��Ztiҧ�<T�O5y ) ��W�$؁?8���M�� ��<ύ.���`W�������0U̬_�.�Y���Iv:D�QP�X��䜆���(ۂ�4N��Ɂ�9���a�����i7%~�ͪ�)/�}��Jى�ߖ*��\4��X�(������@k���ř��h��d�j�^�G�I�S[w��cs?�"��6;�@g�W��D$0?��^ʨ� �T2�|�t(�������*���Ҙ�WqQ&>nE�MṀ��9��{~���r��l�z:e*�H���~��a휨�}�_��^~mJ$��eUw,��τr0���Z�$�B��]�#�*z���h�=ȕ%�8� 7J�C�CB��M��9�QO;z����(A��Ŋ<m�z;�U�4���܃[�$�:��%�#c�_A.��fH΂��G���J����@'��޵�r�-�Ϯ��';�gkh�'*dJe=���Y�ș-\#V$'���j��Ȃs;��[g���c%0~GeË\�L�M�K�}K,��K� ����g�%�����en<��Zc��
�
�+7�)�A,On�l���r+M���G��;�b��7vl�	$��*B=@_m�������s/L֓�5�?Š��G�#��Z�P*+hb=Me���e,M^�5�\s��,�/ �mU�#C77g��Y�BM�O˔�����5�״PJ պ]{d�;��29��rJҔ�kfd(N�iH�t˩ߺTq�[�\5@�Vx�!�f0�8����E��أ�M�]њMV㉦~�� Ϸ��ZhiC
�^��t~��~\��i	�<|���	���-���{{�"�Ś��Ͱ&մ���@�۝�${��OǓ\�:��%��בd�}�W����Wh~���t�;��z��C��AߜYpO�V���o��ck�?�O8a���֓��M�ւoH�4��y�&7��Px��Ycܒ�ȴ4�2ђ����\��«�2M|�*�����lI��.]��&�c7���5wK��5N��<(�NE+O�d�l�&Cw�ӕ��y����~��d|�p���
9���� ���d^��?h�kn&"�ʎM�M�M<�&
��v���}�Cj��$�9�9:w��ّ�D|��f����iF�6r|%reS	�4v ��w�4_E����� ��ūn	�;�n/8F}��d�(�"����3��#ac'�cX�ۻ g#�OC␯��|����N�g��҄!�B$Zlyl ����3��m1�0	������.�սt�t�A1��I��}�����ܙI��?u]UoT���(�����dt4~n��G��x�{c$ڤ�`3�&��j��m��3g��L�ݶÕ*��Nyz�=�s4g��TfY������т{2�^�m���_3��nN����@ �.�!�+L�L�O�O����9��V
<OU4�5�#�{C��]�9�щ��-��M.�� {�0��EӶU��Ғi�(�c��QA���'H<y��6���C�ZP� �d��Չ}l��W��4��Řֽ������;�НżP׃P]�8��Ԡw��G�[)�Dj3�L���Ak4�|��*������$�i���<Q��׫�%���H"F��Y E�=�o}�>9-%�J^��D�GP��K�?WZ�1�/Cԁ�ڛ;{$m��j����ָN�yG
H?�����k:�͘՗n]>p]���ǜO]�Ý���7KIm�4�O�GZ]J����KүmŽ�N1YB)2�W�#3����@����3��X��1&y˸�I��W���)�j� �27(w��/�� +�]H���EY8 K�NP�f/��0������LA��zuw��q<NzN/�=V��W���J���?�V��/e$��d���T��;��u���$��������b�ų��B��� p@P-b���g�4�F2N�Ao�@OA"p_�X���#��b��K����������6s!�d,M�e��h��	ߩ*��D�	R<b��1I�Еn����u�{��������*�4<},<���e$ ���,&Smh�~PIV3���e��:�m���öL�Ų�2Z��	|@����3�(��&﬉�~.0tw!!w���Ώa�j����v+��g�3����+P����k9pثx���8TU��ÃQow��&�jп��� �BC����3������]2��Pi��/����Ow~|�I@fS��-��kۗ%��v�՝������Ձ���{5#��FЧv�տ�;�Ե/	����'�g� š̆�cR�|�[��.��0��v��oE+�B��:a���b�4D3������)�D?E�0���.�sw?m�t�-)ƶ5 �Cd�*���D�R�� �FOz�ɢ�l�	�;���fW�l�K�;�����d\`e�ٔۼfsMX�h����Ԝn!��"&+�OF��a ���wb�t���I	���-��f�[}���)���L����O���{��Z&킼�de,|F�	@m>�������ه�m���2*�{p����B9g_�\�C�x{��?k�Ss�%息�c�R+�@�<�|��"Hgii/�;���i�+��;� >Ft}��>� 8#R� ��e}� �A�)��R*��9�?j��E���v�F�x,��BF����J�/���E�>�ޚ�r��}��w�.��Z��\��bҳ��������K�Bfv���"mb4�ʽҽ�����R��UX��m���-�c!�/�� �b/�@��.�_�qC+�$r�5��_ѧ%�_�A�"�B��?�O�,��r�/�-�x��(�|�^�4.ao� �6�뚊�c���V��0�C%9זp�݁�H����(��7ג�	z�W�@)���i0����v�q�7�s?�2��x��M��V+;@MAK�Jh�o�$��Ԇjb�)�e= �͟ �hz�@��j�H��`D�@X)@C�耕�@���~��C~��P���=z��+#�y���u��Xl���w�8QA��$���&ZT��V�ӥ�]����0���@׈��?��}�T�kJ3_i�qp\.�ʓUߦ����X�ψ�:Kх�#[�|�w��]/�f�.��Lk��e�׉�����	�-�,S�U���>�.�4q��((RAo)^�����Ozēf�#wg�;AR�4-�4=!���A!<�(� (����|6�`�sŅ�J�8��[��l��DXQhأT)_$�{���v��Qһ��qb�R��Y�, j
�8���	ȏEB�a2<��%��s-�z��Fd�_���[S��K{����7�Sv;"����U��a��;|����Z��|V�KaQ0vQ�����8	�)�����|[�H
��<�nC���U���2��cq��P�Qp�:�`hV������2�Sd�xqKԲu�40;��fJS������:&/�����L>� �X:�q���9<y��m�A�4���Z����7U��D�"���Z9׺|2���m�+R��1���VZ�Vw���|�=.@�1��V��Ԟj��x�5��2rM 	^rl0Ї��ͮ
K�� ?��!�Ɍ�"g7s�%k� 4�Y���~�ir6��(o�=mc7��=t�$�i�;_�r�ݮ5��&ڒ/)���T�X}�O��Q�|��x���/�:��/� P�����ںP6NN������4��lM!��i�;V7�v�ʦ���"4�L�~�0>�Y��<*�/0gM{�x�+k��xT6G�dY�s���+�*��v��k�1�+H�8�t�'_�GZ��oI��з���]��[O�����a��q!-�0j6v�#��vPd�|
h��@�&�x��5T?�n�i�>=���@_�2�a�ǀgN@�6�e���l�
�@x��w�;ݷ&xy��MQ�H2AfK�~�N+��r��i��cW4m��	5�W�U��-�;5Q�BO'��� )�7�|	yV�����7
E�,i]�N�Џ��=�7?v�=�l6���kc� ��j ��0��~8����+(�03\0Aj摉�;J���!��7rZ�㭷��GЎK	Ӄ��^n��r¬�����}}zjb�>5�-��{Լ`��Y)�Bѩ葎���Ap�v��I�"�ڭKF�K�����f�G�G�g��ͽX�\�O�����3U�G�7��.��s��O�N����0,
y��J�l����@���v>:0�1u
~h���>�"�C�"���&�~E����/�;%�K�tqP�B���������5�!�`-� ⿸Y"�y���jC.��K��d�9jҿ�xsS�$�k�E�(_�����ˇf%A~qP�P�~��R"/��I�ׂ��!�)��F2����MP�������p�zN���w��/�/-�D�h��ZNM�N���0�� �K�	C{m�4ޔN��U:�������lW,���m���"�iF�`�������q5�m�B)_/
��v*|��'�x�8e����]F�T��Fbi�k�`�K�,�S��,�g��:�$"�}V��c\�8��V����*+O<E�$~i��:3hO	��S�?����}쬛+s����p��9(��#�8����o7�����E0g�`Z��%���s�ϞO�|�4���ږ��,��Jxv��y��gܗ��C�)��#��؅������:�ef�OW+���+nJ�e�6y�0T����|�ԋ��������KZVQ!1��@�/�,�[G��#�iEë�T��\)�T�/"fT�7s�[&��Gy�Yс��^<<@�T�Ak��]�aS&��Y^+ k%b�i���UI� ȓ���7�3�?{e�N;B"�<�_XF��h�t�mn�����5��e+�O�wz��w/���P�i�,7�#&�g�I�	��Ʋ�|��? A���oؼp���Ml�b�sڎ��$U�9�ԉ玷4��zM��g�]Kfy[�G�u"�T�c�R���D�ݫs���Ѱ������J06L\�����Ԅ��mR9�;3����m	!p�{^]�gޛ��nR����#cq7�YK|�NfT�g��%�*�z�d~_}�3#���"I�/a�4��5c�\4�Q�[�M��p��z5d�9�6�d[p�=,�J����Z���In�bTp�ҡ�����!�H�ʘ����36���3Uj`�b���ty�»�}��BPiP�|�ģ��
�a֨��h9�	�l�|�� �ӚN�c�&ͱ'���>{��twoZ��ǚ	�r[��4Z� Q� ,�����b���ttO�^L��e��K��,K?�S�[�겮��ͨ�o��궈5 ���~C��ȷ����7y!�� ��Y�Ҟ)8{A�sE��G"��	��K,M���c�X �`�v�Y�a���m�W.|��Z8[%��y�X͢�$���邻�e�?�(9"6�`p�zEQ�z�����C!OmS�y����q��]�M���xhm8�Pp�&g�6��!���I��4���[5  ��Ðbj{�7�1[�����'�V���*񍐆q��h2�pW���'T���2��I�r�(�#��a��ܾ����6���������P0�+,79�&΢@Z�\`v���Y�td�(}����h��G���,	��f=7	��?s�JV��[�/~�H�~��"��z�;lӉ/GۙXZɒt�E���X4��f���!�ҩfTɔ5��,�-)��h"�D��uW�x�*`9K�x+k(j����e�	
��lY�:�s��^xH"��P6Z�b<��֤�a1
,�bLR_��{���D�q�=��|�a&��7nH���t8�9h��'������I�P%
W�2%:Oˌ|����%z�"<8���6Wy$�c���*Jj�
��ڱ��{�b�9>��kWK(f�@��c�'������³�E�ⶽ	�aF��]��E�e���v�{�P�E���aG�GLg�R/y \ݽ *a���}�=����:�h3�
͌̉� q��:P���$P QD��"(?XÙ�Z�*�X]�H�$-�?�����
�8*�JL�C����	����`O^C��"���_�V��{9������LF��K�_������-��X��H�"0s0��L�#5��ؗ9�6��e�9�]y���-������N[ׇ֟���m��|_�ٱ,��{��N$��D7���%��}ݟ
���.\�~ͨ��r��[�2��b�9�+ҍ�%��Nu��> *�|z����P�5Jz��K�3��;R����sq�j�?j�|��?#��Dhh�EFn+]�s���H� e�j�G}�1��Nm	�;�tU!v�3R�Su��<K�]|�.>HZ��|ː/�kzpAte��78�i��~��G��ۦ�U�.i�2���{�~� �{g�C�GnÂy���)��Ƹʼ������$1�LP/��w/�4�����W��|��mwG�ʫ�!&��\���*�������rRpB���7��ʩ��*�Gͽ.�v�o�6x��H���V;i���|�:�BP�I>,�v�ւ[S�ڎ�
�� �\��h��fn�S�SK+�?�N�� �G3�*k�+��'[gN��4�q���N�x�������e��o�9)1`͢xB�sζ��ޓǀ�,��[��15n�qc1�����\��nm��\o���n�.Ɏ�&��b6z��Y�Yb����J� ��"�Z�e�̺bG���%���L��!R�>��ߢ#��C�����v��ਥ�bz!�Y{���oEn[���
S}JGp����]ܯ�r@ ��	��x6�� ��>��	��Aj�g{d
i�O4>�P�ه���0?���/���Y����|�:�s�C]0#
XJ�y�L���[�|$U�'T��n��W^d[$FC�ј����I<y!ǂ��Ӎ����X�A˄����rB�(�D�sݮ_�P��F�10ۛ�7>�6(��T˔}:?iJvX���*�k2���Ȫ���m`���l8g"��Z�����8�yl��Hv�<*�U?r��ڋZ���ڹ$�M&�n*w�G:`��:
w��%!(Wk}n�y�t����Ŗ��K�ۢ�����>���BR���e\�K�-F�Z���^a�/qEUmd���� P�g�H�'���p��eĥ�Z:aL�U���)��$ ����s���˚�7��gRp0j`�O3d�/���$F�SCo� �a�ٛ�p�{U~Sd��|,�3$�b�sP�E9����C���7�n���ͤ��?Nǥ�E��'yW$>�+�R;@8SN���M}�>�,	�.�~�Ϭ��|zSd��e0�_V˼�«��.vI/+����&�o7�a¥�[�ɨ�R��3�|�΍rg�WE�	(��b=~A
�:�_٫͗�0��+2+1�Zo�C��]�ׁf��H**rW�e:&�G�T^�c���3bySU��Y���3i��ǚˊ.�]�ߥ��h�֌D���Qy��s��6Ir����)�V��x���lavDr؏TFy3!��n�FfH��@I�J��@��a�2��&L�"��G���Kg�^��;_Y�ЕWg�s���d����	�{��e�E�����Ǽ}^���r~��VS�i�:чf�\��'���O�A��+]\ >����w�����\���XP�M-Af��Z*�Q��2C��^��`�s�7m�ϱb�����N�R���4Q6�M���-��#��]�4����h�-��~�6Έ.�Y9S,��^J����'�T'	���.��!A8��뙨Kܮ������w�=���ɅR� �}$M�s`��Y1[.[�?��ѹK��d7���}�3���H�s��)�_;γ�i@2�ź<��[o~U��wG^���E��M�x��;��M�j~����ռk�H��{�����q������Ԑ��1Ě�pj�:pXER�	X�����5*N\[\��݀<I��Y�r!�2aE�BEi'3(��[�(���2O=��d �u��l������.�"�d-ΐ+c)y�&���=��칉�Wg�J5��C�o��nǨagUnesw����Y~��<\�,,�h|�)�@(kw=-�rՑkW7��U�U�����5�e�w���6�p�Uw�x�~��c��ݴ�T��=n��)1m��Yu�4uq�y��J��N�Ӎ^ҵy�����9�1�
�@��K�&m���(R!n�ر����������e��׸'y��x��ch,�m�i,f���`���у$�����{[Kzv~���R� a<+q[̋����[��Wz���8���1m�{'�����WT����Uߣ�y��t�	wsr�.Ml���aH�=b��>(XhC��^�5�^	֯R��������8x��^�,��|���d8<=����+.�J�^%���I�k�`;���n��5|�Ul�՜V�+!��Wr���賫ӈpUKU0�^�(�G���/��O|/Qr��qT/.Խg9-��=ft�3D�7T1
}E�w��#t�7)9:i*>����u�1eb��b�#��Ql�{���&�`�8�C}��]��I7�kᄔ4�)�2
�[hP`^�����o�xÀ,���sT_�Q \=!���v�`�N5/�U�Վ9��e*@�3��@)r���$�R\�8|���Qzs�[�*�r��4&��Ch�p#����5k��f��_(��@�u�����d?g &w�vJ��l�Ew2Զ�_=�JM�F�#o(���WbJ>���)����Qkh�O�A�]dV���"m�̨�)� ޿�R����7��~��L���ܟG�&hߌF����:�����+F>oɏA�%�����rr����Cu�!�n8�w�E�B���	ˬ�*S[W}g�6�_��&W���@1�Ą	��Jba'�$�s&�҅-�� �|ؑۆO���\�f�ׁ�\G����?k>~y����D"S*�Om����:(���z\$����<.�Η+��U�����C*�ee#�!�V�%@�Fam���T�U��?������u��Ɍ��.���Z��eH�%ۦ4�5x��@H0!��B�e��Ǐ�$Uj[�:4��0���G�����{^;q����qy�]H�����Fi�Y���{��e�,�㽌,��JI��&R�G܃Z:�!7KK����s��?{��[P��˵�m�Yԣ�Bn��C�g`'L\�!��`uK�;�����
�ޛ`C��R��퓊��7���N	w;p�iT�˙wo�\��J��п� \��9D����N҃��О�1�����̤� ��R��E���Rd�
h�����
ɺ�XϬ�R��g�)YS|�� ��]5�*w�؀Ǯ��P\�,�(�E��?���{�0����@kK; �Ʀ�m����#����v�o�@�L.䩡ͷ�R|z�"r�D�M��P��dR\�sԃ�	��Q��0�EDX#f0'�_���q��*�D�+�Z� ���M��ܑ����g&���{�鋟���syaR�MD��<�:Dd�����r��*|�K�1�zP�eJ��ݞ��\���$���Ro@ߛ��%iRƾ/�#�),\C;�� l�{,!��Ϙ�\c!�0ԭ�A�'VB�{�`M����T~�s;n��В܈��rt�<V�`�_� ����-�έ�$a|���c��+|̙�g&�&Q��6	ky'�����*c����tbaf��@�uH����Ue��_̀�B���S��g�����J��Wi���=���5�gm�ꉑ ����|Bt	.�f�	:��#�W%��_�L2	Pqt���`�����I�����x��0���j�3���ryl��
a.�^pN(1E��'I K��e�E��a?�l���b�{��LU��o2O������E�]����]������s����Kng����1,���!z�6ඈ�n�h{K��nڥq\�x�)y�cu\��i��Xf���A������_��K�f�/܄�����=�h,#S��r8iTw�x/1_yFF���V9ftmk�t����H�����ljF������_���sf,��y��ԕ��%j��=L�<�b�
N��s1���u����C���7���i$�I��j_9?���W´�Z��vzzá��"����M#����aI%���[�__N ��g\>��N�@Fr��6z�v�Qߠ��5�E ���0�J7N-�Pa�a�����<�-WJ�S�3]����ż|�F�qtI9	�gt��t�O�6������.'��!��b�V �u3y߲�!�t�P����G|�2��D����\��橿wb��g)E�9ǵ�}P�C�f[�~ ���j���w0G��n�[*U����3D�>�%���d���D@���Q���l��ujq�s��=��0m�`�=1&Ϝ� �L�l��ܥ9���=� �V�M�GuOH@Wr`�7r�1ٝ���%p�ࣇ1�@�^�Zv�'/q�M�q��OΫ�(NF�J؀9��B��fB]���u��E�6�S��S�R5=E"h�B^�� ���P0i��K��xJ%�m�ak���g�n^����A���l�/Rlň�b!�u�$�nڂ�).]��-^�Ph���o'����&�����$&ܩ������ج�ͧ��n��K>��.�Tܑ�߂�^e7��ߘF�75+@���@������^d^JQ�e�l�k��J�d�f�ɑé�[�<�;��ei�h2x��J
G�4yʅ�7��+���j��ϴ�c_>�k�?��ϫ�bA�+�����n�ξ��^f�P����x�*�@$��9+}A��3A�)u��5�
n4ӗE�di�F�\Ӥ�������X�8�Lj~0ܤ�Kܝe(E�ØX�t/�.�m�P��Z)k7#�N>�Z)=�$�;!��g?2WJPE��G�����`��L@?����uAw6`��w�1}m��9���=h�#�&tA���D���\�yo
�$�Q�`����)�@����q���`3#�N]�Gc�e��T���r���G�B&�Gw�_0yb�z~��J��jq}��o�W�q��~���x~�M�]!�+HO��ZZMp{<�H���@R�H���qt�V�ώn�����`4#��>5��k������6Y�Ģ]ύ.��}�@��4u����}t!��Y�q�:0B����>�+�����c��~�Z~M�����ط��}:ZC*U�t�=`&�W;�E���/F;k9o�w\���@dI$�P�VU\�d��l�}�pG�S��"$���v�Z�cp���T�q��M֬�x�	x`A�-��%��`$Y≠��n��eY���r�Lf)��u�Z�c>��g�DR��	�Q��w�^5�Vy���3����Ӿ�C	��օ�v������my��bo��ۺ���!d ����0I�m��5}�ه]�������^��&Q�Y�=���X4a��;�kC	/Sq�;%�i�D���m�D'�a�,m�3��ˌGPw��.���k��p�ES~J�˼�ƴd��C�_��TO-��}\C;F�c:CҶ0l�[V���RBX��Ԓw$�{�8�K����5�<�ƿ�!�Fc֖9�]��H�)(���;�������L9�	
:��2.�a���:���Y��A"��6�?]2�=�p��O6-��.v'��	�q��ĮJwPʹZR��sI66ˢ�rY���|�t1�8p����5涓�I�!J0��X��	0B���K�G�m����^5Qr�,,�¸/��γ���C-�H����죎�Mm��Y�m{J��wc���bE��k�K/��]6|�#� ��v`<ۘ���ϙ r�K�F���nבYO5��
"dN�~��1����V+�8�t�Ď�~�cqqh%�=����o(K/d�%��@�x^W/�(V0�t�}��!�sA0wmU�z6<Mڹ@r]Q���p��i
#(�y���3�Z�� G|>��&ئ�ʩ��/�5m��\Ө���B�Oe��=���Ouiv��|�1Ȃ<�Kz�m������OŚe+�h>C�Ō��|�l�9�(Z��s��@=�����*��_���(zt����E�����r��F���r�i��Gr���-�ui�OQe�ˉ����߀�S�T�~&�d��[$�[�6X�o��de�������S������M+�o����	αf�j�[�\T�Cn���9�'?�>t��|�[Y���`��]��a]�L�S�T��+��8����w�~2~��Z�\����o- )�����{��-�CM���9�Q��q\� �8	y��|B�$��Qxtj�Ķ3���6S�F�ߗJl��U��K�.Tn3GZ������h���ѻ�t6zwHڲ"�(A��7f?����7���1A�j��i���و������Θ����>ݫ�وN��tYU����������%����&��9i��$�(��:X�
���AWc���p�?%u�2��we4��߽S��`��F�\P�f�L]�Xы@�9��	�*X�9D���Dm(3;IxxU�f��B}f>����ݸR l��
�s��ӆ�孲�@������"u���_x#݉.�a̹���)�����d�LdzZ�Ђd��g�.�hQ�F�1�VnEB�?u�>�����qs���r���Ɋy�g�y<קAP�(�=�<��O��@3@�%��b���K��S�����t_F�PC5Ώ~�cU)ف���|l�鰙G�5�4%ߊ%YS��ぱ��(?	�B����R����h�k9ٞy�3v�Y���{���Ƀy�����4�I����y�'��Wb�|��84�h ���f8jL��z�~���y\?�b�[�e$��"z���	� �D����9ZqA &mƏ��[9�2��7=ȏi��d�]�Z������s��a�$�Oa'�6^�~9=m�����$��FF��(�����h���T����Q�6ծ�����fMD�9U]�'4�_=��rQ<�cw���(gF�
r$Bo��&Z`���)1���ɍ晽�9G��	��l���87�QV>~پ*bXx�Z�t�Q�r��T\U
jx�I\m�����FM��C{{���YB�z�0��heK��	3�J��������2�<KY��Op׸r�@<�tН̽��_�=�N�$�\��]��F~��OV�W ��kQx�a������{z+�O�Y�y�"���	�	��K����L�ǭn
8��x5���O��B�K���$���"(��a�S]��l�����΢hk�:�R�Y�R���6v/������U��n��a����N��g��X�����Qk�2����Y�kS~������h�~�+�*��-�-����>���I�Y!5�7�D��<O�_jh�|�l�|�k���Ɇ��$Yk�˾(�0M�hDq����o���7Mz�����G��P̆� �=��F+�8I���7D�4���t� ��+`��kMPRLm�C�#�8|�����_���WPlJ�, �w��h��]JU��&�Q���(:���ˮ��p�R�1K�(��o�_{���(�a�Bc5��d�.?�� 
����']�߀Y��_1*OvWj�A��ʰ_��q��g�����p�9zV�H�#�ٴ|��ӷn|<������������q%���S��:�{���˕ g`N2X��-%.���!9�K��o�Uݷ5/�}���n{�?+}���!`V"�0
ÁgT��)��%՞E�8!K��5�7�k����S�*��BW�;�f�B�X^�u��H�&"sE��0���(7�������[��c�~)U�9"��]�qO���k9�VJ�M�� �[q�VO<s}O�yk�-�ۂ��.�u�E�6�I����<��)7��
��C��e�L��u�a����*�!�/��\e\lM�&��b�W��A��Wl��\��OV]��D�W��fhq9FA��x����t�%��h�P���8�����|��l��j{I����)3F�O2"'�;����"3�XW ��i��x��+}���C��/Zڌ����>�m�yh"�mCn��^�8_cvټ��6n��3��Z�+Z��3�\�x�o#�z���r
 ����}�Ȋ����!�":�Q�ǝl��9o�4�y9����|�2f����ki ]s��(Q���O?����"�==�㢈�^���m�rc�#��7�-���9�1DK�%�j��$��z�Y54l��&��ŵէ���IzN����P�z�}��8��J�G�,�7��%*�v��0'��X��yX�[桭�hr��9B:K ��s�����}t_�a�.�{�L�Y�<���b�ߙ�-����2z���b�d���"{�1�X��$�����J�Ѝ<V*[�|�0�z�-�P���V�C�-�P�rf�R��p������a2:��['��۱7(a���&9}8!|����% ���i��{�c�R�:a�h?N+�����H0y�`&~u���<7�5b���s���e�w��@4���_[���C�\��o�rs��ʒ)��M���fϠ`w�Lk���XE@�5�K�g�H?��u��0�%a ����y6%_��b�,��Up����!�����)��;�E�������r�n|T4$���,�G����|�;�[9�gsE+����{���E��k�?3�"�/ֿu��X�!���jY�g�rEQ��+�@�F�2����o1U���@)�D�1�Q�]�n{�f��X~�í�83�Z�lV{�I�*��8",��a���m�\��W1��M�ߪ��x��(����n�Ż7���\��~>�:�T�|��ߗ�F��O�nZQ�T���gM� �4��_{��a�5�t���ܡA(vЀ�V���Ñv��Es�m0a6���
x���t��@Ձ�ǼԂ܊t�n��:���
����Y�p�-E*{��xȏIY�¦}FA8X�N"����94>ǠH�!�~d�s=6�Ֆ�@��u���J�0��+w����`j/���G--�)�8�Ȉ{
;�f����;�H�t ��S)����W+���/F���������f��_�;}�_�Uw�gR�!|KZ���]��g)�	��y@�S���;Mf�I�AHu�mm�g���U��	Kip�K_�h� ��׍�hBi��A]ꈍ���)&�x�Za�B���A�РA8/!bL+Mk�.����=G��;CܖtE�"��~�����?�*��D��:�m-���>2ިt,�p�-����v��P$�r"����Y�s1��Yڒ��J��e�'Q�`|59<[����&C��?1���X�ӸAR˥�+��|�:ʃ�8�<~�O����i+��VnQ��j��l.hqKS#0�Pn����S�EU!5�o���z���L'�G�|����ʣ$�wV7��L��O{�f9&�qOm� �� �b)�Sb�����oy�!{��)���sB��ش���r�~mgYp�J�_���:aG ������ȶsCIvqI3��$i�Dq�ٸ���j��Pm�1�Ê��hF�]���b�m�\�7j��J���i��y��2�����?Οa�qJؘ�f���k$��diۖ��ы�#$�=%K��Dplώ��Vz��k���:mYm�S�{۶$���Z�Y����j������Ǧy���r>?I@�/�?H��@w@��O�B�R�&Ǐ%�U��<��L��d�!y�`[r�wզ�
������ΊDR��wE��Tѕ/R|�GĖ�\��	�΃[��J�g~��?�pV�_�����g}�/˾��Td���;������ъ������-�&!M���$PG�	2���F�=^=%^�G��%ri��a�IA3�6��͜��j���xsL����z�J����ԇ�*��h��ʬ��Zp��!j���zU��lvײ<�b��,�o�+�s�|JT������o,��y4�C�K�����
Bm�YA�Oy
\��t����N����r�?^��j�a�ϵ+<~�6�׀\e�[��r|�(�N�^��zwzU]��i�$�٢�U�=�(��Vw����)�o���^�,�C�(������ӯ(�Z&
�8��)0�ҽݗ�/$s)�kʝ��C�.��Wj.�jbS�T�kh�O+U���F��E��B'W}�:�%9��aíAQ�/=�e�N�2j�Ej���˽#�E4or6��&,�V)!(���|��*�vh��I�}�Ϭ�|n{ڨ^Pl�!�����T��`҆9���TdO�v��TYR�l�1q���|��F�]�k�!`@�
�G�{�2��3&��N��`sD�{���A�Nm|e�LJ<���|�Ǿh�~dC8��[I^�+�̈�����o���A�7P���� ��K�5�s-R{I����oi1^��{>�	A�k2A<�.�~ߩ	��]�U g����d� {�J0�d�3�('^���v.�):������.o'~���Bh�Q��_��a�>X�2�p
L�IDf_t�����P=?�d���-�i�W�v���va-<K]4�l#S0���y�I��;b�4X�Uҝ� !Zi����K��c8m��^��m��QR���W��ƿ�L�G��>� !�V�n(���~.B��T�:�ܪ���'Ѽ"��pF�G��x�Te��!r�)e�& �h`1�!O�J�b�{倶�&F��:�Y<��C��2 �q�;�.%A���l�ܫo\��be�Mb��'�ܰ���]�D����r:���d��,�,��܅�o$�_�1�0�w%�-���.����a�����u��#DbU9���*�;p�wH�3���Ф����ܗ�#� K��M�?�F��I�Oƶ�W�j�0��<���:���j�b��Z%Wg�B>�(�[m�pO�97���L�J���%b�=xp�/�i#ɯs{$�9�v{0$�����#�v�[ 2A���;��ڿ�+��fR����Zؐ�(���N���W�K�5��5$H�5��_��Ȩ��x.ymP���1���� }V�w7�/�L��T�1����&���ֵR��=@4Z�;)1�|n�'�ÈՀ��#|!��$�t��(��߆��۶{ZU�HI�o>��F���]�� 앞I����w���MIb���/[�����Q�4Q��8�<��ժ��@{^	()��6��8��c�^�K��ᝒO���dFT�u�+6^�וc�w#�����ݣ>ݼ��D~�W�p��E�U����x��Qe�h=2���O�8�xp|	<����j���r���Mx����$G�W����˭�<o���N����&�4��,g�h���3�W7��K).�#S@����m�Dߚ�E�ە�� /C�9E)	����e���'���=iX�!n���hcM��@��V�K����N��\
;�	n�T�+�u�~Z`Uà��c���k��}q�.��ͱ��/^��8On��Ʊv�ǽ�c��[�t�t�&"c׽UM7��y����	
<튲�t,�����Bq1�W��R��4@mw���U��'xы]��D
�X/�����d�i6~]R�V�L����0�/�g�G���L���ͩ[�`�ڃO1@�r �o�7�O���1IY��Sö�S��C� U��/��	�;�ٌ�'�kk�b?wk��e��E.q6�ܬs_�����֘}*e3��������C�}E�W_��'I��	�����Q����*�{=���4#3k�C�F�r�ag��рU�yI���)\Q�] b���e��v��D�񃒑�z���=q�*�h�s_�A�S*�����(��تb�X�	���b�@�\��.Z'��º�����y 2V�*���Us�o�U:"([עH��^��� 
w��9��R�%�N�	��Rv�g��hd:���6�5h}�'+]6�4*S.iI����� 0�Ϳ���T�O�%-�E��lZ�/V���d^��)x9O�5t�u�@W�8��1U�\���d[`���X�-���79��&{�3�"}z|�L����w"o? �%ܻ|�;v�S]��"s
܆�m�B����&��� m��	:�U���m�3�9S��'��~�B�g�{:�s�	����3���;!CM8�C&��z��4�m}�SX���e�L���4��&%��ѹ֕�W��C�<c�@֨����®A(��9��W�SG�[�DD�-!��c�Z�':�VzLa�p@�]@]�`�� n�� �
�ؤ���u@�q�N��"_	ؕύ�3��a>��� `�+��z��S���;�@Ӵ���Ԗ��n���Wz�Pl����5�d|��!�y�L�	`��e��n7��I1����P�	Lf��t:\?�4dTs���Nⲷ��t�k�_2���Zt]b���V�����i-`��N��m"d�tQ���>6lj3(C��N5tt�%B�4�֤�/e%Pҗ��|�[�ё���E�7�L"�:u�����}8�hO�貿d,�_g�ȶ
�ۤ����9uJ5(��c���#���f{���%P/��q��΃V�toE2��7�û�¤j�([��	r�U'��Ɇk��)hÇ������M��#��*u�u�l�X3�x�
d����Q����Q�Z��v��L���=p����̂��*H���T��aĿ1fȷ`<�-帻��Y;���Z����&��O� ��F�QkQ-�g�K���#
��y
;#�2�R��W��U�̴i9g���hT@� ��^B�Wo��m�:��ErA+wh�bY<{���V���K�X�h=v��&��#:/��뤺��.Ȁ�wuR��%lތ���I��>�B*9�^�ǰuf�'���u�d� Ujx}m4f��x���[$�-{�7��"λ�|�>~�\�
����"�����H\�A8��v���SF���t�#�Dz�3������5�RmH�4י�,Ց�(*=/�Rr��\�!��=tc�LUl�B�y��)V��ԩ��?eW|�+v�7F�����^W�U����G��8�恂��"��;�2kɜ��=F�T�TW����.@���-���Ǘ�AJ�32�v=ʫ�ب%�E �&����N��ɩ��Π��2�X�.5 �"�l�"rA��E��uA�P�6A*�d��X�B�	�E���r��m�����~�J�O����3$���w�B	�qt6S6�����^1�ԛ��P��?��?GB0՞���U�Jg�-�&~5�����JY�l�0bT�x.�v��:�L	">	j_mp�@s�������J��I|Ƌ�u�䶤�=e�Ϛ�C��-7�X �ʑ����˫O���-�SD�)ʼ�g��ޫ���a��Sh�����Wz�s� Fr��]j�ҁ���E7wb'"�o����Y(&�4�xt�� e���T<Ѩk��gb�ߥd#��w$��9~�a�d�E�A��h=���N;�sr+N���ԫ���I��s&G.�4�Qf _�D��M���,��*�v�>�H��j8ؓ���)���+;M���6B_��6+-Vt��Qu�.
V�����LO���f����3��AW������<Z����Y�!g�����BN<z��)�1yCB����%�ѐb�M�t}�l���jxpqaB�6]���0'PV��s�j�"�U�<+x�qt���)���p� l��N��I��:Å����V��EW_a�n6�s�_��U�����T ���02;��[_��ۮ'p�P>���,Dvd�D];듸Pߙ��E�R)vd~��$&9�\��G�>O��u��-g�c3��+�A����d�c �_��b)�d�f�]K�%���9��ud�����K�QHM	���=t���FR��bi�8���#oY1-�����b�U,�]h�\ Qe�J=\霼���l�w�H���Q�r�E�Ԅ8-���� �tE�?��%���ůHq����x�hݳ�jC~	~�j����ޓ@�d�*@h۳ش@Ar�����	}|z�#��m�?rY[���ĽG��u�������v�e��I���F���k�����"d�[��إ�*)��^�SE��O�������&-�,���2i�@�t��.�+��Z���5�ǟ���z!/Aa�]kFݬ�%�Cx�zWIe�q]��"�w@�xj������'��/L�T�L1o�w��S�?�l%(�����Н��	|�n�'ߣu�2��m磃�9�e4a��a�����M{1EY��c�5.������!�
��8���+�j)�2��k��
�X��k>�淒�~4�}��V�z
̒r��p��/Sp9\� ,۪d���#�CT���-7��K�-N� pj����w�hY���v���so��^��V�Z	\I���:�'��y�ˉ���LwsXe,�d_r����-�&���IkˈtZ����I����
2����e)���}!+�!��5��8b�!�,7�A/�j ����E�|��Pkչ��bo��`S)�Ec�����J���\{��I�m"�D��(1����V����qp,h������d���|9�qjN�YI6`�5������9a�BV�A�����!��C�q��������
������C�����_�Ӑ�B���.�E0B:G\�c��bLo����s��S,���e6�^^W��$�.0@}4�G�4��5�bԺ6������{���e��\�yS�.�^?��|"~ՄO�q��oE�ugY\��M��r�̂wF�Z,����|�Y�M)�S*Z�c`ڟ3�@D~���&�N2��lK1�y�#��Li�ɀ�'�LBϑ�K�\/(�	tKoYS��v��o۰��Z�8A$i`NԄ�h	��8q3�)y��B43awMi�_�uXFw]NNsE���#o*�8���'�)���P�P&EIg�P?!�AS���U�*�>�fh��]�2q��OoR!a1p��Z$���C��;J�I
�+�J���x<��T!�s�r��a�v'{��v����|��?0J��}�MD��x��L6��|�Rͺ"?H��]P_� ҦQ��$��x�����hq��a��y>�����F�5�[�W�%T�����"Γ�J�����Ů{F$&�>("4Cs5���ܒsl������6e�����|<{�P��'��&V|V����{�!�����E(��Dt�4�y�Y4�9�Xze����@����"{,��-��`aY�e�z��q����,`6ķHN�S�zJ#M��=�U7,�q��|�A��� G���d�M
G0 �K�����4�G�a.�-D-1��~�n�H*�ҝM����ܖ�v�$��49�?`NUkP"�!��Ⱥ�:�S
��G�:/�|���m��	V_uPHm6�9(T�S��������JG��o�+MC	#���j�HGу73?d�kx�H+1D��V��*	�רlɄ�(8J��t��d�<�7F�=�H�bz B�����u	����S���e�����Xa��U9��]�3�#}��?,Ww�>�3��Ou
������G{l�]��ƾ�qC��_Y��#:�B�3��s����kw��-=
齡��=�	0�)�$v4U!

��Ԗ��������u�b-/N�+Vj@R	���m�A�/�(����ZJ��ɟ!!��zd�������mi�~60�7�Xٵ;Y�O���ކ��B�I���|`�ͦ=`�鮞�I�K�:V, �(����(��)�\2.;S��ߥJ*�)c!���ұ�$s)�� �l1מ�P&*����kKt��{�=���'�vU��v?�F����X���'蕓/0�״��!3�+c�p��#F�P1�i�����y �ʩ�SdNx2���KH��������Q��4���C����AD�v���W�!�t�)�8���jY�VMZka�@s�(�j���I��d�p���Bzi/��Gd�lL���F�زAĊ��M�R�w=��:
yWs��wWb�'���f�p� E���ȴM�,�?�,��i�j�rg��4�Q<M��s�bH��|}O�1�5�R��r#R���K��2��̑�Pf��B��~��6I�������<��Q�+L�d�����5�g-8M��u�p���<������������
�\�����:3Ԫ�$�%������]�-�4�DwB� �Zy�jWqcg~Pn�� �2�R��~?��^;� �����dl��F~z%��܊�!����s��x؞�l8V,�Zj�Pm�1ß6��4��)���7鶪F�pR�u6�������Tz�c.�c���kGlSg�$�r�x�8r>č�.~<,(�y�Ņv9������ wN{������y��6�	e)��y�j����Ó�u���<p
3,��HX����qBgI��.�I|`���j�i�=z8Ы��t܉�>j�\�#oLg�W��!�w����	��{Wk�m��7�����5��g����
�I[��=M�`��1�N�Y^��;vq�2�~��
��j�"a|΍!w_6�*t֟.
�HIl�G+�l6��a������k�k����T\he�N�������f���>�i��@$�m�O^v�8����Wx�
����*�:���kG"a]N��R�m[Ã��*:ק���B~{071�"wS�!~G&�]��xR��@�5p����	�Ľ ƫb�#��N����F��O�;�r����Z/�4i/�o�����A޶���_޵;�m��K7���si��.*>�^�5p0��2\�/͆�RY$���6�|<1��c	06$���/N�?}�w<f�����r�����d��f�U.�+v6>�7!HTٛ��Wl�z��v3{��QIB��Ɂ_��������ɔ+RǼ���=������Xq���<Hٽ?�z��D+Ь��!q�7�������q@��Cթ���U�F�d8z2�u����p�(w CS���7��?JƒO�55����olsS�m9M^0�qmV��G ����ٓLp:��0��Q�>l�� ��*�z��k'@,�k���v�#�F�8���2�0|��m�D��JP�D�0�~�I(���F��2M�M��eN7�+�`]�4����7)N'�_�0I�х@d��t�nJN�b�K%�;�Z��xh����:3c�7����&��+�Z�����}����.F/�$
���e� `�	�<P(.(���>��O[�)H�������'%bewB�&��L�����Yb��e��1�L��&����O���bd����n�@9���=��#TO�t�D�4}�4~e#���>>����z�Ӯ��A�������7���P1�C��N�`��؃it����{ʋ���f�\�at���=�'�P�.�[P��^'P�X+ӱӠw����x�{ 7��!�߁r��Α���h � �7�ٝc��gY�OS�f2a9��_�1�� �Z6�䬝�I~\��lj9�*�k���ݎ��
\$�}fB�\�l�s�kh��O/B\v#U4j��������nwB���r��ߝ�޽��NI2Y7���"K��My?�y��j�Ƣ9����}�e�q��1��hWH�9I�R6$]�| w�.��A�Q{9�/��L�d��a�dC���|m����f��${���@,�j�� ��J����E�֥!R�Z�����Y��*�$;���>'�D����觏%W-�n-C�i顖���|G>\��:���hv^)��\q�C�r\��z��3V�8f�/�*F�hA}�\��X��h�e�*��H�����JVK�����S��C����I��vI:����ԛ�84�<��O��+a�	��`��v�9>��#��D�g���;C�����\U��6bm�}X���� ���.���c�-�<�#��ʄ:Ï�Ζ��V"P��|�R�Y�
��L�5�ڊr԰��<��2M����#��&�`�蹮є�9��3p݃�$�
9L�a�?�vv��.�-�m^4c���b����f��G'5�!���4]�ա3X��_^�l��WiG)�b��#�+2��ߣ�d���?��٭��.�����g��K�@�Pt�$]�:%�b�B܎E+M�,I�ͺRF>+���bg��9��.�}�b��:~���j]���;��jpi	�]IsN�������5�,_�2q�Qn�:r ̴oaum�7h�i��#o�_���m��M���6��8��B�������l��p���Ib�>3_$=ئxKR�(�1�U�놖Sc�IU��L�,���d͈W�/ 3;����Z��ff@wk���A��f�e����za�\��e՟���S;����U�����'Z�.ZJ�R�&���ڳ�h��P���5�{��9?��U���!є��,Zq�ȁ��r_JH�H� �?lH�'��j���S%��a�d�$�F1��S���.����OJ�w-�?:`�9��m�O~e,�	���AŹƠZ'H��a�=��+����-�s|H�w5���]������o����Aכ�W_��:&o��sN���C��[S�� ����^�`��(�R���f6�ƺ�G���F�ZB��&��`���yJU����菁�����q�p^�]q&�z���:���I�`Xe"켼d�pt�Ol�r����3/*���w���g��1]Ę_ P�f�$k{.D����%m���&��͙at��.y��h��Ǡ����� �Li&�	�����O�����;��zn�P�T	���VM�pR�PM��bfB��0�W׵�W��6pRƫ��Ȫ��",+I�����e&�����c�i����ߙ��H�������IWH�_����3TO�=�@�융�zǗ���5��&hջѼ[�	���ff8�C���_w��x���ۙ]�~��ր"�pT���x.H��{;t;4���
����R�E���,#�]r�>�����1�/��1ñ�(	P`0j�5}�	j7�Є	G�Y�bw&}��d�Y��:Y�����T��2��ip�����"g��ɜ:>��ao�io��<�"��7{.�顅x�#�t�T���b�p�ĥ�Hl�������*GP�AR�oB;���V���g�D�2sQu��z�Z2��vX� f�����so#�ؿ�=����w]��(i�Ů�TK��!BGTo���#�\� �N�fĐ�����MeDթ_�:����9���ė���~�npYN��z���`�X���8u������.�%�����������hF��E�x4Q�F�*v!F�4����8e{
f͘ծO�� p�@Ԣ��7t�#�H1툱����uԄK{,�<�\g��q�;l
�M�:ĕ���w���O!�6�������������X�;�~.~U[Y)/P�sG�Z�s{�K�Ú���M�9���-?p�
xX��?.��D�-]P�%#��b� ��V�:��	�YwRf�6��cV�,�@5{��� Y�t��/�[+@ʆ�cC��D�OLNd� ��D�2`�)Ke�ա�1D����f-'�Xm����d50�_��&
��(�Q\�cL��.p/�u"�S�g���[�OJ}�թ�S����3�J�\w�Y�n��Q�|~n�ށ`�2�^G a�\֓�4�^��Ȃib���k�c
��J^�cmݮT���vC7�3��F?")�St�g�'������^5�R=9�H��u�'BSI}	F P�[�<��-���n'MV�O���w|���F�=����-�(����U��sF���y�4b�Ӷ�c��]R�D��_���ʈ�o�h�Ķ��l��	[3�?U�VB��� /�L:��4�gXc8G ��7�"�UU��!�g��21m�4����%x��u���Hᱜ�Й��dJ��p9qgq�'3Œ��h��F��<��'E�`f=�m���
�tW�����)~EƬ�ڵ�NR�����A�x��*I<Ph�ֆ�FSa��҅�T+^�P�V�q�I���w��uv3�F�ң^ʹ��)ꐩB���vU̥�f'ٮ����̦���.�A��N6r�Җ�Dj�����Н�d���+ۣ�c��������2Jz�pu�����؅[I�%���}$��U3�r�~P����@�F ��9���Rc>K�4���x���V���g��5{�R�[$f~M0��,�~�U\�q�]��2$�[�ûF��y.(�.�-@�rP�����R�_!*���i��ϕZbY��Ú���i�[�?LEߊP�
ݰ֥(�)�v�B~��POw�2��x��s(�����I�&ȾN��*������2di
S��	���.>�R?į���?��A�GMa���8u�cAͤ�5��?�ٵ��e[KU=���Ã�:�R�v��9����f�|���|k�W�]G�V�:|h7A�ga���5fp]K����]��_��
�">�
r�$�9Ȫc6��AC�¼�dGQz*���[GљT$-�&�ՠ7��8����K,�r�% �цb�`ޣ��*�`~�p��];� ca��Ə�n݃��S���@�Àg7ȿ44Ba}F6r.	�8粧���[4�Ϋt��m�>U& ɿpS��i���N�c6�󑆢r]���9A�=Nm7rO�U�;���<V~�ފ�s���O���pZ���Ed�	O�b��5j��,{>1�U����?������������k�d����+� W��S2;1�_�8Yw��r��݈�����v�}��u/L���Hh�v�n��Sg��e�׿R�h�B,��o�?��L�ZW{���dن��ȣjz�a�v���#H����Ӎ�?{�X�8����X
M�l҂��&�/��A�ͥ����sQ������HXb(��U�b���8�7*-ֆ�9�4Q9!���!T?��]��ӵv/n�U[_�H��5)֝*"G
ٽj��Z�m�e�7>D���Z<�Ω��K��bź�E"�d֩1KR���4��}ք�.� ���s.fہ@G(DiWڢ�%�������G��k�*����Q�^WE��R���?έhX_�pݑ�ԧO:�D?01�O!,��}T7�VR��rY��ߛ�lUg�·6��$��`�z�u���;�'�Ur'Ёp���L?��E)5�Č�:�侓��!ttĜ�Ԡ���T5	ˤ�V���ᢒaB�0�k"#�I�lܸ�7���kr~m�ML^�������jn:�xH�[>��j�@3"�Ơ;�̧�������� k�\7:�����T��˖S9?�˥c��Ր����"3!�k����c?-���-H�}l�Y�ǖ�(��}G�MMC���fTؓ�s��l�!R�.Ih�����ƕPj���7��)i�U��+�` ��vR�C���z����ZN�tzܕxY;\+-�P��,;n  _}^��IfA��}��!�YS�]lD�S��$`\��&�7N&ɥV�\�RS.�&C�@��۷hC�&��f�����,��SGXR�R���}A�<GN�!)�k-F��o���S��o��NlE1(�gq�:� \��ƾ��0��$���Q	��E�nq��2�����2<yv����LN���:(�h<�'�N"�x�Yf�P2�/����s��B��~Y{��������rG��.�#�H��/�C���[��P[a��.V��!H��!��!���-�b��RL���B��3O��_�=�pW�-%(��āl,X=7����yτ�(|�SP����gUc����Ͽ^/x
J@��0hg���V��Ki�d�K�U��-`�����-���B<gѲ�����I�ݮ���%"Q�=\A����5��~
]rL�i�	��)"g��Ow�B�m��C����	��Y��,=lF��3?Qp���!a��i�ɼキ�5�w��ʰ���ж��Je!Av��aj�5"�9b��:t������/Ύ+��7i�6�L��݁UYSXu�<]I:˪�_e����y`L������:�u��*;�cV>X$���s��ZV�|�E��񫥖[��rR>`��(ր����LJ�,u)�
z���B�FB���
��G�*�\8?{$^#C��b��Y�F��S�)a����{�B�μM�r���e�v�<�>�Ny�p>����c6��5�������]:�U����C!p�\Śǜٓ��$l���g$+�L�~�|����=A��͚�e�؃0WA\�~"�����<7�VV�Ǜ�t���d�>���(��b7J@�3<����ݤ�����U��e���a�N�A������v�{��ݱ�n�C1g� ����a����J��ks'`#��@�w�R�SG��ԡ���N�j�#�coi^sv������B;��۶����h���# N׏�c9D���Wv묔��Gc$�Jϡ���۪7N和���+6��'�oE��f4��/��B���+|�a6�X7��VD�����1Z�E���K���wP9�U��ۆ(�^�M��+����-fc���
�#�:�d*�2�;J���7�wtY�t�p��K�aH���d���2JK�T@�K~|c�+�g;P�d�V'iWw��L̍�CѮ�7D{~ҷ�Alq�bb�M�>x�tt`�2!�~�=FU��/��|�L�쑖�m��`�k�J�� �I��dh�����;�B��.�HyV1�Ԩov!�:�7!��Nֵ�t�a<D���~�EK�uh�;b'�V B��d��{Z�ȎRIx_��j4��i$(q���L#�Hj�he�.�[������dֳ��#������,-[�瓨���b*�d��F�aWd��+�t�i}%�r�ґd�м����c�w���+(<t[�	I� ��r3��OR��H��ؠx�J�v$o�����6���.�N<F�6�.��x �.�N����6.��
~�e�H�]��a�R���j��d:���D�YX��}s����|�|��!.�x�R�����Y3� *^$���?�bu�lF�j4��M��iq�Q&�T�OI"�؜��B�Ց'=�U�]J;֣�R��D���kM��x_&|�L[���!�(��ٰ�v�Q��f�A�����"�ʼC�3t��1L��)�E�E�=$z�v�4�_)� ��m����'�MՄs!�!������/�D���,��O2_�:L��)Y���v����L^v���֢/��h���ƪ�#k����@z
���3�=[:�!����Z%�dv�|<-�<n���T
mCm�pF.�u+Ä��̀AT{˥��Vb�B�uY�kO���:v^�8H�<�x'���	�����z�	���*�$o����:��p=��a�:d>WLS2�93hL� �{�pz��hj��2Zw��a�I�Uײ�e��و/sS���v��O���N� ��e0��x��x������ŠH�n������I��$s���s2"�ij8(acʎ�
�2��4����uN�H�^�trXTo����`���չ���d�N��/[�cp�kً�eޚĤ�m�8�C�^��f**13��W
���.x�lL�w�"��:W�q�9� u��+~&Q��y�0
0�w2� ��F7�A��E&����+Q���!I� �TL��$:��=W./lg���M�9����J�|ԶBtVd?Jػ(���^�4|J;�[{2瀼����.ʊ)v��5�BG�y�����9�kz��X�z?8����!$���623�g���Yߧ��m{",g��{i;���XN����e�Gn���) ��T�^�Iؐp�H8�����	Dʠ��a�� �#��G��0���Kѳ-׬R?\��cR���!��C.�un�����h@c��P�|;��E^��e0��I*���vګY�֊�$w�<�z~�J���۫X�`V����I�b�V�~C�ҏ��P;�
@m�-�c�<�W����.���4^k�� 6i嗡�$�~ְJ�nA:�i�=q���y�a�<��q�Ưk)�@`��;�|a`�ƃf-S�C�5b��8i��qX�<@>�WRm0���}<�NE����f�O���33�A�-&Z�
���(�e�<��5������(�p0&��2�^!M�=�����XRw�Ū6�IL��`Q������S�+����^i�o'��	��^�*�.m2pzeXV�A9ft*2��9����d(v28�r�vb,F�v�yT�2�R��Y��HTp�HTU�T�*��M�9 o��fX>��*!��P~���H�[���wA������ػ`�?^�@�貙>�&�}�$��ݳ@���o�b����b�]*=\��L�XA�����Y����&+��F�C��	���ե�����}B]�f٤<�.3�MD���1�������zΊ%ǉm�Q�h�l�Q�Hb�=IV�UEP(R�]H�М���?͉\�u�.Pd)^�ẑ���l&e�LpTh́Vk�N�=�O8��/�Hv -�4o��
�H[� b+�5AW�A�;.��T�����] �%Ma݋NA�;����\�l؃�.N i�G*XO� b���q���}�	#�E628�C/��J�(��2��mȾ��Ě�����]��Ϡ����f�gE9�!�{m�D���m����37U�����؏:�T��ۏ3��
k�w�h�����"��yθ�{����4i��Cr�ob�w-�Rg��L�UT�F�s�bٳ�����qADL�yQ�:ZUMl/j7�N_.%�gDJE���P�l�c][u&��`�_��al����zhA�ء�W}�K�(��������yg�PQ�����*��u�xҧ�j�^�1	H��i�!����!���s}���=�N����7��63X1D��-O���|s%,��2�/��xlutѩN^���+|�l3��YJ�g5����l���J�o�0�ai�����N�"��|2�{���qW{�M�0��N ��'P��!������S���Y� M�$@]�,+rیI��9V���p/�oȌ�,�+��h1��*D�t�� �0\��\��2�k)[����f�zJ5���fP�����osLFj�b'����eE�N��%ݵ\Vy�}��F��Aӫ��72��G�CO�4�<x��Ԏ��<��E�\4��fS/e�{�͒�	;��~IY��8�z�~�yx�}d�����v�ˏ���
�;�9�]�ʲ=�%m;Ȁ���㗎vM �@����s����Gk��������0��}�3Ҕ/��=&u-�s���4��>�j_Lk<��o4Ln㣿�6�u���f��A����D��wC�{P� �J�BL����Τ$����H��"�1�Kw"����!������4�.Ɇ���,:�.��_�mHΈL$t�Ki���`noڨS���OC=�ŵFt&VV��t�VG����<#�.�lNNb\��/S>	#�"���nm�\��O�������v��DI�)Ƅ��Z���R�(�&%��w�(G�v�s�1_��>��U'(2��r @�l�A�7�#?���f��Z��G]�:�R�w���n�BB���)�ÆR�(H_9�
qwＢ	��F������<�"j��9��8�#�@[\ʄ�	H����jb\�2�	�N��rX!��a�BUy�
ҕ�CR��z2����»��5A/u݌zY"7�1�)m�n�x�Y\�3݈���/��d@��A�&6�芺 �Fij,���_�Y$D�����r?�O����ҷ�����Ġ�)Q|t����dȴ4�#B.�g�G����*%�x�]J+˅�/�bK��a5�A�i(3�b���r��a����݅������=���_�	f5T��T��!����F�g2
��oh\'�q���X�F�pi5�@�ޏ��������e�v��B��Z�,�
"Uc�i�����s���)ϸ��{�NdBf���-�7��h�fbH�"�zq�\�4��s�2��)h"���ê{��FW��tä��`�#F�JT�����T����^��/-%��ic�!bd��'���1h&�����Z�jwK���{0�6�|�z�<�'��x������cq�4e�"
��*�M��J�ԝ���l1p���zȮ܏�S�i�N�F*�'45Ǝ�FN���z�m�޶��H�b,3P� aw8�]&˙��d[`���5�Y�+#����L����}Nj��ok�Ħ1�SǪ��g@�{���R��|O���@�~0����:�~o��O3�k�;^����sx��,V����Cw@M>!O��)}|_�ͩ^HG��(�3���j����L5o�Y�蚨�ɿF_?��ŞDN���ju�-��i�\���'�w����&�p��"�!T�߄Mm����G��|�9�C�F:�`�ɕ^�����lx��+�OQ��ծa>���|F�>��e4�J��%�.��F5!��H$��SrUH�x�9k'�x*I���{��փ��kl܋��E��D�8�o�`���c����O�.1L�3@��R=_���A�U�`��#Q=�>蒑B�� 2�^_(�7�2#k�R�������6��:��S�҄Q'�54��v�7b��sgsX���f�\,	\ �öa�Q�
��*'�]��ݝ_2[& B�2�־:�v�ِ��R?��G�UKJ�L�����;�g����D���7���0�9�n��B:�� �r��"��x�4p��D�H�RZf+9���O 9�U�4%����h�F$D�:�h���CR�bT!�q�t$��ۧ�]EI%b3R���d�����#����,*"1�����z,z&�AĹ6�Jd�*Ʀ'��[�rTn��h{����O��Z0�m1��!�a/��>��r�F��0 \��ɩH���LZW�W(�^�L�`2a�!��f(��h�MJ3[ё�we���]+`��a����b�;q��x��b��M�?6D3��ڻB 8���K*�v�]�l��ò������I����d8_ڼ+��.B���$։�Q�Y5��d/50�XLϢ���0L���[n��.h��B��o�B��+<�l�L��K�b�x�R��6�I�A��V��Q*tY�v��8���f?�i�	�Ve������IѺLx�?M���IQv�o�x����u8SW!���k~p�)J�/;l_ژ )���C�O��!�>{(UJ�23ő��<BX��Ē�,y��n`��Mul���X����'o�]����$S�z��ߦ*�Q�{A�E,�s�^9�&�&/֞jj[.��^z)�;H-ކ�c��i5u4�b�\�R��_v� ��r�j?õV�e+���\�z᭵`��n��s�֞�Ը@ߞ|�9�CyJ�De ����w������b���
����*�t$5���fҎpbomr����5��/X� �q,`�̞�3��Ӧ{�iw�7l��,�����W�Lw�Y	ǀ��س=ɋ�*M��YZ����4��o��{>���y���w|C���x����M)�Q���jZ[��>��((��p�x�s��p�N����<�������4�����,�IY�Yk�nae�4�YI����#}Փ���x��G���s{J���\��G�{�6�=���CܝV��x����γ�z	��1��M�y���g�*LSh�9�&)�2��R'd	r,��l�Ϸ/w5~o<9bA"4ƹ�PM\�	s.��o���`8Ԓ�����Q�Ia��B�!o�6.Nd��ޯa=iv�ti����=�Ն�_aI��_������=�2��Aj�ز�����W��������$Vm�Sg*�ԕ5������P�b������!�3����� �5]v�]HP������:\�� 5JF�_��_��0a�%#<$�e�G3���E�y��BIl�-� =�s ǳ$��!�~a���J�ۇ��m
�����9�šD���L�����xv�����tg�h�J9O!q{�����'�0&�m�zG!�mD���Ʊ��I�Dh���ԩ>+ϥ�����յ�L:��J���Z�\u4(�Ɩ��p>ڒ��f G�m�@s�y���!��8�����=^1����Sd81��d�:�^�Vʠ*?i��Ԟ`��>b*|��XT'�'t[#�lCB�� .��z''�y�������ʹ?�.��^�3���B�����r�^�(#�!�?��1��6�'�HP��X����7��<�=;1�A=׽�u	 >3D�]��0���F.� ��5�9������:��u�s�ҀVs�܄L�	wuLȵT2�򩱖z�k	Q3�`�,��D��K��EH?,�"ˍQl�����!<��;*�S��y����V�hP
$� �m4������� �`�vD�Ϋ�m5�$t��8�G��q���8�
9��+ӏB�$�g��ϡ0�uǙ��~
���f��ձ](�٣��v���n=h8��="�E/XцD���F���V���Us������nH*����U��v �\Ҥ�ec]����_�_�:�S�ų� h��b:]T<�����:ϔ@'��e�����.�k�u��d���?=�����@z{�b�*�٥3x��(g����N�0Al�aM\���^,�b#����ߵZ�]��L��l�K7�`cx�[�m���c���z��;�1�{[�z�/��w�{Ey�#VU2�K���j���ݖ�K��n�ɵ��]�z�^g�6�U�`a���� 5�`�'R,���5|GI�:L�Վ9�WO��	��I��qa��~y)a�nG�⁰�keyDؒP�}�d���sf������BFGŢ���qxu�������7�TP��~_{y�~)���YJ!@���5�xT�m메� ��"���@{���8	{�ԖP9~f�{��O�>z� �{b����w�QZ�%�1O;I��m�yu���zHO������f�ʇȼ�P�O��0�*t�R�$���VxU����tD]����QDo��3J.:|38@�y(F�=���ܫ���7n)�B����r�g��|:�K�.��MH*����}D���:.dW��9l�O�����5�\�]��p*��~Aܳ���tw�@D��W��v~m���X\X9�=�&���w_xi0��Ac�5eI�0KH$H�ϕ�N���O�ܶ�����.��Y�z�\��& �($ �G�(ooZrX�f�B*�l[��I�|���H9��t��"���ۿ��4�2�I)�Lt�O����3��i�����ѽ�t���H���~���4ꧪ����F|�=��o{b�A��NؕD�8���ڵ�Y�<�	=��tzv ���y�~n�kBI��N�������Mё��-7����*���9%��U��ę���#��/�&:��L�Ⱥ-[$h��m��/��c:�ғ/,�%��U4�4�ZP+���t�����Ԛ�8�#�Z"����ߎ�0��UzKn�?�F����f�Dqȷz9���џM�JgSQn��D~!��C����*�YIJ�:Ad�Z紾\(��ob��ց�(�r�b&��F3�;O<����N*1�����'gQ@��Н��Jjy�Q{6ݽ3�Ne��0� ��:̥�H�Rn��wU;������/�4��h���݉"[��V���s������Yr0�d-