��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q������o�/�W��s�5F��C6�B(�@n���V�����mQ�b�/ bz�\�����
��F�
��&bD�ߌz���`���� ����G��LL#ר(�����s$n^�Ǿ]~�����%o���@�I��.�46��LV����m��}_�Yc�ȥ3��3-�l�8L�٤[����M�b��PKֈ�V��`|��|��ҎO�� kn�����VZ�gAO�Қ4 ��	�����鯒8��(�ɈlH�HTt��V!ܷy�v��x���y��e[8���_&�����Ilǡ�N�c���B+�8����Tpө��V�+7��+��s�����d���ͮr��#q߯6�A�6q[��M?�9��ŵL
��_�d`"{�f�[�]���Y�C��6�� /�h��U$�j>�*s^�Շ���KӍ�����Ы.\��C	��˹���=p�����l�����{'���]��@W�����/�Q���2��n"��5:�n8���Z"�`F&�1�8/j��ty�5
�6�Q���
^�7$"#RaT��ʇ�y� .L��μ��s�h�1�/��z,ʡ"V���4�\�_؆�2���Щ�;�Dǖ��i��M����O̖a�
.
����[�6��.�z�&� #�����4`\'FS\��sr��:��{���<$8���T67R�V	��.�J�AXu��~���<- T���d'�ƹ£��@��3mȢ�ܱ�}�a�q�(XR�,��oR�'�	�__�,�@�?dr��ȕ�o�R��6���"��P"-D.v?;o�'�uG��)�
�K=��ƎN4N�eSڅG�m޽��H8c�#����W&I�6ȩ�k���@[:��qU��>��E����9���3�TA�����A,?�)���mo<i��S��c:��}G�)��6JѶ}��,x��w�4�J0@\f�TJ[#�d�:3�7��&��i<w���-���/շ@/�lj�sL2'��N�Y��yZ��K�zR���U�Н@؆�Y�?�M�W���aq�kgޟ'kW����lP��z,�D&����)N�(�]�Oa��A�J��WI�4��V@��wAhF-t�K���%>5������,�iݥ��)1��9�$���1�!��G;���h_5{5��I���'ps�D��:>��%@ɸ�9�W�$>O&��IaUN�=�����L
_�
-���h�c�_�BT�}�@�g
�-��g(���J_���[��<�z�[�_2p��tI 7���'�ȟ��!.�j=�}�D� ��s�3�w�>ٖh��?@7�H����a��b�)��M ���3�,���Xj��������{�w�_���'�;M�)F�ߋIQ���@X�lP�r�P%�s�g�z�i^JNAG�c�r~��a�n�(�v��J�K�O�D_ta ��5����Nw|ԥ��#��[@b:�U��֧�sp��k�e/Ǽ�����w��l"�خ���OQH�[%"�ť�X-�f6�nӎ�aZ���V6����Bؓw�A�T��&�*�XPI���doϢ����-�A�4ĵ[n�t�{�_Y�-PL�Q��3��|4
�d���O�#�zD/��n���ws�"���{�e`�Y@�ŗ�g�)l}�P��5������a2M<o��=M"R@���ڿ8�7���]�[��{�l�"A�)�g!��������1H|�L��m��&;�b_�Ԟ�bFmCƵ�ɞw��{u��1�&|���SM�l�zڝ?���1M�S�k&Ǜ�T�v��/e|��v��8���-:�J(ȥ�U�$��wY;���y�fg�_Yˏ��s]�C��J�?�15��Y��8	D��W���UZj-���ﾞ_H9�U�#�u�1� m�B�j#����@��<�K�I��U�.�C,�g���n ���Z
�?�ҫE)�*��zBM~j��8��6��݀�����se�p���Eq��K�c@��������h�p�I.��CzAB�u�W�ً�F<c�/9T@km�ةZ͍w�5� g��niլ=����EĪ�f��h�����"����� Pr�� ί��H7e�,��G�{.���ۿ�0����:<�� ��pp��Y݌��Cm�rG^u(�9�ӆ��%,ʕ��}�xi���[��f�a^�WI���HףL�,/:��M��f��q�HP&�T:k�gL|+��S�|�Y��Y�������P���B_�&� �m�f��&�����9��~�%O$)�@��i\�3����g�5�Ä�VP��n�(����[�,��FV��n���2W�[o��a���vC�пaA&��7�v�_�E�d�o&��'�=�9S�Hro��X/�N���;�:�r��Oe�q^�.wu10-Њ�Sz��P�85Jړ�L!܀��1߫u�̀`ZJ���Dh]5����z�3A��w��T�sM�煮��$"Y79�'����EZ{�]��)׳ګ��-�^T�l��P�۲d>*X�E�ȧ�8�M�ڮ;j=�:��x�Tc|S��֐��r8������6T+��ȶ1�9A*�
R�շ��Ȱ�Nf)������BX��@�����k�� ��X��x����'�(4���K
�qg���p������ʆ��ҒΊ�QC���J�\7�[�N�s����b*��\*c�Y��$�����)��d��>���	(�R��F����䘍�=��n�7r|/���ס߶G?6������m�R��/��k[���WLeiy���#勨�J�y���h;�9S5����)�z�I2�Ư���)̣��K1�Co��Gf��	?'�ϯ��/��M����4�3�B�N"�R��;N�+�&E2�R089/d�U飤i�ܐ�<�7ג<�l!���V�#�g�(�NA��s�K�H�	���T�M�㣹��x�fe�����©	.����̝�;��	m`M��L��=%���()�/uo���\��d&G0i���.c����]0��F����M�l/S�B���	ǕȑПf��:�W�̱^/p�os�~�e�:��h9[�P8Ξ=wv�r�֠I�sJ�ПP	-(y�K�'ztf��	�y��]�/��b�E/:I�����J�Ү���u�"�iکD�j���7��Wu������/x]�t��g��H�S��GT�㔗�<j�O�ir��N�������t^K��.��N�'�9;QP� ��l��zh�r��j׃�ڼ�'�n�]7��� ,�:�@tQ�����5�Y���]��:�'%l�˺h����i^0h&��(�N!����N��MqC`r��J��*�O�һ�����8Iz�=a��ʱ�1V>�
��T�k�?��}�_Z�&��x����*r=Ѿb0WR����-��S5i�����FG�y�[9h�P����	��������ȾSd�|�H�Y���fd�S��h���!����G�l8tH��Og��[-�}�Fw+����H�Q�>K�w����?�9����@���'�O�q���R������vڋ#���`��(I'm��!2°oAD��'B���Ptl4<�0q�<�5-�.���&R����J��,:/bȊ�� `8�E��o�b�P�����oP�'Y���bm� ��Y�pi3+Q����ik;�_B�=���<����=���E�p�yu����@O�Yv��S�AV�4�&z���Y�o��LGt��l��)�(�˘��ƃ�=H��o���3^�u�ܥXP�!3ۇvo�|��袃0��Y�-�F�������e����K>5�J����7l��頨��eE�z�\M2hA�X8�1�&�7'�;>��9@�uش�
L�mL�O+����j�R3p��Z� �n�
��f|>�$��o^3�G�x��Q�"0�g��Q3a������80ܕ�(����Q�#�/����)��n��������,,�nc�8�[�q*)=q;	�WJy�R09�z@������ĝ+��
�vQ�c<�Qp9�ؾ��h#��<�P�$G��T�����Ѥ~���<��88��C�Fs�&�is�Ƨv��
���8���* IS�9	����/�
b�c�ѡ5	^	�ۍ3��������0�S$��gv_uI�q �z{��Vc���s�,7�$���=��])3�q�ȫ,�<�Ë�����Qȉ�������Kf��R}͚��6�9�H �Q�g�%�C�\��"�OA�eа�q���0�
	��Na�)�l�Ppl�A0=�'���ГXw(a�&b:�/B�����f�HPߑ��2�ς�
U�x�`����F��^-���s��w��W�|�����-�'�0���T��ԑ�
)ua�K�U���2�>��>z`-"9_�o'��>X�H(�5?��D@�>�d\?�W��J���Fډ�6p��s��e*ܝjI�ȫ��Y5����rg0u)����J����,#�P�����,�X+��z�z�}�d<�@�	� IB�2%�o ���|Uq$�k��Y�c�Ə��ɻH����A��̡��+Eʹ�t~��8�o�B��� �j6����� T&3�މr�t ������X��-Yr�1	*�O�����.o��ʇxsl'�+0�O���!�^JRi��h��A�U�(��H��m���r�991 k9���^�"R��Tq��85�����#y-��/��[�ep�����r�'J����a2��^�İSVQ?�{V��2�9�Ӧ��1�`����$����f�̂�v�'Y�q��]�XYB�Ex}��>�{�c�ɨc�D���