��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M���
Q���m@���c����j$���3�1b����}E~��}Ͻ�����8�ҡ,O��@��X�BEls��7?��PKG�UET��B��E|�(ۦ�@Gݚ��1��f\�����B
]�qN+[�9�|�	�ײ� �J�k�H[×��/�J�z0����E���FXO�+�������#��A&0у0��B�>��X�����Ŵ]3�m���;G1uܣ�,.��D�m�d��/G�Uu^���<�,bZ���J�����qj-�b.�g��+6��y��
m� ƈ����i�+O9�g�َ?��qf[��I������?�mW�X�Y�B��MR2�����N2��ֳᐇ ��ݛeØ��G^�x��HN��j#�/�7����4�����u��<��%'�6��o��ZJ\�P��bXME�Y<�PgG� �YZ�>�W���r��@/��
����z~��[!/���ɉ?�`R��)����r�pg�,�R6��|�I�[��yJЫl�ΡF�K�8�4{녉w`�&M�2��j���Ȋ$�DBc���Z�LN!mW�v"����P�5�(�e��x��c�{݉�B����deI�ܢ%���;V]�)l_p�D��6>��#wyJ�$s�(r�N{R�~+�*�9�A����iFVC��G<s}yu��?)&-T0䍞P�&Bs7@h"F�ĩ�`&�Ƕ�*��T��xi�G�1tZյ=�l:�a��0�������pZ�Z`�X$C~�,���h�� Z�>z�C��k�H���f����.�  �+6�P�ڥ��g�������>�n�Wy���[��_��Q����a��� U,.��i���x�y��y��;0&� k������"~���U����Xc��@D}nV�~���#q��޿�� 9�0iY�v�?Hu��R��~���3 !�k!R�E��!�2d������uȉ����[Ɣ��y��٤���|`}��`Nڈ�w p��,ɂ�O�!ib��b���9�Ã8Ai\6�|2�F�2c����O��Ǡ/;%�;��k��Jg{�{ꍎ?��;�ZS��ױ�aU_UX��@�������׼�	��������8����E]Ǌ� Q�z6 K��{#�R��v���P�����_2q�(�;�����2�)7�ۚAOȉ��l�=�!�PZ�w�Z���p{��]��Γ�ɺ����7rrI��}�`�AՌ����Uܢ)я�G���z��\Q�>��/@l��;�uG�#��c���m�Ǟ�����:cT,��(�k�-��ϛ�J[0��z���A�gQ&$�z�ȈfbQ�S��f���Q{:��M�&lQ���&&�i3ٰ+��Ü�x:���N�6 ‛g�״��I�h{��{����C�y�ԅ���ZR�Ҙ��0 ��iq�P#T?��#-�� � u����2�y��*��1⾩D�,v���5so��������e*a����G�[��G�g�(�9xg;�=	u[�5�@���Ϟ�=}��)��%S�f�-�@�'v�7���p`Nzf�+��;o,	
���&�������� ��;	4���<� �Ȝ]��@�-k�u�lI.2�� >
>.���,�,����������"���쮎��^�iy��6�\?�����ֿ��A;�Dv�lQ���<r��{����e<�}M]��*�'}�L�����%�ŵ� ��ϥp�,��Q
k;t	M�(o}u/���3���h��k�dĐ]�9�w�J�e� �}~X����x�P?�Ȑ7����J�m����Oλ�Hz0wO��ˀa3�m��kgm9�?���	�Tp��'�l�@���gq1ԸLjL=
�l��v��jW�W<�ݢ�.�uo�kn>��e���Kf��w����g(�������;<�~l��������U��(��<�E�!��"�|��N�� ��+�X(��]�����a%#����Qm�(;,׺�[q��Ů��5U��c�s��T��g�DǱĤ���
2�ɮ���{��@�7)��+�� ��}O��m� �ԩ�ʤI~;��-�����=�U�3����;aDC8˩��Tt3b�_��9�;�U@)0Ykz��=��4JY�e ��_d�(�G&��)�E	h+��r�a��!�:�w�ԁ��T[��I�׵�_[a�ea�[��c����;����Ǐ�hV�N����H����� 