��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bdc��NAs|%�\�4ar�W����R�fԊ�@~���R^�ԃ5�9�j�d��Δ�A��$�"�pX&�	�����w�/~�>`��?v&���e�!��u���Ǝ����x%!�c�?�?ln�H5a�˘�l�Oy-�B�*��<�kNsԮG);e[�����H���%2zV�6S���\��m�\���ۼcZ�����M���ѳQ�4~'ť��x�dg|)�p��bV��er�л���$�6��3��Ӌ�J��!����*���9̐�!U�@��=�
�J��c7b䪈<��#�tgX�:�A!��R=e�Okc��]�҅ob�*�?k��4�a�����J�������T�p^o�T��A�t��E�����y*�Z���A��N�z��4��m���Qsk�?�?0���D���ŧ,߰[�8��:`����	�Qp�qc:JW	��M,|T�s���ö�}��r#j�0uhO�?�m�h1*	�>r*<�e"�T��J���P��=�u�D)X��r!��Ӧ?��{o�T������?�D�T��̸D���ґ����!5w{�����>�S��b���y�F@���>*ra�0����ɘq"�w�6k�Փ�F�̯�w��b^i$�qE*�+��[یPBoy� Xfn�̊C�B�;���@�,cٜ �s�5T�~+�J>,��O�Y@�ȁ 0��ʏ����
̰�DS@�ډNz�~�.���w�zW����9\g���2� �S��͖x�:OĐu��}��w�϶�����Z��>lIu��ET�Ih��]��Q���K��v*,m38�|�T_3�ء�a8J�ܟ:Ϗ�|p6���h��r�a�>���l�n��q���h�_��H����������jP���>c��WJ��۹p������'�/MW�'ݎoJ�u[�=�9^G��v;B���2D�*�gY��S���.�I<<��*� Z:���
���&q��u���7�Ds�eSZ�χ:T�hg��fpǤ��e�Q���p��u�d���kԏ<��4��T�Rb`zf�,���d�ID%��W �4pZ���Z�P'��g)�k�E��Й��.p7������� �Ҩ�r�` ]�&m�_��%����8z�6��V�n�i�T�ΫR��)���BcY��o>`��j��C9��k^�7���+O���ڟ�Y��D�|f�-�,Q2�y�(�p�
D����"_T4WOm���T�֋�Uװ䰹`~�`%F^fY�ي�
�q|v��nqi�ZAX��] \�2�4���nJK�١@3�Po��"���O�:����	{����k���6�+�Z.#�	p˹f�)-���;�E��E�E:�l���u�*E�~�H�X��u��dS{��C�X��ݷ��646���y�Fu����(*LQ<��4o��&J̳[ē�7�K\ڢ�e��.%=��e�0���y��4�#h�
 ���W�Kݖ*��/~O�fl�$�5nn�>����:�8�������|�5I>��oV�_!P~0�����k$��WgH��՝7_Ӳ��$]�#�)}R9#�X����O%c+����K�%x���ʚ�����Z�����+R_�]<�A�6�:�)O��6��8l�=N��@-��;
gv�غ*��
�5[�ֆq.�y��򨔩�1���z���� ��a���9 D�v?�mQH�dڄN��("eb�ȵ�`4�A��ѣ��E�64Ӑ隿.�������ȗ��w+�gS=����L+(� �Ex�2E;??��ɮ|w����1W]��*�W����+�Լ��@�a[mW5�BD��SᑻeŁ�c��3���������"��r&C8j�,l����aE[]W�oԢ`]�$��@����.h��$2GD�.uÂ&[�����\+�>�-R��Q^5<�T�݁�����|��5ج>�i�vbp_�N��ݖ�؈4���K��m�>��ar|�q�X����'H2�{<�2.�Hz��(�{��`��%���Al,nm,*WI|��΁yi�}_4�����~���RQ۾w\V�W���t$QcT>Ϝ:�����}�Wy�GE"��?q`�r�1F����lj��(��rs�ڛ���[��3��:;��'HKz�37ESv]���R̋b�l����g8DM����1�A�l�K���!΁�O�G7NJS���BB�0=�Q�У�t��Yу�7�r��Cg��{E��w�oŷepTVx�����n��ݪ�A�p�4	��(�y�����v:�B��H��i��#��'�0B��
���}�wᓠaE�<6̀���T�ccYb�M�5�s�cm�P�
s����B?��3,�yW�N<(>e�qj�SU�]����K�sa�[dȬ����Z�s�j�Ȭ
O�}���"�}��"��M��M�lEk�Y�Ҡ�BZӺ�w���V���H������B i�E�l�rT�W�%f]*����Z����Ap����>������i
���I�������3�SxP|�Ed\��j8���R�-�q���&�DA�9�*�����[9�|�Mxj�6T�c���8�Y �E�m�M�݈H�}��Q����?]�L��O�����yҳ5*�KH�u�����jq+��_,��6�����FS����TM�MV�%�M"lg�
�o2��m0?�$=�O��fd��-�}�#�-t��%I��w$��w;T�K�.����}U��P�}<<�k��&D�:�j�������. ��^������]���vH���Ji�kE��6�!v������+�1]��hƞ@@���q�=^�k��+�wk�&5PV��R@}F�ܐ���#���%Ѧ�����ӎ	�&2x�!�f�eH�/�}��� �Dc-/�̮A���L��R��NgR`K�ޔ7\�.�jx֔}{ଙB�Ȧ��sݴ-�I�-f��z��rLG1wMA��D~�&�M����oA�艊�T�q'��d_����gߠ2� )H�	V��snK�gj�m��,�t���٬wu�T	j�a�i�O�z
L�G��^!�Jp]q%����ȓ!�����wx�-@�Il�q=~��YL�E]��S�;��V�:QΖ)�Q6z8Gg9_���N�����X��)I�y�����b�㍤~�����R��~%�g޹?�P��7q�w�og8[�*
�$f;��f�?��"�3�Y_�&�Sh]pRb�(�]h�=�w���uM�ϱ�Ȥ/[���0�t)���_}��b��;ߠ�O�zV��S'7�S���{���N��L���	�h���c�dm��+�����Hw���+m51�>o��采h����|C�o�G�H�
��UC�E�I�$�#s-��"����C8�MW������A�8�C���F̈���D;��c��^^=�;Z�c�5�qI!��|����uո$n�=A��>���#�V�Ӽo�|�e��0�m>��5E���u�k�f�w��U���I��㨇/�8����:V��v&�g��G��H�!�$���H�ʉ�jQh��x��t�uU�DS�c���Չ�'�I�*��6�Tݹ3v�9vO][D�s$���񎠓B��?��XTd���}ză�^��XS������
��B�
GCb0'��XO?�5`����Z��n4ҙ6xjP���"���D�x�stuA�MҔ��D�ш��4�S>�e�oS� `�䐸��j߶�:cUf�,�#i�ޱ�V��qړP��e
83�б�"� ��?�չ]��,X��]*���]dR�E�E��PhЖ��M �sC�g����➮���p�Sv	�Upn���D�@����:�D���Z�7�UK���M��@�����L�"�`h�c�KZ1�fv�U���7�,}�ѯi�槤lD��BXht��ʯXd^�h&�垨���S�4P�\����oR����b�۝��7�!��W1r�Ry�$E8r����[��!�__C�z���!��Gf-�9Z`�D>�99b��\L��s�ղ�y�bә\D�S6J�?��EY^�/�i3i��KI^�P]���>���t�C�Še�� ��w�w��4);7i �ƽ
_��(��<e�L�}�6�m����*�?t�m
W�c�������A��������'��/-��D+�����w�wVģ�\�9! �um�����������T�躔h�Er�
zr޲�2�Ё0��Ѳ\J9/�/!�؈�6�{�H�zMj�΄S_Oe}e�������M��$�j�{#/��Q�F�Z�����2���Sfɠ_Z�3��z�8Ƃ�g%������2;��@�qE� 1;z��7'�0�a���y��sA�}�!��YLnZ&$=͗���$�u����De �V�!��S���7�ǌ��1��T�!���X��������%��+�ÒMFӾ# qH�%b�M����5���A����V���G3n{x�T��	~-�ak	Λ�C��d��8kU~:����6@C#����l��f�g/#
6��]�������a�������1�p�jh:���)<�3���m��r��׏3�c���qY�8j��X����p�)��}s�u�=�.9��l�i! �ۅ}�r�#g%z��?&mK�iJ�~��өp�}m=<d2��g���+:K�0�MK�����yp����a5W�/�1fnq�����[���aVe��7oO�ܗ�,�S��V��&�c�`��q�ݣ~$������k)�Q��Ix(H4��=�W"��gO� ��b�[��Ņ~�I�͎�҆���Hu׭���>8�j']=p��1ujl��S��%5��b�мd`��KL2��L���k���=�M+&��O�����įb�Tc��M7H|])d��VL �F��(��R����Q�f�����HB��ξ��4�Պ�������-��"Cǫ˚�֡8�
�0�&�,�
�(�e����'�I'��a=�!,[lR�3��7��H4�$D�+��~F+t7j\8�
����x���71� �֤W�|c��F�$HM0���L&0������R�	�#"��Q�l�%7)�<�u0<��P�vc��{Xh˹*�z� -�=����Cn؎y��Ic�����е/��~^~zb��ڂ�Sn?��� ��-%�(�+�� �SpQڇ<㝂�2����c�u�����7��~%�'yQ��艛�QlK�S�Ue�g��}�8��A��ԗ���؀}���礠�,�r�d�Cj��vv�aH���ra�)������I^�-���H�e�JEPgRcjp�j�Qq��M�z�0n�<PE��i��(�B�`yߔQ������{�b��'��}��]]}�`qP��x�cL2}��~�ȟ�_�9����Qr��@�7�(=��Q�e1_k��}��E���ZQ�)�/�@`F���x`1�{!�����F`�Ko�XgE���i�	���$��z.���ʹ.�l���<牑��Z�82=kλ�K�w�JB�nZ]ٍߞ8��rp�h���;��Jir�m�O���I!���Ν�	�=(Q� [L��lE	���>Z����=��f�	� +��q��Vz�IdZ�Gf�n�Q�4[�8�L�7���j���2lX�a��	��,Z�E�s��8|�������/E�-0nG5U����ܵߗ�$k*�b��As�v�]i�9��?KK�)wD�:muO�4�q%��*���5fY*��l'�V�xRJ�Vc��
�v�X���WZ~��׽F�S�R����2P�F�J��K$�t��8hKM��O�S9T�t�k��<T9���2U%��LUI0����T�iK�4f�(r��TF���>G�Dr����X����3��1�j�=�<s�B��0>����73��G�EQ&R[��g�)�Z�s)4����8�l�zS�
	v������{�����O�u��Sd�O*����\�鞶� ��Mq>���f����5�NHD�>YZONi?��E�~.�l������n��MT�1�Վ�k7Q���BDPDv:���y7��8�$c�:ن�E���˪i���GDK�b��p~#<�C!��������U�lޣ}�#
�]��@۵����h�_�梮��qI�--p�l�uoG��٫�����(��C���o¥}滘��0fZ�P���ٶ��#8J�L��v���D{o��R�|�(�S�YW���WދN'�lW�ֲ�������{�/���b:釆����92%�MIǞ��B���&[vz�2>�l��(��qd��Q,[�1�*T���L�7Ѱ���4�{�l��Q�"Z/H _��)���<��MƯ"T�� ���E��Ձ������)/�*(EM
eRʨ ��{V��Z.�/�S�I�J��� ��C+�S٢ȡ�#�#��ר|=�H�����Rg=���J�i��Cw�b�[s��MQy�l�+�Q�ٔ/�J�/X3�)_�S��XQ�P;��U!eC�u"�����n��C�$f��꧂��8X&s�����Е7�R��i�(�@��xSBOwQ��1z2�S����r��҈����7��p 6+�F��n�l������:&GҪ���"���� ��6T��:��d��P:���Tp�)�}��^�L:�zAb�ud��9�#���H~���u�zfx286{�}���\&����
/ʲ�Z���z뇴�{+��v[Cm)dj�P�|u��T8r�$��¶3~���1�t{����.q�����keK
��A�3g2��i$fΒ��[H]gtV}��йU2��0{c����`&Pش���"P�� Zg��]h��Q�,������"X�0>�qmH�4�P
I�L�w��CB(��pu�*;���U�{�V븴iF���(����e�T��y�fS5��ִ�1�f�/���m��I����N���~��o�V�ɽ�_������*Pf��*��:y'г?�#K�a�vj��T'��Xw�KI'�mt�s��.�Ѿj!^������%���vЫ�0/:���K��**����NYgY<��� �w�]kLȪ���HE�����o�00�~�{h�'�f���ּ���LPv��G�[(�>fa] ��
�[0=�<�s�8w��M0�&d���]'����{�k5b��#H�A����ˡv�1�k�����|�j@G����i&�f-�2�m�{���!��mI��8��z�l{AM����i��O��^�fuKc���N�d=3G*פ�S,�Q'^Yc��g�m����u��8:�ic�ѝ�e��8;R3�-*��Z��]`N��T��V�]�ǰh��}{�+�~P�Vkz�¤AI��#�[���h@	�:
��$�\��e���Z�'&8D՗�p<�Ź��{�[4���#���ێ��8�������g�����i��6M�6Y����,pۨ$e9��g�����	*
ՠ���b��X���	����DӣҪ�'@Ӊ��=�pE�e�u�#fV%�b#�[_O��:!.���>4U�Ԋ��Wyvg�ӏ���
{a;���僚��U\^*��~8��LL��9�i�!$ ���p�X���&�4�ҷ�)Pg�$��Vq�=���B��e�E<��>V�h�4&��T!&�}��{��Nf�#RH����.{��y}Ö���N']��-1~�"�w�dBB��<�[�{�ö��#��Z�rVw`�6�+����a�V�S�uM%��a�A����xn���2}H<،�p�&�a�<.�n�媇m�r��ۙ���c�J���N'�45��&R���Tv�(��2Y\jZ�v��!�]LO���/����;���4�gmAִF=� ����	y*m���/�x�g��j�0F��^.*XJsn��}x��S��/,<mk��!LO��d	Rm�xt:	�6�"����{��J%�}�>�&S��l<�X�+��X5���&����c�h_�7<a�mO��[����'��:{��[%�Ic���Cvm��.Wྛ���G�x7�b4K@^|������	vo?��N=�h��k���7�7G��2]'��x&0�*ۥ�s#0E?�!a����eأ
�n�8w�(��Q]ӽp���Ƌ �Тo"���鞡W���%�8:�l�����z���`VHV>89��D�b$�4����>oM�V)��?V����;���$Ue���W��M���{�eQ\��c��%_�X�WO��_|�����^S������s<۝\��VW���?�l�܈h9Q�?Pꘔ��
ɣ	�bϸ.�4�l;0I7�
��R|������#hߖD0Z7���S�uر�(�}Zԃ�o(�jQ"`#d�fZH�9Y��MJ��d�����)|���t����^�Ɏɺć���+m�}[N�.�Jч�\��a:x�r�寇+�^W�}���&&�]3��¤zj�;pV��
��qh��S�yb�5�gaa���GHB�{Y�7 Φ
i������� ���٩|�u�g_�|�|u�v�i��Zh�g����}"[C��:ʸ<��#�.�DY���^bQ�8'��t��)����ya&)����aT(���O%�˓�ʴC��ץ8�6�$��j\��u&�"�����������ч{��Ҥ��}5�rX&[�h�3�(i4p
f;�d�͉H"���8+�Y	7�^�飦&�D���訨/Zsڞ��V��r�V��,�K-��}1�k�>�Dى�HO�@�wC������)'��l$��C��p��ڏH�	7�.�5s{z%5�\P�����{��uk��"ْuwf?O��x�ld���X��
�(1�\�Ql�KKXM��)t��TA�K�4fuh��S���4wZ��ҚP� A����!�J&�)��O.N�
���A2�{8�5�\�������V0VD5r<��g�.����Z���sޯ�wj	7�Uz��P�[�1�����W�s�eZC���{�D+��L��a�B_�LiA3�ڤ��
CԾ��*��ߋ�/��
��X���-3lT���
�r��Z#�l��2�¼5Ȣ��������"�O�����.�V'*�G�r�8i�K%|}�LNZ�QH�����c����yhI�'y�65.8E��&N�8��s	)���C��Jic9�s!r�ah0fr�(O���IQ���yZķ���A�U2l�p:�l��.�X�4��ahh�D\.9$�0Z�R�ITB�>����Z�W�����5>)����i�G�7�hV��2�՟�O�&��<1R6Q��B$�6�<��,��1�"5j3k�5������	E�B�����X����+Dͷ�܌EҥFN�{��G�'�J��1	�0H��f�+̖f����J�Q���Q�P^��qs&	[��1�VxzY.8y�S�k��н?T�6+�G�PB��sk�[q���^���E���X�7g�h�tS�1�Y@�S���A.T,7�����������%F������T{�~/>~��Y�W�4�*�
�TN^�q� �-�!)�۬(p�k���l��}s\ R\&V��;)'u�:��oE������b>y6�Ru��`WC{Duͧ����9	ϙeC4�ܴ��D��@�Pk$�^;ئ�t�F���]pqBW�4ʼ\$N�Z�!��!�M��"n�(9l D@�	N��8 ����7�3��ɏ��0,��I�#%������S���a�>k��lr�ͱ����B?R]�N:�s��џ9i�0��_*[D�;)�63.[�7r��x��&�`G�{E�-��E�ѐ���C��C����Ḃ���a�H!�	H�&�l�<t !`�e���$d�1�J�LQ����۝!_J�1��=O�j5}�ScJL�ԫ�X�+ַ8�t���u,Q�r���˼�K*�jkL�-���:��T]����,0�Y�r��p�Ω��&�N��nO��8��f1�D�i��[g��Έ-�T�K�,�Ѹ1(�eL���JL�>�g<)���*�g���a�I����RF��o�fs�~b��+��Xl��?h2��Ƥ��+��Te���	4�Bi6�K��M���)ۜ澑����ꛄ�=�y�h {ӥ��x�1�P�o^����v����^S�����F��A��,S�D��ua�g��H>����U��7�(��aL:��u�I1?F𧢩?Ml�|T�j~�������h�8�J����kH,<�}�1��Q`ڃ��qs��[Q��Eϭ����m2����\��O�ܢ�0;1:�W�P��=M	Ê�[d_P�é�,�)��|�$lҪ�� ��2�o0ٮЌi=x,I�ԣv-46ٕ� �f��%�/a��G?�A�a�s2b�k���_c��W_\_l��]@���fjE��>�M��k������,s*s�90���q�A�G�q8�ʣQ�9?�U���^]��ڜ���CI��.bV/���eۡ�<�t��������>|���3�����l�e����^��~����wG�(�t�[ ���55/�N�"�y��c��õ�ʞ6��y��ٮ�8��S�� g(9(�0��%�`Y/�|C"�{��ɍ/�����쬮��/�)U��^Յ�ZK(��V	d��3Qj>"�?��	a��x�8i^ԩ��vX�BY_��!��H�՞y�䑟�Ц�r�1��栄��,3�~X�ߛ����Ψ�?�-5�9�7�g�+W���o4"X�$�(=Z�6cVN��{/����e��q� c���_�stDs�a��}"�9�����4W3����l�^�. ("���.�H���m�m �@��X;��ݟ���'�s	�lVcYW@q��	