��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q���u�W��R������`�LU��4��I�9���v��{���A����UM�X�c8%?<�gŞ~�����Nu�6{f�Xq��?Uo�u9��Vl��K�,�}PΟ�������Қ����*�9m�"����(w�f�A�@Q��Sb�%�~��\�
m�a��u=��֌�G/�n6�1z`ݹ�/�� K�r���/g�+�����c���ޔ�ο�ي�s4�b�=�Xx0��R�&� �m0P�&�|�D����Y��h�9m����N��EPA$9��Kj�'>����ْ2����R,G7����Y?B�(� ���ڥ�n�J�"�7������ۖrv~�}0��[�
���NSw�A��Or=.b��J����a]ZJ���Z&�)ix1{L��O�_ ��k�p��%��{����&#�l�6]�S���nJ����Z�	�:�W�F��E�t͆��BߠW^�!lu8���Z�cg�;�
t��܉,�q"f�n����y�?�DTC�q:l,��������SV� �0�#�&/Y�`�*�S?t���ÕG Z��� ��ެ��R��$�
ݖ`ؓ׳j`��=��%l�ۚL��첓ńI�hd:�r��r��D������D�S%�Rϗq�9���1-�m��rލJ=�<�Zlu��5ֵ��J|�Q8��*bWqӤ���������_�d�!��|�B�`�y��ʃCJ�R�k��&8L����/B��jh��o���ր� `b��Be�2޾�`�
��-5k�	g[*� �D��k��l�o��@�h�i���Ⱥ�rJ������r�C�Ҽ9��纳;�?��L=gܝ��=	�������#$x$�+{{�p�[���(?X����T))F�h�b�{?������q�|�Eܹqt�&Z�g���B$U�Q��; ����gx�\I;��8���n5�3�c��lN��{�����!'��^�D��c�{\sY䗨�2�~5�HQ����_�>w�D�dz�1D���ژ�H��28Sq��y���['"(ϛ9���ʸ*���nl�5р����p�n���^�ߠ�F=&u"�gUh�R� �;��A�A��Kw�w��IL�L�s�m��j���uBs/��?�O�����V,h�'Ѐ��_=��/�Va�F��;��gVG�iM>W�l�-|B��0K�,�њ	M� g��"n=��ڎ�ɣق��'����-�M)k+%�L����u;Í��Ȳ�6�σ�J�(W6���Х���'З�;֔��1�jɿ}�C�)n��,���1cki�\_�[�q4��9w89Smi�\��S�<v)��'�oH��7x�o�����y0�j,�3=Qh=��26^Ǽ�bX��>1�a�G��.���Ej]8 l�� )��E���[k����=Z��懼�<�t�)�J�=�M�:4x7{���m�.p{ڊ�|�� hB8�h��8q�?pn:�<��ܖo�v/nc9��a��$�_m�5�7�'u�����K��J<��"A��Ѫ��߆+G�g��@1��j�W���o�� ��v�k1�*:�f���5>�'B3��a�i�?�0�9n�h�?�ᇼ�tk/`F���o���0�E��r�������$�4 �.����Y��Zl�^S�f&&Pn��Y&��YE2���%��� ��X���Ha�Sk��Ki�$�2���<gD�J�'0H�N�����PnF]��� �VH|H�=ީ�>Q�iV�_�X�g�;Q�W�����+(�ެ̋0��A3��hx	=����<Z�'_�km-�;���v#��F�a�8]��	��9��3c%��A��'�c*f��b�@0p�t��m|焌V6�q�a2�;�E�r��z��H~�<��Y"��>�`��ʃ�������R��!�d��z�OB�������.�p�+���c�4_�"QJ�H���@+~F����%%/eU(�;v���TE�jY��L�7ƼQ째�Fn\J����hƮ��'Cz��e�X �-V��[sWĭX�-�p���
�{���C��0pH_߈��6��՝k�rs�ob��$�W���=PO�v*q�HJ/���
�Dk�)�sJ��0�[����JR����	v��d�X,��֙�0��XE��]�dW�A������#��
V��������쪂����|��x�,u��䐉�8�j�,
�E�T�m}3�\#ƍ���N����싫��+���b���:h@��7>�x�*�\�,D����Cy7�WA ʤ��EU�T��f����}��;�n�_��'e��%jU��4c�cA�o&�J�[�8Cg�J����QC���`�F�B%ΉH�������[�g�^�8d���|+l�i]��Gξv����5�v��0��=Ȕ\��'�:&S�|�ff�ヺ�.�s�+�#yVy���۵�b6���賰5֍j*?����.¸
�n�
�޴)
 xF�n�s8���
z&��1�^\<4��QM����`�n6��!"����w.�ڗ=����=19Mc�+'�K)�n2�ĴР�#?5�6�g��;��vhg;��z�ҙۗ����Ljxt^����
c���mW)�5�,��FZ�E�`�a* �J�	Q&����ڪ<0��.�֪7�Ԅg��8Q����2��9<��ߩ&�)�H�J��k�v���c���6t���>���{c��t���'nڦ����>&�c��g3檷 �ɿF���3�y`���q]e�XށEVQ-Cm6�h�.x��D�YT�� 3gS��D�DRU�ӓW�����B����~���i�W��U��Pj�k�_T��G�Xƍ�;�j�*��\���l�ϯ:l��Ќr�0peߧ��R����E'�4��u��#�hB��۸����յA��_ъǲ�=��D.��/P��kŢ�W˻�E3}��h�q|N8jW�۹�H�;����P�����w���,VO�s
��'w�r��k���%k5�TE�[����z���T�$g�o���m��;��މ#R}��k+�gC��V�����8���R�w�)�;���f�x·�I~����<t��;���d�Ο'5�.)<�%����8�h2�đ/`I����ǘi�7w2�usGQ�{˛��8"�U���h/���Fqb�2�.\���z��5���]�dp��Zi����N0V��ߜm��>��K@,�J��2^/�T /-@4ﴐ��:t�k�<Ko��a�t�F�X�Nr{Y���Zc�S���t4�u2|�������-�+������ȶc��g���0>����^����0��0DЎH?�3�2�ܔ���M��o�J�:V�z[M�q�4����UF����p��I�"Z�Х	q��n6����WNO3w��&��qz���C�X�W�[$�Z_�"-�~*�kEx���W�[�s[;�Jb?* X���e&����ӵ�|��+̀j|������:P��߲�)*,26�6��i�-�"\��f�������
��2���v�U���>c\����xw1?qjo@�*]��N�mK�.�{r.J௷����/��)ء�)#�/4N��g��YL8�^,��dl�E2 '�!�x4����/5��h�В�+���f\Y�r���������	]��$�����0:E��tNQ3{\C�LY�V�)Alm�	wM=�E�a�At��JW�\͞ka�/��^�@�ֵn��e ���r�������}x7�3vj��^�=�+��1�\3J7ڲ�
��m��Mf���`*���z"�
�(�#J9��0��+H���x������M�X9���a���m1y�� ���=�N���{k���:���#Z��r��gl>ݯ1t���/��9qo�.��ʓB��4�d6&dӡV̽�OYx^8�!Xa���Զ���p�'q����̈�k,J���LZ�~��ڤ�k ���iAՁ.d~���U���*�O��DIƝA��rdU�G{�o��߯��@�Íj���I��<9�@�58d�6e.��.��E�1s�R��Ɋ��YH9.%�o���������f%��Ud~UH��X����$�I���YU����X��h�Fa0𢡫�h��X��|}e�1�x�ۙ,]��9Z��+zb�v��ߣ�H��:�ؔ�����=�v�܄��B)�JȐ�c� =Є �ސ?
1�b��U���q�}��A���[�ނs�]s0�GV`8�Ȯ�����fl։�׷�LG�Kv�Wp��C�D&SQ�$}�u��8{5uS����s�^p.A�ԓt��%p��s�n��ybD�Q ��
�ǰ�;�/�Do�����j��F����KO���ũ��,ځ�����nb��+Vd(Đ��l��G�
Z�HDh޴H�+����6�Bױ�B���E<��n8��]�m+�h�l�-�i�M���|��U���B��{��,�;Ʌ/����l�,�1��'޻�/Q��
"{8N1"ѕ�31�m�Ԙ�� ����q��Xa03n5P�|R���VϿ��X��pD!\^�i��� �r�������cZ���� G\.V��%��[AE.�L��K��x!M���=���_V��k?��:!_,�kսc.�ڷ�X�dP;*�*�m�c��٤�]�4����o�Q
��g5�y2�I�ECT��&k^35<���=>og�$�Ơ�|El�BA�%��n��(F�Ȅ���?ߙ�m6�����w�ӰW�*|c�٩�:Q��R���E����W���thi�Ć����������^�WT)�����CLC�`������*S6�"�����|U�;\4W/�������80����Cv�zf<v�0wTo���qfއ�5�~Y'E}+�>�3��♻7��D�U m����8r���Rp�'��@s�
㔛�c�T��2���7�V��]��]rnd�]�e�?B��O���А
����[�$��5�p�NŻe��c�@�Ȟ�C�po�_sZ	��oP���3�R"�X$<?�w�18��#��h�:l$���+i�Ud��P���<GFB���X1�@V��ϟ�!����\��;Q��R
Z��뜒�k6>X�{J6���锏l�>�����S�(Np�rY�K`�\�*X���$�TOt!9���轆�ka�P�ds��ԐCd+ZE�j�����d�T�"C�#Q���!���'"!:�b�����z~v�iŰ����7���>�pD/:#��Ӥ�[o���*�M 8]���N*�[��t�e�?�;i쿵��IJ���gh������'~�"�:���7���8Ņ2!79k�� �^��8��!,v�Xgؚ����m�|M��h��ꃙva�oa�f�s��S��F���&������}���d����W�Y��YpM�~�B|�oT?�����]$%�?����o�]o]��-e*���tifН�@N��Ϋ�֚��$ƞ_�P�� %��T�:�����LLaq�Gc�g��4:rC.�(�!}=4>*å�msР���A���?8����O�@�����9bx���0�#"�z�-���F�+M��H��KUi6�G%9*�� ~Ȧ(h�\�+�EӝP�"���
�G�T�z�ç;��*s�)��i�M�����=��q0l*����/�C�9:W��'���rѻQcM+��~S5��_WP=�0��x#�A�,Ӟ4ڎ5|*56������ݫ}f�[&\X䓂�Hw��m�7�y
@�CE>E�K ��^w��I��� 9J�*�_�#��T��<
�ݽx%ym����Tǰ�7��-��O!�SЂ�X\I�Wm��X����È`^Ny�G��O;ErH!����֯�ċ|�������h�������c&Dg�L�v�5�1�����[L�r��D�:�V����/֐/�x�/�]w�)8q�,b�Ȓ��%��p��X��,�> J���7M�o4X<�>����B$�\.�O�a'�N-J%��pl�)!�O{'�o :en��h����3zW)���p��~3 �1���^J �j�� t�+��<���$�H	��.N�ݬ���)۽j�3Lٶ.֏��/u��
���h��C��b ߇�?���j,��T�Mh�˯�� ���@���+���I������H8���&�˭���c޸���v�������S��(��I4`��d0��6snH����bqH`��m֩nT]wb�YWU��9j
>9,N2#�y�
xE���vxO`i��8Ӄ�7HD��W�Fe��N$��� ��by$���UP؎�(t_��iܢf<j=��`Y��	�ɱ������Ϊu���6�Q	��zI��,�^�l_S�<�{l�@��]P���&�=t\w+ֻثʨ�]�
����/$��2-'�, ��N�Q�ao7��O�,��!���v��)�a���46�e*r$f�ίo����La�o�N�'f5�����θҥ0pB��n�ٓ�V��S�%�C7��~]�ӟ��a\�K�	*�!�?Pp֎���?�D����pe�"'}
@bq��o*S����9?�D��x���&.7����w͖�8Z��3�/�0��#���/N��$�,A�I�{��l���Z���̐�-��9n�Q�F(�B�AO��h�@T�b��=�r'O�{{�`do�u��E_,�IBcjc�b� e�!X����4�MO�V���~dE��m��k _s�����(T��J�32!�����XƊ��AD��$�a��.��P�B�<��4/�>Gi��<�-~j2)H]�䂡g���d@ݛg!VPM�EɎl�e�����6E����:
�� �T