��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�=L��4�.$�!��V	�jӨ���'��A����`����������M��D7�.�A6w@Nk��Z�)_}(vB���H�A��U�Js졀C4��i�|�)O`�G�?�4���!�x�i��y����B*A:.�T�]�(��=��m5�����z��F+��p�*�{��k�^�އ=?6Lf��$�R�����Q�$�C����7� �P�~c�C��.�lGaw�~ꖤ0�/�hz=-�'���Ul��\VKMU�z鷃ʴ+�L�G�������uRm�	!���%�HI5�+���E�D͗��M�l]yr�5T5In̮����G,��# X�E��K�!��h��Uj#� �4����y��DlW����%��~���a�M�YdU�$>�ޚ�u��WG<tӫzx�í\_�v5��7�3���y���TX��a�c���v,}����(��nVp���:	aÏ4�v��+Gߚ&���*�I\�|�weKQt!Y��+C{��:DG�[+��*��#YR������W�[ۧ�*P�F�v�p'-��A0�tz�	�����)}A,~�	?(ˤ�%b,�F�]���?�����Iq=����/!& 6e�C^/0�unw��fP�'!i���Xq�`��䥔F��g)�fl3R;�0��e��Cܚ��s��ˏCC�
S�����j;pZ˒yߜv�gUt��R&����$�������<�7��ȷE�D��~�T		��v?3�C0�7�I��]_ �툑��twĪD��H����UQ+_��g�='�	���8�H3�h�,���ś.��iD!�p�+�Cw�G��W4��!_%g����zRN� �6}���N4pUߡ��#��ĀY ��T�b���V�c2Q֐i��-rex(�ц}�'T3��;�I�3�ċ�=�S����!�&�ѷ<Д��w�1`0}j:�t-שy��X�N��8����� ������q4�n��[5�Buo��T5�G�3��3ۨL9f$�`Ǵ����N�����wC������u�Y��?]
;j���t�9ؤ��z�P
�NӍ�|W�Hn7ˡ?����?bT>�)'l�۞ܲ��<�h���^�	a�-������*�,3����b؝�a�����݋��Q���O���Q�O��m��>:���\ZJ���w�^	�}d�WۍEy��!���x���w��᪹>��c>���!��g�d�$ R�����B��>��y�]�"�[���P�3�~���&C��L�ma��T�'�� _���e�t�������!+b�ᚐ���t�/H�n^yÖ�S����4\Hj�j��j:��R�x���T�s��yX��r�2YK����;�0dq�'x��$��� ^P'����4��%į���`���:6L�"�?yx:D�y}ߥ#�_��l�������}ik�=j��0���g�Oʔ����Š}i	=��Q�$��8�>��pH���+��u��,�Z��z���v�L�v9躐Fi0b��L+��)aw���i��%�N`��(�2e�������`d�q��ק�Uq�l@���&JI�8N����2�����ѐ۰��U�>�Bg��Oȼܦ��C���j
[�x�K�p�	�4�S�aᘝ�q.Qpz�!ꕴҰ�]=�:��m҂nB�B�g�xY0��jф�t�To޾(���O,GV͔����$W�D�+��"��s���%���T�W(NUr�����s^h3��^������DsJk�z���n"�����m rwiC��T����3C/�*� ��̗��'�gAzi�X�"F��8���ȈR����X��K��M���A8�kpN(J�sΤ�%��bGO�ҥ�Qvf:R'�1�����fs�۠�7o�Zi�uU����B� �Eo�-#���VY�Pެh�۵t��w���7v�J6Ys���LAA��ܠ���|������0}Aκ���'9��vy;�Z�[^<L,���S+�+�Z�l�e�s�au��U6�R�k�3n(aǠk� ���-"B���'��JrL���8��T���I 2�I
�`2~�G�H���D���ǿ|�!*˥�r:&�RS���{d|�N�R�LH��Pr���vu5�⯛�>�C��	�{%`ۤ�\5���}��K`���m\�A��@!��񰔸v�qj�óe*g����Vt���yf�������[�^(�V-�!Q҅3JKle�R�.�y" �b�����cG��Sarߙ�xT{�,;>u�����*8aD�?'0]
e7��(� <�����}��l��@!����cM�X��MS�z�����8�~�y��=�U�_0b���c�T��"�+��q3X$��߉���i��/�@�mpvy��ׄM]��hm�ҏ���!�ehT���U���ZW��}4[~�N�1�z-�u`�oC����Ca"����l��;d�;�+�@\W��Ra�,�����Jw���R�2u���;�X����RÄX�����^�p��z���ݚh�ZY�� (��:�����h������D��́�'�7�{H��s�Æ۸^2���;�}s@N���q�D�-2��}�i�N��-����+�P��jOt)q�p�S��'B*u�k\�����2Lpg�V�n��H�~t��ڽ������d����>2�N��]�7�ե���'+.1=:��yNB��1����2���_����'аX!�;�)������p�Պ��Qv��\K�k�,�C�l�g�՝����z�4�FK�7TNlK�:�4�~����j��R����t��i"j��\uލ��ý��I�vQ�K��q��ݙ)�hATo/�ߜ�h�B�\�����S.�"A����| ��D�#�PQr�5�I��X/ܶ����w�
iL)a[s���Y#�&%�y�t�ә����9Ξ�	%wEjW����R!yÓ���pA'��>�V(���=F�����O�~ms��luc�fh��7�4A����3J;�)4�4���6����e}؟�m"�&����-j��}�m���R?��>��[��(�\W�E^\�I��z	X��H<�"=s�3���s2 n��n�^6@A<y~$�����zŒB@��@�|l\{iv��� ���@1m2H����t0�H���)��Ms���7Zl��)�I�eQ��@�a�)��\�_��S1^�ֆd��	�iԥ���Y�z��F��(.)�QfQkK�\;������f[��qN0����RS�r�{ڠh
��d��*�r�z������H]��-g�J_�ǧh�[����@4xS�	��I���v��@���N�ϻ��L�`�G]����*�;$�W�i�v�?��v怲c/B����l~�K����_�7Ps�\�7v���$J���~�78���9_��R�(���:�SR�N:[��dg�;.h�=X{����$5���ý7��M6��v��&���J<�i_��k���7�>��ü�8���I�'�m]&s�*�ٝ R1�j��@j���O<)m�;c`�� �=G!��Ɖ#}�.Hy����^ü�z4�t�S�a��La`��z�T�)Jx4�@�nq�D�4�1G�!O�"�b3���S��[��p-4t���U�h�m������D�e�	E4��$"P���0M/�� ]؊ܓ�X�<(�/d&�f���VC�NP��o'�#�|��d/N0���l��R��)l�YY�t�Gp�J� ��ʾ�q��S���\�T	��J�7��o+߅�����*���r�`�U�B�E��!���ֳ:J��Ի�����,�}�[w~�v�@9DR����(��L��0���u[�/'{�g��������@]xi���`8̿�������(EcmB�P�a��������UE�u�0�ؘ�qȈɕ����dK�DY|bY�fP���Vj$T)�G��m8q����w���tE���#�xk���_�;=���XH��g�G ��&i2?)�~p��Si��k�����8 �G�:PX⻁�[�����[�iO��s���rGBuߘm1{Ԍ�^�6�d�����8��_�n��%+:�v~"��|ؔ�\YNe��,�m+-��Y42o�;��=q���Љ~��?��	��#��'x��m_nW���)l��m{�