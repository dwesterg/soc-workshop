��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]c*x|1�88S)n?��m���|���a@�� M�m�,��OL�:��9q��f�|:j��~��$�}�`�;�=&��P)�C,m,�X������9���	��u��K�NdS�8J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\�������@�"ϧ̈́�>�~ط������qjSY�_�Bd71��/
S%'���@H��P��r��ݛo��U-�:0����XS!C����j�{�,��a"t-�P��v/+l���X^�[�Fwi�� y��o�5�3��Ą��YVsͳ'F���E'����	�_1;m���N�ɧ���py.	�[S�{�j�KYL��"���`yj��&Z�p�q� K�V���0�XNN��@]���>�.�CwG����F�@�W���ѥ�Y۩�ޡ��|�uv�\�Q�G�8�{j�޾��Cp��&��j{�V#c�ॉ'�v���kܯkCPŏ;���%lg��$���s�h��n�_
���E�:=]M�#Q
 Z&��nJ�}��\=���[�������[.yK�>G�l�����K�5�i'N���9� �
!jM�j��9�<J>�YB������ˌ�9hr������0}�~����|9�QG7�.�%j��f#�y�m�M��cb�A�k�Zդ�[�vٙ��)��;�v?{�+�U{�ۢm-� �-�{�E�/�@�r���A�ݞ)?`?�h����h��׼!��T�6~wV�����I�䀝ԓ�r�-+cȗ�3A��+�k�B'e�b���@��$�<ҳ�s����5ף<�ޙ[�����_��;�/���Xo�懶}#�;J~�@0y�T����ι�ހ�V*���;#@��F� �떶�̎(hBx��;}`^'n�'zB A4xw��;����Y�� pd�<3ڴKq&��mQ*pa��¾�#�[��R�f� ��.�,�R�A�X(b�u1�v��Â�=\��`P���C4�{kO��ݨ�{+-d���rK�N�K���N����D�
]�FQU��j�hn���g3n3�2\'�V�6�x�=��?#I(�&��Z�t������4��W6<W�*��C)�dRF�q�D
zֲ��Dq�]�3�|�a�¹g�זG�"A��3T,sa]4�s�-�]�&ˋU��I=z��H��HD
d�*�t)�g�z�����R�Ne&k,ؖ��7��Es&%Tvy- ���8��[\x����MI��L��'ۮU�M�>�g�|$ȍ�J@��wR�=�p8����Ұᙣ�*���CȻuA�"�ENT=�7ݐr�H>�MfV�[�H�dZ�Yp�^s.⡷<zU�>�U�3�L���"��뗖�#��:sW�Hz/��~K�7΂�y?�R�
�.kb�'�LȨ�3����&Gnu���o�r�-�4�}�S3�y�:�8߆ �k_b�ұ�͍��84v[SgE�AB�;]��]�^�i���3�1�����T=�O�Aȸ��-`��HB���K�ءI�D<y|�o��#�+�`�@����V mw;h(	K�+:[�fc�Lx��*kL_r�>.�9��6O�OP���W[�C�!������W ����,�W�3b[���/%��cpZg [��.��BW]5�(�I^J��Y�	��x27?�3I �h��j[�bկ5dHB����6�Ϲ��O�b^RD�"(��2g�j�@~R���\�%f�b���]B'���s=��ֽ*����nni�B�0G������s�8��^/C��?�̄M\�b����w�X�����/�s�A"c����e�;3Ky]ϒ��0�	-8�4I�}�5m���Q���~�y.m�'�y"�쁭���������F�vc�o��l�V�����,p��N��0��$���e��!�;ͣ��J���%iƠ0�1^����r�H��;��A�ݜ	^�(p΄�+J���)��6�s��0������E�uy���b�Q��t;)�~��&T��!��"�Ů���zFV�cǜT���`5�����H��O��[:][�`W���B �S;:'��3�*�Tp�@��	_����;\�K��9����>�Έ�#2r��i�J�uX��
֋t�-�wFP���Y@����<���'�8�f\� Δ�6���>�
L�(����ޮ�`5�k�?���������y*_�毖�4m<I.@�B��hS� w�`���`�6�[(�T`zR�F�$}V8�8�̼
�j.�Xn��m�oLt(8t�g%���Y4����,����QR��&��+�� �@&��hu���X��{��jQͰ�Cxe+l�ïB�|@[�@X�\q��W3w�!�X�w�����&-���-�Q_]���.��Lq^��Z(S��'d��3�j��oŘ��N�O#A��S-^4d�*�!4����OЉK�h�������	�]A)1n�%�@:w�|'���$�-UL`%�ꤦ`��-�n��*C�'�TS3�hb�P��,-v��u|%r<�ѣ�H8�������4�|(?�bIQҡ�G7J���H�]��gPw�Rym�I4�kJ�?N�`Wh���.�&��T���Kg�� �d*u5���gۋ��aJ;���JI=������I&l]'F�|��F�F�}'�T)��6:B�A�?{H���2�q��87�Ux�E��e)J�\����-�"ǯð ϷYe��j��WnD��zz4��vpI�ăfC�u�mx(�(��N���yA�J�~��V��{�c�2Xi�Nf9����{�����u���C]���������Q7^�9Ĵ+63���B�~:��J�iA͗Fm��]=?�8�	%�US��f���C����#�N1ܧ�x|�H춁��!�Cr�y���@.^aok*4z�V��U�vR`>�;cM�)�jA�w-�OmlMj�')~�b��
�x8��6����3��X+��"`���䯦�Y�O����.6"eFB��EYB�dB��8Y,��Y'.���A��8	WC]�>#n[V��8��z�I;Túp[�0,ɜ�7�7[��86��I��u5tC�(�����|���6���E ��>�����ͦ�#h���W�\���ԅم�8}ԯ��>No�'c���!�4�М+.+��}���l#��,2(�C��kk��ln�8s"x$��3�/%��c����:+R��#VP�� pP��œ��,(fwo;��Cf�j N��S��EMv\��L]ˬ�]b�a�(���rg��J��'�w��$�,����l㻡�b��OP ����cϳ���X���g�������,�B-y������M�YS+��X%�B��v�-���چ��tb��,��6�<�zB���gn�r�J�Vøhp}��OUt5�C�xq�[�"�<,�e]��C��&5eh㟚����ׁ�"a�&���G��k��sx
ZX+�t":G���1�H�(��Y����sS��c:�9���>�b���@�?��]E��T��8*�:��x
��xֺ�F�5]���Z�g�WO&ĩ�hK0N*s�Zn�N(��ZG�,��q+TS�
��f��xh{�,r���m��r��MX���x;��WFB�ʞ<.�z�^��m��Dj�!���h�U�1�R�Q��U
qt���"��ʌ.�l�1 ���a��Loy >����X� �sgMj��y$-RWk�cR>|m����ʢ=�+��$K�R�w�9�*�#䞥Q��Kt8<��NRB���%�4�?)�5��m��[�)ah&=�R��#�1lL�[	 �$)	@>h�4�ϤN���ͅ�t_2�9b��$��*��XӠ)��۬��a���]�<�
��q3����'��B�Ml��W�����~*+ѯ2���Ҷ�&��[���6��[�^�����muņ�!�q��փ��$���/����[�{�Z4]{�t�,��+~ꏤ�1M*���{95Z=�a�&yٹڞٌː�������1��L�Q�ȧ)�9�|`_��4������M=��S �(/�Ɋ��������q��t$\���e�y�	��0�^z�����?dSeEF���(]Z\E�"]p<7D�-���l��
.EMv)�>|���Xӷr�7��2N�$�ę!p��=D[F�l��W����#S�z"��E��K��0�%�?/W^���+T�̉ln,pLvw�8�����gL,t��[�ˑ�U�����@�����P�5����]�p5Z�)O���P�7��ĕ6�.Q���)L�O�p���L<��Oh~�w~��-���0�:i�����O�w�c�j�xO�S
.>��l⸖���9]Gjʎ�TG&�7��
���ST~H���'U��^��n�Qo���Ȫ��+�U�'��H�|�䫺��� $��?��i%��Q�
QI�� �f/X{$e�y��L.�.+�|ݸ��D����&�7t�L�	̆�][K���Ø.#�d��i��	1��`�I��5�,������އK����WmB?�F�O����FDj�sz�c�i&�\t�}�2?���N����I�a�X���a�*T�l�u��k�⑔�r�����{OV�s����RC,��Ǹ8�
�/�NG;x�$G��^5V���,	������=��<Ca���Q!a��7��s?��%i�t���Kg�C3�O����GQ����'6TU�=)*��c/��g�┃�V^m# �R֒�C����@�L���t{�-�6s�8)�$��n7 4RR���<7]��ŖƬ�2-dX�����X��ߗ�"�n���Ɇ7���T���ƽ�G#�_��J��v݃�$���D�����[w�J	L]=��n�9s����c@q*�0�=
鸖��Q2�Y�!:�� %����y����A�3��Յ��f\��)�>�CUE7Of+��훂`���L���,�@5ڽ���h� ��r�H���'����,; a5:_�+O�|��@���B�~'t~��ȴT峠v;nr�6	�j�Vԓ�`�k�> �:��F���J 
�ӣ�<�v3�h�>�C|3��[_� ��#���N1�7l�u���<{�>��^��d��<��1xu��6��g���u��"���b���D��*�^��O;!Āy9< z^z*+����'�(ж.:n�R]��Ώ�^0	�Vi�	�M� U��hp�����!�Y&�P�����e�nжj�1��������0f	V���xy8Z�	�jh��ؑ��{� �߭ID���_�j��g5(H:F$c�n=�$|/D��'��F���z-��o|��]c�\t�5�����0�	��֫��X�����ԟ0�|�`�z燅��]cQ�ӄ�9���'�Ԟ��c�Ro����,�3OLO�]��*̵4�I��b�z�z=�6��+�J�C��6��ŗ@=�D5-: 6�Y7��a�/��B�u�T[TX�|��9��>����A�ҟ�#���.U ̅�	.�G	�Y ��!�Xv��n�7$`K����s�A��3�޾c	�����TfŌusi!���`������L��Ba% �;�u�?����8_瘇j��XS�J$������R}i�_��Q��j[�y��-�I�ĘP��y��e���d8e�K��]��ȟ��ڴGA.C5�m��M��	1)���6-�GD���b���H�A2`J��#��ƴ!�Z@[���r��/3,���~����Ú��+	�W����G�E�u�ڋ��;�I��iM�%�&�9�>�E�lk�<��0�s��0��j1 ���;�_�=�L:a����.t�9���
ʖ�7��ӫ<��W�FN�j`� T/�?e���D0*�����Q���s;_�{x��nxm~��������9�������������i���������o�Q��
4XtfiGL�DĨ����QC�8�kqyY�S?���9��шf�R�@$� �f�vDLߍ�X����Z���w8m�p�
/�e�s���+������Z�%����E���K^q�%��u�����2W��� ��h'2���[������T}۲�l瀚A"R�Ҟ[���'��s���j�'��L��{A���݇>d3ebD6#-�q�EAD̫�^�Sܜ����K�0f"���%(���J��9�b�ݞ�Y���0�-�g���]A#d�^ғ�����/�4uv���7�ؔ^�+��C�����X�O��	.H�|X��v�4�V`����~��8n��3`U|o��E0'��q��u,� =������Ks�
��i�\��N\��g%��u���._�
����o4�g��/����ޛ� Y�[$�rfR�IN?�zV����<ؙ��PUj�<��o��� S�C�Z�2��u��	�\^�`_l�:�b�����@�O��+~�)�	��;Z�>w�ކ�`E�5���R���9����'n~��|t���14d9B;&5�[z�A�g�ڡ[�N�0�� T��+H6�WEœ�(}:����|��Ɨ[��\�q��g��)L@�U{x���sY��Q���� 0��x]M���N(z�Q�@������%�}q�bN�K#�Mz�Td� F1�2O���/�'�����c�M4Xڲ3�������!��I��?]'5��:��E�զ��͌U�Nmd�x��l8R���{��J}�"�J���,�zX�ҧ��8M��g�\y�_�;&��.T���˜�2(7���tXП;
Q��ZB�X������/�J�ݘg2t�z����Zc���8��$wR9���ϧH>{�;�Fc/�M�{]g	�i�#�pJÐ�e��%3}�z=nnX���5H���1Q0�ka���b��5E}F�ao�9YiI���af�)+��+����K���;��^'���c\7�d�7/;�f�ִ���A+�}[�ď��:ٳ9Xfo!լ���c��O��z���a���'-v�M�D��[�u�m>���O���PC�cv��.����J�%�����o����Y�z�yfe�|"�����1�&FR�����~�sB3z�Iu�B��1�}�%�j���gEiA�&�qD�^Q"�is�Z�.	�a��h}Y��-\b����^��������8W�O��֮Oh���(k�r��S��vs���Z�@��̪h���3�� Ɨ(߻p�r�K�p�͞��e`Y8�&�Ը��A��$��<k*R���%-vS2`n|r��&�]=��a����
)n����WDE��lƬ�-V\�?�Xl��>x3�������mԕ��8C\�S�X9�{��c~͚s#���U�෌ovZ@|Al�zt ��}b&9���kDdP��ōn�y#t���_)�-ӱҿ�R>y�!��a��H�����_�����XNc��gx�w�tG�Y���sz6�v.}�NC·d���,9��tGN*A��(���>�L9݇�+,{�.�_��F��<�I �7��r��P������^���Ž#�̖���yt�6�߱
xI9�Q�i��N��mg���g�G{y$��grr�\�@:6E���h�ʵ[t���㪂��W�)a �	��z��pv�LT�m2r�'�@�4S��kU���,��m��O��#�#��������=���,�;��c� �N�=���Ri��:�,�}*ts��림�Gd�!�/����hB�>�s�X7s���!��v�<lE����(���W����qL~i�v;���R�&)�d�� ��۹�
[Tn;Up����5�|e�Yn��c�%���9��b}�#�_3Ŷ�iJ�:4/�%0\.� c���q	�-*	L�6l؈j��2�:���v����MjH��!Y%8q'o�ֱ���:� ���W2�#��"Ƙ�k:���`��Ϣ��t���N�I�HDg\��?Ȍ7۞ @��������MNU#�q�:JP�?D�f�H��w�yN��VE��82��p� ��﫷V#0�	S�MW�P�K_9���O��?^�.�@�\����,_��CM/�Y��7�p
Y[+P.N1�j8IZtv��U��?�b.%?J�2��jS
��x6�b�+t�r�mIZk�+s%���H�2o�(x.X:���{�s���Jo�~�F����=�:�Ǹi�� �\k	��2��ޮ��4.��!����P�����@�x�w~S���e���蚇�iȏ�